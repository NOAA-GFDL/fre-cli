netcdf atmos_month.198001-198012.aliq {
dimensions:
	time = UNLIMITED ; // (12 currently)
	pfull = 65 ;
	lat = 18 ;
	lon = 29 ;
	bnds = 2 ;
variables:
	float aliq(time, pfull, lat, lon) ;
		aliq:long_name = "Cloud fraction for large-scale liquid clouds" ;
		aliq:units = "dimensionless" ;
		aliq:_FillValue = -999.f ;
		aliq:missing_value = -999.f ;
		aliq:cell_methods = "time: mean" ;
		aliq:interp_method = "conserve_order2" ;
	double lat(lat) ;
		lat:standard_name = "latitude" ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_N" ;
		lat:axis = "Y" ;
		lat:bounds = "lat_bnds" ;
	double lat_bnds(lat, bnds) ;
	double lon(lon) ;
		lon:standard_name = "longitude" ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_E" ;
		lon:axis = "X" ;
		lon:bounds = "lon_bnds" ;
	double lon_bnds(lon, bnds) ;
	double pfull(pfull) ;
		pfull:standard_name = "air_pressure" ;
		pfull:long_name = "ref full pressure level" ;
		pfull:units = "mb" ;
		pfull:positive = "down" ;
		pfull:axis = "Z" ;
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:bounds = "time_bnds" ;
		time:units = "days since 1979-01-01 00:00:00" ;
		time:calendar = "standard" ;
		time:axis = "T" ;
	double time_bnds(time, bnds) ;

// global attributes:
		:CDI = "Climate Data Interface version 2.4.4 (https://mpimet.mpg.de/cdi)" ;
		:Conventions = "CF-1.6" ;
		:title = "c96L65_am5f9d8r0_amip" ;
		:associated_files = "area: 19800101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:code_release_version = "2024.05" ;
		:git_hash = "5d306c05d9fe755cab04eedc8fd3de0d3c8355a0" ;
		:creationtime = "Mon Aug 11 19:59:10 2025" ;
		:hostname = "pp033" ;
		:history = "Mon Aug 11 16:16:54 2025: ncks -d lat,,,10 -d lon,,,10 atmos_month.198001-198012.aliq.nc reduced/atmos_month.198001-198012.aliq.nc\n",
			"Mon Aug 11 20:02:14 2025: cdo --history splitname 19800101.atmos_month.nc /home/Chris.Blanton/cylc-run/c96L65_am5f9d8r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run1/share/cycle/19800101T0000Z/split/regrid-xy/180_288.conserve_order2/19800101.atmos_month.\n",
			"fregrid --debug --standard_dimension --input_mosaic C96_mosaic.nc --input_dir /home/Chris.Blanton/cylc-run/c96L65_am5f9d8r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run1/share/cycle/19800101T0000Z/history/native --input_file 19800101.atmos_month --associated_file_dir /home/Chris.Blanton/cylc-run/c96L65_am5f9d8r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run1/share/cycle/19800101T0000Z/history/native --interp_method conserve_order2 --remap_file fregrid_remap_file_288_by_180.nc --nlon 288 --nlat 180 --scalar_field (**please see the field list in this file**) --output_file 19800101.atmos_month.nc" ;
		:CDO = "Climate Data Operators version 2.4.4 (https://mpimet.mpg.de/cdo)" ;
		:NCO = "netCDF Operators version 5.2.4 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 aliq =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.031242e-05, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -3.526298e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -4.556498e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -3.004034e-05, 0, 0.000136373, -6.854834e-05, 0, 
    0, -5.697318e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -9.464145e-06, 0, 0, 0.0003027733, -0.0001057889, 0, 0, 0, 
    -7.459467e-10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.47481e-05, -5.539358e-06, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002248975, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -1.079074e-05, -6.699383e-06, 0.001128023, 
    -2.658448e-05, 0, 0, -0.0001016447, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -2.415745e-05, 0, 0, 0,
  0, 0, 0.001441931, 0, -7.000007e-06, 0.0008300915, -0.0001407763, 
    -9.438008e-06, 0, 0, 0.000478413, 0, 0, -1.56304e-05, -1.81322e-05, 0, 
    -1.787011e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0.0001312646, 0, 0, -2.393607e-05, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, -5.373598e-06, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0003400902, 0.0006594859, -5.393656e-06, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0.005057988, 0, 0, 0.0006399896, 0, 0, 0, 
    -6.459188e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -2.269641e-06, 0, 0, 0, 0, 0, 0, 0.0006637969, 0.001294392, 
    0.001585289, 0.001386604, 0, 0, 7.645676e-05, -4.137244e-05, 
    -3.787704e-07, 0, 0, 0, 0, 0, 0, 0.00203962, -8.412631e-05, 0, 0, 0,
  0, 0, 0.001871323, -3.574727e-05, -1.32363e-05, 0.003009877, -0.0002749608, 
    -4.925872e-05, 0, 0, 0.0009390195, 0, 0, 0.002100706, 7.071897e-05, 
    0.0001778454, 0.0003411351, 0, 0, 0, 0, 0, 0, 0, -1.861847e-05, 
    -1.282381e-05, 0, 0, 0,
  0, 0, 0, 0, -2.805291e-10, 0, 0.001306059, 0, 0, -7.707778e-05, 0, 0, 
    -2.846266e-05, 0, 0.001420725, 0, -1.617998e-05, 0, 0, 0, 0, 0, 0, 0, 
    -3.673723e-06, 3.780113e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0006781553, 0.0007617081, 0.001298307, 
    0.001256644, -9.800518e-06, 0, 0, 0.000621867, 0, 0, 0, 0.001036861, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 9.910822e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, -3.899855e-06, -1.726435e-05, 0.001638663, 0, 0,
  0, 0, -1.933265e-06, -4.801379e-06, 0, 0, 0, 0, 0, 0.007855057, 0, 0, 
    0.001595624, -8.862073e-06, 0, 0, 0.0006190252, 0.002313426, 0, 0, 0, 0, 
    0, 0, 0, 0, -6.754055e-09, 0, 0,
  0, -2.709311e-05, 0.0001137562, 0, -2.718594e-05, -1.092396e-05, 0, 0, 0, 
    0.00369861, 0.002634042, 0.00178005, 0.003970406, 0, 0, 0.0007768043, 
    -0.0001033827, 0.0006734019, 0, 0, 0, 0, 0, 0, 0.005570251, 
    -0.0001457037, 0, 0, 0,
  0, 0, 0.003704477, -8.562727e-05, -2.190997e-06, 0.006054154, 0.0007716815, 
    -0.0001624652, 0, 0, 0.002913577, 0.0005159847, -5.480596e-06, 
    0.005474776, 6.288811e-05, 0.0006760852, 0.00194721, 4.179011e-05, 0, 0, 
    0, 0, 0, -1.691992e-07, 0.0006503824, -7.797182e-05, 0, 0, 0,
  0, 0, 0, 0, -6.394059e-10, 0, 0.004283353, 0, 0, 2.684377e-06, 0, 0, 
    0.00198654, -2.56078e-05, 0.007012126, 0.0001450158, -5.060079e-05, 0, 0, 
    0, 0, 0, 0, -3.856489e-06, -4.000557e-06, 0.00119855, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.001444583, 0, 0.001350008, 0.00178241, 0.003116708, 
    0.003460702, 0.003759295, 0, 0, 0.001706085, 0, -2.357618e-05, 0, 
    0.004618625, -3.842257e-05, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -8.778976e-06, 0, 0, 0,
  0, 0, 0, 0.002851595, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.990394e-05, 
    -1.964154e-06, -9.022303e-06, -1.967683e-05, 0, 0, 0, 0, 0.0001500941, 
    -0.0001009434, 0.004253115, 0, 0,
  0, 0, -3.401325e-06, 0.001596875, 0, 0, 0, 0, 0, 0.01059098, 0, 0, 
    0.002170452, -3.101725e-05, -9.22965e-06, 0, 0.001962234, 0.006231906, 0, 
    0, 0, 0, 0, 0, 0, -7.771783e-06, 0.0007294245, 0, 0,
  0, -8.412508e-05, 0.0002598817, -1.327953e-05, 0.000499098, -4.537284e-05, 
    0, 0, 0, 0.009762335, 0.005321773, 0.001833001, 0.008173849, 
    0.0004068609, 0, 0.001103982, -3.169771e-05, 0.002127811, 0, 0, 0, 0, 0, 
    -4.364314e-06, 0.00794105, 0.003307279, 0.0007417429, 0, 0,
  0, 0, 0.00829406, 0.0003150337, -6.138675e-05, 0.008031086, 0.001291359, 
    0.0001904804, 0, -1.41059e-05, 0.006037233, 0.002224813, -2.192238e-05, 
    0.006889635, 6.212351e-05, 0.001263552, 0.005330333, 9.731822e-05, 0, 0, 
    0, 0, 0, 5.34015e-05, 0.002357366, -7.69918e-05, 0.0001989994, 0, 0,
  0, 0, 0, 0, 2.660541e-05, 0, 0.008740665, 0, -1.783854e-06, 0.000910498, 0, 
    0, 0.0043055, -7.099228e-05, 0.01117124, 0.002852027, -7.7242e-05, 0, 
    0.0001435887, 0, -2.056286e-05, 0, 0, -3.856489e-06, -1.809526e-11, 
    0.005707842, 0, 0, 0,
  0, 0, 0, 0, 0, -8.391077e-06, 0, 0.002183241, 0, 0.001584957, 0.009861733, 
    0.008179534, 0.004046062, 0.007306968, 0, 0, 0.002780168, 0, 
    -0.0001154973, 3.290394e-05, 0.009980203, 2.822379e-05, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, -4.780547e-06, 0, 0, 0, 0, 0, 0, 0, 0, -0.0001482368, 0, 0, 0, 
    -3.386326e-05, 0, 0, 0, 0, 0, 0, 0, -4.436569e-05, -1.084148e-05, 0, 0,
  0, 0, 0, 0.004497755, 0.0009773379, 0.0004790708, 0, 0, 0, 0, 0, 0.0018177, 
    0, -4.414801e-06, -1.332604e-06, 0, 6.400149e-05, 0.001182552, 
    -4.627775e-05, -0.000359652, 0, 0, 0, 0, 0.0003009377, 0.002657189, 
    0.009679044, 0.001369806, 0,
  0, 0, 6.889351e-07, 0.006665296, 0, 0, 0, 0, 0, 0.01218756, 0, 
    -1.178213e-05, 0.004619655, -9.801673e-05, -0.0002237953, -4.557577e-09, 
    0.008616415, 0.01336409, 0, 0, 0, 0, 0, 0, -5.919504e-06, -0.0001160156, 
    0.001774996, 0, 0,
  0, 0.0008783364, 0.0004330094, -0.0001029449, 0.00488302, -9.158583e-05, 
    0.001096585, 0, 0, 0.02041615, 0.008415651, 0.002695009, 0.01427534, 
    0.0007693804, 0, 0.01249601, 0.003388085, 0.00399686, 0, 0, 0, 0, 0, 
    -2.552358e-05, 0.01265537, 0.006272876, 0.003120587, 0, 0,
  0, 0, 0.01262023, 0.0006248466, 0.0002516886, 0.009491638, 0.002672906, 
    0.001215588, 0.0004420281, -2.331061e-05, 0.007891608, 0.004041512, 
    0.0002251716, 0.008726074, 0.0006998989, 0.002678533, 0.01136868, 
    0.0003335103, 0, 0, 0, 0, 0, -6.842476e-07, 0.007406715, -0.0001026105, 
    0.0006796707, 0, 0,
  0, 0, 0, 0.0002541424, 0.001173798, 0, 0.01888907, -7.130036e-06, 
    -3.041958e-05, 0.00375054, 0, 0, 0.005007324, 6.76553e-05, 0.02047872, 
    0.006431526, 0.0001926289, 0, 0.001540269, 0, -2.779096e-05, 0, 0, 
    -7.941087e-06, -5.03065e-05, 0.01298359, -2.220846e-06, 0, 0,
  0, 0, 0, 0, 0, -8.391077e-06, 0, 0.004638549, 0, 0.003702182, 0.01306008, 
    0.01149125, 0.009141521, 0.01147939, 0, -2.878647e-05, 0.003309219, 
    -8.096825e-06, 0.00129472, 0.0001088596, 0.01455136, 0.002609059, 0, 0, 
    0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.0003958938, 0, 0, 0, 0, 0.003352923, 0, 0, 0, 0, 0, 
    0, -1.829256e-05, 0, -5.771366e-05, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 5.590417e-05, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -4.53332e-05, 5.85107e-05, 0.0008223545, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -6.127851e-06, 0, -5.755333e-06, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.870928e-05, 0.0004027202, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0.0008577809, 0.002618924, -7.432612e-05, -1.59695e-05, 0, 0, 0, 
    0, 0, 0, 0.00542727, 0, 0, 0, 0.0004248736, 0.001703562, 0, 0, 0, 0, 0, 
    0, 0.000168397, 0.004722255, -6.006483e-07, -1.696194e-06,
  0, 0, 0, 0.004813678, 0.006243368, 0.003434441, -7.140858e-06, 0, 0, 0, 0, 
    0.0070761, -8.752932e-06, 0.0005429583, -1.328411e-05, -5.24391e-05, 
    0.005023008, 0.004567261, 0.002244001, -0.0005081207, 0, 0, 0, 0, 
    0.002020946, 0.01665987, 0.0112311, 0.003301313, 0.001099729,
  0, 0, 0.0004731021, 0.01385983, -6.131199e-05, 0, 0, 0, 0, 0.01363405, 
    -2.192499e-05, 5.577348e-06, 0.0158064, 0.0004700648, -8.437954e-05, 
    -6.635268e-07, 0.02584627, 0.02883746, 0, 0, 0, 0, 0, 0, -0.0001035138, 
    0.00012617, 0.01298759, 0, 0,
  0, 0.001976664, 0.002318355, 0.004063013, 0.01402067, 0.001730421, 
    0.006535065, 0, 0, 0.0519182, 0.01596337, 0.005112318, 0.02796909, 
    0.003448071, 0, 0.04873737, 0.01245631, 0.006070104, 0.0002543605, 0, 0, 
    0, 0, 0.002582385, 0.02010924, 0.02019376, 0.008479808, 0, 0,
  0, -3.339906e-07, 0.027969, 0.00446011, 0.01169429, 0.02511636, 0.02606366, 
    0.002738609, 0.001108051, 0.0007640316, 0.01024269, 0.007973609, 
    0.004201525, 0.01541748, 0.003817382, 0.01117341, 0.0199791, 0.001983967, 
    0, 0, 0, 0, 0, 0.00122282, 0.01856513, 0.005993462, 0.00458108, 0, 0,
  0, 0, 0, 0.0004470558, 0.006275546, -2.887378e-06, 0.03700218, 
    -7.341986e-05, -1.375092e-05, 0.01073, 0, 0, 0.007175852, 0.0008901841, 
    0.03173523, 0.01308444, 0.001961723, 0, 0.004661222, 0, -2.148395e-05, 0, 
    -7.912988e-08, -2.453833e-05, 0.001066758, 0.02528918, -1.799678e-05, 0, 0,
  0, 0, 0, 0, 0, -2.076191e-05, -6.942878e-05, 0.0139739, 0, 0.005906735, 
    0.01767876, 0.02225427, 0.01938672, 0.02284183, -0.0001152263, 
    0.0003999007, 0.004995417, 0.0002615281, 0.005366876, 0.0005160327, 
    0.02235299, 0.005308246, 0, -1.549617e-06, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -1.406564e-09, 0.002841444, 0, 0, 7.268204e-05, 0, 
    0.00666745, 0, 0, 0, 0, -6.084629e-06, 0, 0.0005814361, 7.852938e-05, 
    0.0004650641, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -7.253904e-08, 0.0001334755, 0, 
    -6.276219e-06, 0, -1.613177e-06, -3.963938e-05, 0.0002796351, 0, 
    0.0006265536, 0, 0, -2.548131e-05, 6.481865e-05, 9.045427e-07, 
    0.002435717, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -4.037102e-07, 0, 0, 0, 
    0.0002216251, -2.124831e-05, -3.219534e-05, 0, 0, 0, -6.956751e-05, 
    0.003656478, 0.008832604, 0.0001423761, -1.616953e-05, -2.621581e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.515128e-05, 0, 0, 0, 0, 
    0, 0, 0, -5.792726e-06, 0.001698509, -1.975184e-05, 0.0005227479, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, -1.006698e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, -9.048618e-05, 0.006330249, 
    0.003214725, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.049277e-05, 0, 0,
  0, -2.428167e-05, 0, 0.001215382, 0.004577314, 0.0007327976, -7.316683e-05, 
    0.0002889289, -3.281146e-05, 0, 0, -1.32784e-05, 6.038822e-06, 
    0.01318981, 3.796444e-05, -2.23637e-05, -4.283169e-05, 0.005263642, 
    0.004364987, -2.299759e-05, 0.001711245, 0, 0, 0, 0.0004762974, 
    0.004209742, 0.01891248, 0.0003045212, -1.150204e-06,
  -2.010964e-05, 0, -5.149612e-08, 0.007411194, 0.01149501, 0.01619671, 
    -7.870104e-05, -3.426976e-06, 0, -1.275145e-06, -7.003457e-07, 
    0.01307762, 0.0008419832, 0.005673671, 0.0009492589, 0.0001713629, 
    0.01030375, 0.01293157, 0.007850606, 0.01041945, -1.856584e-05, 0, 0, 
    -1.53844e-06, 0.005588454, 0.04292559, 0.01546812, 0.004395408, 
    0.002332075,
  0, 0, 0.006997301, 0.02496688, 0.00349402, -1.20665e-05, 0, 0, 0, 
    0.01564634, 0.0007347991, 0.003001402, 0.03476197, 0.001048506, 
    0.001417192, -4.813345e-05, 0.03786615, 0.05199378, -1.429885e-05, 0, 0, 
    0, 0, 0, 0.001543626, 0.003654463, 0.03160518, 8.932118e-05, 0,
  0, 0.005223952, 0.009719543, 0.008602826, 0.0221892, 0.004844641, 
    0.01205558, -1.607413e-06, 0, 0.08564024, 0.02860149, 0.03201464, 
    0.0535591, 0.01613074, 0.0003243686, 0.08505151, 0.04456345, 0.00996939, 
    0.0006230657, 0, 0, 0, 4.377504e-07, 0.01206392, 0.05752998, 0.04778002, 
    0.01764179, 4.918155e-05, 0,
  0, -3.350269e-05, 0.06707957, 0.01700777, 0.03717114, 0.05240111, 
    0.05145375, 0.0253362, 0.01377798, 0.004000224, 0.01614774, 0.01213383, 
    0.01771154, 0.02226299, 0.03972331, 0.03086161, 0.03717805, 0.003297784, 
    -1.865353e-05, 0, 0, 0, -6.200306e-07, 0.02009745, 0.08730662, 
    0.01571701, 0.01351138, -1.019132e-09, 0,
  0, 0, 5.477564e-06, 0.0005533585, 0.02620506, -3.173409e-05, 0.08789323, 
    0.002302417, 0.0005094074, 0.03854923, -1.131652e-05, 0.0001033964, 
    0.01415013, 0.00684574, 0.0622047, 0.0197434, 0.004141928, -1.408694e-06, 
    0.008951358, -7.832692e-10, 0.001741926, -1.413326e-07, -8.390874e-06, 
    0.004734713, 0.003713523, 0.04091076, 2.253488e-05, -2.386747e-09, 
    -5.623104e-11,
  0, 0, 0, 0, 0, -4.322865e-05, -0.0001212362, 0.03022385, -3.8077e-05, 
    0.007847385, 0.03177189, 0.03675582, 0.04896417, 0.03100744, 
    -0.0003487375, 0.0001360526, 0.00917691, 0.007131144, 0.0109006, 
    0.001989717, 0.02709691, 0.009788091, 2.333885e-06, -1.11696e-05, 
    1.484417e-09, 2.680149e-08, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 5.539167e-05, 0.006568928, 9.304885e-07, 0, 0.0008007079, 
    3.766519e-06, 0.009686558, 0, 0, -3.66634e-08, -2.672771e-06, 
    0.001214953, 0.0001438156, 0.01652999, 0.006764972, 0.006571102, 
    3.322863e-08, 8.576198e-09, 0, 0, 1.399959e-08, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0003536931, 0.001619301, -9.448978e-05, 
    -8.031574e-05, -1.667947e-08, -0.0001405112, -3.864975e-05, 0.003996003, 
    0.0002146456, 0.001875401, 0, 0, 0.001026237, 0.0002450967, 0.001938396, 
    0.003939075, 0, 0,
  0.001044756, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001211814, 0.00173118, 
    9.69409e-05, 0, 0, 0.005776905, 0.005043855, 0.00119218, 0, 0, 0, 
    0.0006846487, 0.009397505, 0.020691, 0.002599592, -6.381433e-05, 
    0.005185514,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0003462734, 0, 0, 
    -2.460645e-05, 0, 0, 0, 0, -3.03115e-05, 0.003480577, 0.001861204, 
    0.003694297, 0.001704244,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0.001894392, -1.285405e-05, -1.502717e-05, 0, 0, -4.778033e-06, 
    0.001663677, -1.850388e-05, -3.548476e-05, 0, 0, 0, -0.0001021546, 
    0.01094645, 0.006992452, -2.274547e-07, 0, 0.002752156, 0, -1.188557e-05, 
    -4.417511e-05, 0, 0, 0, 0, -1.430914e-05, 0.002695798, 0, -1.207506e-05,
  0.000480319, 0.005103309, -2.359728e-05, 0.00587821, 0.01244328, 
    0.01332051, 0.005504979, 0.004962577, 0.0002828209, 0.003647258, 0, 
    0.000287802, 0.001072225, 0.02581781, 0.008369779, -2.341517e-05, 
    0.002708195, 0.02056802, 0.01112929, 0.002728307, 0.003927482, 
    5.8535e-05, 0, 0, 0.004465845, 0.01181419, 0.02945868, 0.007715635, 
    0.008982581,
  0.0001376187, -2.247243e-05, 0.0003050519, 0.01602275, 0.0247145, 
    0.03262456, 0.005967617, -5.595521e-05, 0.001189121, 0.001883144, 
    3.895492e-06, 0.02226802, 0.008487527, 0.01546391, 0.003360353, 
    0.002651965, 0.02040034, 0.01831551, 0.01243834, 0.02917234, 
    -0.0001345571, 0, 0, -1.53844e-06, 0.01076238, 0.07235911, 0.02343378, 
    0.02119472, 0.003359612,
  0, 3.530411e-05, 0.01769511, 0.06578395, 0.01977609, 0.001273358, 
    1.863302e-06, 0, 8.700582e-10, 0.02899329, 0.02966261, 0.005351246, 
    0.05056082, 0.008115686, 0.004220338, 0.001080048, 0.06576254, 
    0.07897183, -0.0001475067, 0.0002458447, 0, 0, 0, 1.185936e-06, 
    0.04275419, 0.03652814, 0.05521159, 4.902284e-07, 6.606339e-05,
  0.0005781139, 0.03327363, 0.04870749, 0.03276725, 0.03865824, 0.02419687, 
    0.0282358, 0.0009900681, 0.001237036, 0.1494645, 0.1223593, 0.2014815, 
    0.2101947, 0.1733692, 0.004237191, 0.1413766, 0.1890041, 0.02282632, 
    0.006219763, 0.001151519, 5.394787e-07, 0, 0.003394868, 0.1612424, 
    0.3636693, 0.07936168, 0.0222362, 0.0002206467, 2.074422e-09,
  2.116789e-05, 0.0038562, 0.13392, 0.03458858, 0.08337176, 0.1188134, 
    0.0839933, 0.1321275, 0.07673074, 0.0828308, 0.08464128, 0.1004333, 
    0.1576038, 0.06039786, 0.1765341, 0.2085624, 0.09972533, 0.005177381, 
    0.001114486, -7.014045e-09, 0, 1.550452e-06, 0.01829002, 0.1497892, 
    0.3737766, 0.06225493, 0.03335679, 0.001336829, -1.5161e-08,
  3.110834e-06, 4.273831e-06, 0.0002888687, 0.001309547, 0.0378665, 
    0.004877751, 0.1507241, 0.0414666, 0.009604026, 0.110546, 0.0005336666, 
    0.003952444, 0.09174461, 0.09013069, 0.1637584, 0.06688996, 0.0043861, 
    0.0009502077, 0.01562182, 2.491308e-05, 0.006803697, -2.008404e-06, 
    2.445688e-05, 0.05708706, 0.02759182, 0.06305692, 0.003691301, 
    7.461726e-05, 1.260395e-06,
  -7.699029e-12, 0, 0, 0, -1.368119e-08, -7.56433e-05, -0.0004323374, 
    0.04189865, 0.0009375052, 0.02887629, 0.07547558, 0.08361408, 0.1753017, 
    0.06895324, 0.0007861647, 1.080529e-05, 0.019167, 0.03039036, 0.0216518, 
    0.01629781, 0.03537129, 0.01743002, -2.645597e-05, -2.70461e-05, 
    0.002080734, 1.19482e-05, -2.977583e-05, 5.571879e-06, -3.647673e-07,
  -2.268817e-08, -4.516513e-06, 0, 0, 0, 0, 0.001011634, 0.009056396, 
    2.723732e-05, 1.329231e-07, 0.001120432, 0.001817941, 0.0128999, 
    5.299732e-06, 5.575467e-07, 1.739377e-06, 3.107612e-05, 0.006488723, 
    0.00311014, 0.03888565, 0.0287707, 0.04173865, 0.0005826385, 
    1.354923e-05, 5.465148e-05, -9.739442e-08, 2.348846e-07, 0, -1.69382e-05,
  0, 0, -8.191251e-09, -5.487548e-12, 0, 0, -3.715013e-05, 0, 0, 1.21872e-10, 
    -2.462036e-10, 0.009708377, 0.009045804, 0.005238362, 0.004044292, 
    -8.5491e-05, 0.003045129, 0.00473819, 0.01005243, 0.007378473, 
    0.005271012, 0.01130079, 0.007282336, 0.003924779, 0.008619336, 
    0.02608779, 0.01552576, -1.111762e-05, 0,
  0.004227054, 0, 0, 0.0001538788, 0, 0, 0, 0, 0, 0, 0, 0, 0.001335419, 
    0.005468472, 0.003606915, -3.761359e-05, 0.0002156662, 0.02651202, 
    0.01062639, 0.002696448, -5.17719e-05, -2.477418e-06, 0, 0.003021198, 
    0.01866523, 0.04359412, 0.01695774, 0.003926239, 0.009990091,
  -7.263008e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.612397e-05, 0, 
    1.235519e-05, 0.002273633, 0.0005932745, -0.000100816, -1.327345e-05, 
    -9.067003e-09, 0, 0, 0, -6.224385e-05, 0.006267952, 0.006799832, 
    0.007140953, 0.002579121,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.00107171, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.001994516, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  -0.0002398836, 0, 0, 0, 0, 0, -1.062297e-05, -4.431461e-05, 0, 0, 0, 0, 0, 
    0, 0, -1.757539e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001843266, 
    0.00381864,
  0.006750029, 0.001458276, 3.976561e-05, 0, 0.00446598, 0.003188563, 
    0.008205518, 4.701193e-05, 0.0002833544, -4.314431e-07, 0, 0, 
    0.001371633, 0.0156843, 0.01383801, 0.001842628, 0, 0.00668454, 
    0.0009504608, -0.0003563198, -0.0001382482, 0, -7.605021e-06, 
    4.396923e-05, 0, -0.000102231, 0.005699925, 0.001027006, 0.0002586435,
  0.004090916, 0.01216741, 0.002986378, 0.01790701, 0.02985531, 0.04157859, 
    0.01900716, 0.01675701, 0.002536027, 0.004886304, 0, 0.0008558914, 
    0.01331308, 0.05412336, 0.02453016, 0.002683886, 0.01101867, 0.03131551, 
    0.03631725, 0.01170072, 0.01183778, 0.009252482, 4.919337e-06, 
    0.00465885, 0.01184462, 0.0198944, 0.03921854, 0.02368802, 0.01961044,
  0.01180546, 0.0004838697, 0.003300688, 0.04468461, 0.06590819, 0.08946783, 
    0.0547096, 0.01773968, 0.006103409, 0.0189036, 0.02241671, 0.08501838, 
    0.05185228, 0.04396554, 0.008641678, 0.01865762, 0.0678245, 0.05697606, 
    0.03301391, 0.04124653, 0.01296035, -8.864889e-05, 3.99991e-05, 
    -3.308413e-05, 0.015246, 0.1085642, 0.04448019, 0.050595, 0.02384611,
  1.717936e-06, 2.530854e-06, 0.109025, 0.1037282, 0.1363407, 0.06724241, 
    0.02665292, 0.02497779, -0.0001091458, 0.04866206, 0.131682, 0.04904887, 
    0.08269396, 0.09066202, 0.07530417, 0.05748407, 0.1628677, 0.2077961, 
    0.1170055, 0.02445186, 0.002152737, -8.402266e-06, 8.441497e-06, 
    2.644305e-05, 0.115873, 0.1718285, 0.1492272, 0.006065301, 0.0004086621,
  0.0001299385, 0.07156887, 0.1949624, 0.0526013, 0.1131998, 0.08000924, 
    0.1064381, 0.005026801, 0.0005765061, 0.1147467, 0.116759, 0.2020413, 
    0.2591248, 0.2396996, 0.02293536, 0.1726509, 0.242412, 0.1849166, 
    0.182324, 0.02674044, 0.0007364207, -4.857227e-06, 0.006756531, 
    0.1423879, 0.3280472, 0.2434626, 0.06475966, 0.04037404, 0.0006989401,
  0.004264024, 0.06209442, 0.4288662, 0.2156403, 0.1332313, 0.2315827, 
    0.1664678, 0.141682, 0.08465379, 0.05335507, 0.1033719, 0.07945242, 
    0.1254686, 0.05308193, 0.1413365, 0.1935088, 0.1520695, 0.02749644, 
    0.01232736, 0.00788823, -4.429193e-08, 1.278163e-06, 0.04208041, 
    0.4425554, 0.4794622, 0.298704, 0.228803, 0.01478834, -1.291342e-05,
  0.0003158649, 0.02018438, 0.05686961, 0.03456764, 0.113119, 0.05360938, 
    0.2871258, 0.07285917, 0.146715, 0.3167641, 0.02803779, 0.04886332, 
    0.1249435, 0.1224959, 0.1625182, 0.07223116, 0.001757329, 0.005217026, 
    0.02401989, 0.0006662981, 0.00218494, 3.233879e-05, 0.008192024, 
    0.3120646, 0.2641205, 0.1029156, 0.02347476, 0.01074316, 0.01265689,
  -7.322318e-05, -2.624217e-05, 3.933125e-05, 0, 8.77748e-06, 0.0009807851, 
    0.0317729, 0.06952706, 0.004703029, 0.1143667, 0.09393443, 0.1038401, 
    0.1806398, 0.0745744, 0.004301274, 0.00423413, 0.02807443, 0.05148232, 
    0.04047907, 0.0995971, 0.1422667, 0.02822467, 0.004193994, 0.01356554, 
    0.01534897, 0.0001008593, -0.0001485458, 0.01131808, 0.0007679088,
  0.0008081434, 4.107755e-05, 1.125848e-06, 2.099413e-06, 3.976193e-08, 
    2.134331e-10, 0.002133064, 0.01154592, 0.001230692, -2.78047e-06, 
    0.00760534, 0.004017457, 0.02102032, -2.080217e-05, 1.661185e-06, 
    0.0003009939, 0.002706399, 0.034956, 0.05774232, 0.09883808, 0.2013261, 
    0.1553772, 0.02310804, 0.001716907, 0.01115894, 0.000159793, 
    0.0002854491, 0.002017409, -0.0003349896,
  0, -2.265092e-06, 0.0002176506, 2.678037e-05, 5.919548e-05, 0.0002483703, 
    -0.0002142791, 0, 0, 1.09324e-06, 2.187816e-05, 0.02113484, 0.04975968, 
    0.02703717, 0.00813963, 0.002020259, 0.01572665, 0.01852458, 0.02948491, 
    0.02169924, 0.02382744, 0.02075524, 0.02205921, 0.02171835, 0.03406733, 
    0.06739799, 0.03704241, 0.0001300063, -3.015128e-07,
  0.006972607, 0.001554034, 0, 0.0009916698, -1.780234e-05, 0, 0, 0, 0, 0, 0, 
    0, 0.003923582, 0.0151391, 0.01134792, 0.0003443758, 0.0123889, 
    0.04427839, 0.03170381, 0.009008583, 0.002142675, 1.358135e-05, 
    0.0001772014, 0.006829399, 0.02736602, 0.06481104, 0.05244874, 
    0.01840853, 0.01801703,
  -2.991467e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8.970423e-05, 0, 
    0.004476557, 0.005931336, 0.006798713, 0.005634072, 0.00018674, 
    -8.492218e-05, 0, 0, 0, 0.002617741, 0.01638313, 0.01857561, 0.01314321, 
    0.01161184,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2.222757e-05, 0.003489666, 0, 0.004354576, -7.599924e-06,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.01012084, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.044465e-06, -1.290717e-07, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.008861385, 0.001095972, 0, 0, -2.532962e-09, 0, 0.006477216, 
    -0.0001455888, -1.546441e-05, 0, 0, 0, 0, 0, 0.0002518971, 0.0073707, 
    0.004642643, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0004276453, 0.006317056, 
    0.005727021,
  0.01303795, 0.008218053, 0.002508656, 2.169805e-05, 0.01462425, 0.01268496, 
    0.01241713, 0.004583968, 0.01317334, -3.849707e-06, 0, 0.0002589377, 
    0.00349397, 0.0191486, 0.03036312, 0.0113558, 0.00222406, 0.01645656, 
    0.01117584, 0.005964985, 0.0001485378, -2.344885e-05, -4.98777e-05, 
    0.004476048, 0.001938612, 0.0002709054, 0.01574553, 0.009886015, 
    0.008597972,
  0.03050725, 0.04196437, 0.02594152, 0.03955084, 0.08906053, 0.0894649, 
    0.07627521, 0.05260788, 0.03452352, 0.02026551, 9.107612e-05, 
    0.003030323, 0.03371153, 0.1040291, 0.08047046, 0.04443476, 0.04757564, 
    0.09430154, 0.07465948, 0.04577155, 0.04854326, 0.07623529, 0.02378768, 
    0.01844907, 0.02362202, 0.03980953, 0.05952036, 0.04887958, 0.04296788,
  0.02927397, 0.02102106, 0.02415493, 0.08235814, 0.1301242, 0.1403611, 
    0.08278997, 0.02678315, 0.02224338, 0.04352778, 0.06865417, 0.1624431, 
    0.1312717, 0.1715935, 0.03424663, 0.06455858, 0.1207289, 0.1373219, 
    0.123573, 0.1515671, 0.1174872, 0.03968948, 0.03245459, 0.001585779, 
    0.04461673, 0.166184, 0.1061881, 0.144759, 0.03691865,
  3.031413e-07, -1.403671e-07, 0.157338, 0.1023942, 0.1210474, 0.06998271, 
    0.108513, 0.02700267, 0.003462665, 0.07805286, 0.114811, 0.03840681, 
    0.1116311, 0.1190153, 0.1129889, 0.04251197, 0.1602667, 0.1906223, 
    0.1556893, 0.1859675, 0.03780149, 0.01358705, 6.19013e-05, 3.931559e-05, 
    0.09998573, 0.1631781, 0.2006152, 0.02704463, 0.008459918,
  9.677717e-05, 0.05698159, 0.162974, 0.05350477, 0.09018145, 0.06831868, 
    0.08765234, 0.001444525, 0.0001670854, 0.09521931, 0.09879537, 0.167284, 
    0.227186, 0.1938784, 0.01463291, 0.1540888, 0.2165487, 0.1365416, 
    0.1736685, 0.06623669, 0.0629146, -1.538521e-07, 0.00106782, 0.1325697, 
    0.2665656, 0.2330786, 0.08365094, 0.0584521, 0.004579347,
  0.0004361032, 0.04386085, 0.4181174, 0.1637674, 0.1012151, 0.1725253, 
    0.1402184, 0.09765044, 0.06274307, 0.03521001, 0.0655537, 0.06218699, 
    0.07682566, 0.04068243, 0.09771972, 0.1416028, 0.1086371, 0.02222479, 
    0.001487914, 0.001076513, -3.122501e-07, 1.488231e-07, 0.02965197, 
    0.4296911, 0.4615011, 0.2698953, 0.1777836, 0.01313374, 7.427175e-06,
  0.0004355149, 0.008143644, 0.01359909, 0.03131611, 0.06805327, 0.03508081, 
    0.2358774, 0.05218082, 0.09896841, 0.2651633, 0.01567993, 0.04029545, 
    0.09230871, 0.08054497, 0.1323167, 0.06006759, 0.0008269316, 4.93819e-05, 
    0.02145224, 0.0003327488, 0.0004498432, 0.004073411, 0.00270372, 
    0.2244351, 0.2027602, 0.09566417, 0.01295444, 0.01591483, 0.01218581,
  0.002745572, 2.873854e-05, 2.44714e-05, 3.806631e-06, 1.594602e-06, 
    0.002632813, 0.02115496, 0.0551754, 0.002416593, 0.08614226, 0.06793613, 
    0.07371978, 0.1523536, 0.05866375, 0.004614444, 0.002089585, 0.0156671, 
    0.04215267, 0.02796186, 0.07207364, 0.103294, 0.02748789, 0.000389567, 
    0.009746588, 0.004918355, 1.052702e-05, -0.0002593535, 0.002164789, 
    0.1272842,
  0.228955, 0.02120834, 0.0003083922, 6.735146e-08, 1.635802e-07, 
    5.815604e-09, 0.001280078, 0.01511121, 0.01790782, 0.0005442834, 
    0.008165067, 0.00202413, 0.02069737, 1.651013e-06, 2.625686e-05, 
    0.0009009737, 0.001191365, 0.04657453, 0.04438028, 0.1029545, 0.1845701, 
    0.1624531, 0.009485417, 0.01371715, 0.005526222, 0.00788918, 0.02971238, 
    0.00171874, 0.03448775,
  -3.814813e-05, 0.01930882, 0.03188302, 0.004983678, 0.002564934, 
    0.000958332, 0.003807728, -1.32427e-06, 3.303908e-07, 0.01663668, 
    0.01029594, 0.03233129, 0.07541401, 0.04650757, 0.02353877, 0.01329888, 
    0.03743554, 0.0384206, 0.1024614, 0.04646371, 0.05059883, 0.06610082, 
    0.04515018, 0.04050364, 0.1150893, 0.1479816, 0.1486606, 0.01094606, 
    0.0006181282,
  0.01708651, 0.01076601, 0.0006577059, 0.004352324, -0.0001181879, 
    -6.429629e-06, 0.0001179631, 0, 0, 0, 0, 0, 0.009373583, 0.02753236, 
    0.02829051, 0.01023355, 0.02940908, 0.08019105, 0.06105405, 0.02769545, 
    0.004147334, 0.0006272719, 0.002045106, 0.01617014, 0.04545766, 
    0.09354989, 0.09259813, 0.05224806, 0.03173266,
  0.005974905, 0.0001908998, 0, 0, -1.702003e-06, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0006829477, -4.531837e-05, 0.006960634, 0.01176567, 0.01690797, 
    0.01075986, 0.001248194, -0.0001582129, 0, -2.370933e-05, 0, 0.009401907, 
    0.03551312, 0.03857388, 0.02893593, 0.02669678,
  -0.000105231, -8.147629e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.001521613, 7.366179e-05, -0.0001281482, -2.235308e-05, 0, 0, 0, 
    0.001535818, 0.01348621, 0.003622024, 0.006847163, -5.59153e-05,
  -5.420765e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.01542759, 0.001379554,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -7.38772e-05, -6.87471e-05, 
    0.0001291277, -9.820765e-11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.02420489, 0.02205963, 0.01413839, 0.003351572, -4.029742e-07, 
    -7.078633e-07, 0.01010538, 0.0005204577, -0.000136477, 0, 0, 0, 
    -0.0002523385, 0.002937234, 0.01140039, 0.02384759, 0.03021977, 
    0.01961497, 0.02266525, 0.01294738, 2.592584e-05, -3.277417e-10, 0, 0, 0, 
    -1.004777e-05, 0.00049498, 0.00882639, 0.01065341,
  0.02261878, 0.04289868, 0.0405122, 0.01084832, 0.02143286, 0.02671579, 
    0.03288676, 0.05756041, 0.02879596, 0.02772403, 0.01166599, 0.004817916, 
    0.01605931, 0.02774661, 0.04615238, 0.06619241, 0.04958751, 0.04175945, 
    0.06299102, 0.0489105, 0.01759056, 0.01565795, 0.006884498, 0.02338806, 
    0.01407415, 0.00793215, 0.0349988, 0.02701994, 0.03159292,
  0.08403455, 0.09398653, 0.07988276, 0.1273202, 0.161471, 0.1455221, 
    0.1014405, 0.0948506, 0.08424044, 0.05104613, 0.06659738, 0.06055342, 
    0.0793845, 0.1675685, 0.1713935, 0.08110797, 0.09531575, 0.1604101, 
    0.1344132, 0.09532845, 0.125721, 0.1335927, 0.07593387, 0.06075835, 
    0.08922734, 0.1242857, 0.1226503, 0.1143967, 0.09888644,
  0.03241577, 0.04349153, 0.02109675, 0.07628263, 0.1179873, 0.1380262, 
    0.09482055, 0.0521638, 0.04837326, 0.04690181, 0.06714424, 0.1386289, 
    0.1263411, 0.1534445, 0.05122915, 0.05626451, 0.117598, 0.1196349, 
    0.1179436, 0.1583357, 0.124273, 0.05652944, 0.05268147, 0.008715215, 
    0.06639417, 0.1658091, 0.1118308, 0.1463609, 0.04394746,
  1.255662e-06, -1.318306e-08, 0.1605301, 0.09903442, 0.1240907, 0.06032201, 
    0.09302855, 0.01697458, 0.006434306, 0.07639706, 0.1103725, 0.03352724, 
    0.09947179, 0.1376313, 0.07698514, 0.0253236, 0.149037, 0.1613358, 
    0.1141701, 0.2012988, 0.02500732, 0.022421, 5.527021e-06, 7.763154e-05, 
    0.06782164, 0.1507486, 0.1598467, 0.01578702, 0.003903297,
  1.44188e-05, 0.05154026, 0.1372469, 0.05527909, 0.073066, 0.0548496, 
    0.08533784, 8.334484e-05, 0.000347188, 0.08350784, 0.09232476, 0.1325203, 
    0.2091095, 0.1660818, 0.01564933, 0.1424974, 0.1897065, 0.1315029, 
    0.1444308, 0.0361458, 0.05541091, 1.079018e-09, 0.001358628, 0.1184349, 
    0.2053278, 0.2303236, 0.07041454, 0.03401245, 3.677362e-05,
  0.0001497591, 0.03304183, 0.3806709, 0.1433882, 0.08604794, 0.1377723, 
    0.1347101, 0.07184746, 0.05739762, 0.02294269, 0.04933198, 0.05434924, 
    0.06000912, 0.03929692, 0.08090598, 0.1323695, 0.09883947, 0.0305997, 
    0.001350695, 0.0004300969, 9.71484e-09, 8.657221e-09, 0.005945884, 
    0.4146424, 0.4313499, 0.2267962, 0.1209297, 0.008402631, 1.911076e-06,
  0.001770592, 0.004802009, 0.005301932, 0.0187369, 0.06048233, 0.03211094, 
    0.2207762, 0.05224242, 0.07931406, 0.2321759, 0.0091912, 0.03800701, 
    0.09278404, 0.07562, 0.1253437, 0.0500877, 0.0007141253, 1.378613e-05, 
    0.01586355, 5.944907e-05, 0.0004010306, 0.0006296959, 0.0006868067, 
    0.1616171, 0.1663566, 0.1188785, 0.0189972, 0.0268661, 0.003840063,
  0.001679644, 9.614823e-06, 6.633815e-06, 2.149432e-06, 1.058608e-06, 
    0.004443137, 0.007924726, 0.05650957, 0.002306294, 0.07955206, 
    0.06271288, 0.06500138, 0.1333274, 0.04867042, 0.00343262, 0.002143635, 
    0.01361062, 0.03782644, 0.02459808, 0.06471639, 0.08549594, 0.02698899, 
    0.0002272441, 0.01072706, 0.001153074, 1.292299e-06, -0.0004258325, 
    0.004868966, 0.1339405,
  0.2117812, 0.007912654, 0.0081346, 2.880805e-06, 1.20209e-07, 0, 
    0.007489387, 0.01802968, 0.03608442, 0.007861828, 0.009144921, 
    0.003387561, 0.02090056, 2.761162e-05, -9.629297e-06, 0.003783795, 
    0.001249392, 0.04631824, 0.05678723, 0.1235041, 0.1760733, 0.1133481, 
    0.001816103, 0.0186842, 0.002999375, 0.007747864, 0.04883087, 0.01309819, 
    0.05370496,
  0.01459246, 0.09070139, 0.0374978, 0.06603032, 0.02232642, 0.03325787, 
    0.08055352, -0.0003173148, 1.379504e-05, 0.04083763, 0.02164151, 
    0.035275, 0.1140389, 0.06008888, 0.06335795, 0.06052001, 0.114322, 
    0.1765045, 0.2422671, 0.1180859, 0.0339449, 0.0695031, 0.07243405, 
    0.06330568, 0.1739704, 0.1973781, 0.2082411, 0.04248746, 0.01583513,
  0.04471761, 0.03240261, 0.01295311, 0.01028735, 0.0001036738, 0.0003561566, 
    0.001536185, 0, 0, 0, 0, 2.973424e-05, 0.01822514, 0.04284225, 
    0.06882556, 0.0379022, 0.05125273, 0.1342749, 0.1019236, 0.05506808, 
    0.01133109, 0.008498305, 0.02344271, 0.04714873, 0.09065592, 0.1644014, 
    0.1591721, 0.143222, 0.07845775,
  0.0177959, 0.0008795843, 0.0001232512, -1.448415e-05, -1.133308e-06, 0, 0, 
    0, 0, 0, 0, 0, -2.300509e-06, 0.01982809, 0.00040787, 0.008547424, 
    0.01646825, 0.03786495, 0.05759637, 0.004191731, 0.0007889209, 
    -0.0001801229, 0.0001948782, 0, 0.01832805, 0.0686914, 0.07728842, 
    0.05261735, 0.04467965,
  0.001106022, 0.000122997, -0.0001291446, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -1.803541e-05, 7.212504e-06, 0, 0.004969968, 0.003458839, 0.006137066, 
    0.002935911, 0, 0, 0, 0.004008568, 0.03136522, 0.02331509, 0.01447878, 
    0.01038177,
  0.00131713, 0.001652403, -1.409181e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.00020727, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.408264e-05, 0.0001797954, 
    -2.11145e-06, 0.01929983, 0.002791352,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9.893284e-06, -0.0008022294, 
    0.004486058, 0.00790402, 0.00646332, 0.0004116306, 0, 0, 0, 0, 0, 0, 
    -0.0001169236, -1.328349e-05, 0, 0,
  0.06783874, 0.05156364, 0.01319059, 0.01736706, -0.0001606598, 
    -0.002592329, 0.03962559, 0.002592367, -0.000298125, -0.0001346915, 
    -1.669683e-08, 0, 0.001507688, 0.0425198, 0.04853063, 0.04829288, 
    0.03118038, 0.05473615, 0.02764739, 0.03047685, 0.02816738, 0.01249038, 
    2.791309e-06, -2.017418e-06, -1.00557e-09, 3.579041e-05, 0.01090809, 
    0.03192684, 0.07397,
  0.06660354, 0.1054237, 0.06691085, 0.04482209, 0.04001807, 0.05415886, 
    0.09480424, 0.08428376, 0.04188687, 0.08950553, 0.06559891, 0.04296569, 
    0.06540508, 0.04745612, 0.07544216, 0.1279609, 0.1085888, 0.1060444, 
    0.1074021, 0.08012439, 0.07016232, 0.08548819, 0.06852379, 0.07324778, 
    0.04847921, 0.0919507, 0.07808353, 0.07145167, 0.06940727,
  0.12318, 0.1231961, 0.1455428, 0.1662791, 0.1768364, 0.1657843, 0.108855, 
    0.1280814, 0.1431097, 0.1006885, 0.1378523, 0.1036598, 0.1168384, 
    0.201904, 0.1755327, 0.0925006, 0.09116043, 0.1507045, 0.1226008, 
    0.1190038, 0.1449646, 0.1758237, 0.1614551, 0.1120202, 0.1506885, 
    0.1517316, 0.1589171, 0.1277966, 0.1284734,
  0.03187616, 0.03945896, 0.02509984, 0.06824639, 0.1052735, 0.1251406, 
    0.08683259, 0.05770458, 0.04223676, 0.04023366, 0.06755945, 0.1167633, 
    0.1059241, 0.116965, 0.03958568, 0.04049106, 0.09501999, 0.106445, 
    0.09537897, 0.1496707, 0.1127935, 0.04396001, 0.04969358, 0.01104416, 
    0.06186041, 0.1288191, 0.09665117, 0.1322608, 0.04511369,
  2.184967e-06, 1.729007e-07, 0.1483624, 0.07955361, 0.1368131, 0.06159436, 
    0.08351142, 0.01351512, 0.007415411, 0.07706925, 0.1114503, 0.03086378, 
    0.09916107, 0.1265229, 0.06013138, 0.01644552, 0.1327593, 0.1448191, 
    0.08542625, 0.2158841, 0.02949736, 0.0145028, 4.151332e-07, 
    -5.297867e-06, 0.05262876, 0.1439202, 0.1343466, 0.01281511, 0.000296114,
  2.808152e-06, 0.04812712, 0.1207189, 0.03792662, 0.06388218, 0.0381469, 
    0.08036011, 0.001214586, 0.0003007245, 0.07032564, 0.08653022, 
    0.09775869, 0.1909077, 0.126449, 0.01117537, 0.1273536, 0.1650085, 
    0.1225638, 0.1191843, 0.02223814, 0.02719164, -2.150055e-09, 0.01603245, 
    0.1017969, 0.1457191, 0.2443231, 0.06069428, 0.01599528, 2.574639e-06,
  2.226707e-05, 0.02573087, 0.3376652, 0.1094412, 0.07116976, 0.1012674, 
    0.123412, 0.05273095, 0.04384632, 0.01578611, 0.03285172, 0.05122731, 
    0.04245306, 0.03679679, 0.05689027, 0.1249536, 0.0831144, 0.03088068, 
    0.001103563, 5.384186e-06, -3.82466e-10, 1.123986e-07, 0.002327767, 
    0.3509074, 0.3916523, 0.1916142, 0.08292927, 0.002700758, 1.544449e-07,
  0.001401512, 0.009127505, 0.004515599, 0.004445807, 0.0591195, 0.02177233, 
    0.2086146, 0.0555006, 0.06041669, 0.1879133, 0.007033889, 0.03180097, 
    0.08581632, 0.06070245, 0.1103831, 0.04491255, 0.0006063314, 2.85975e-06, 
    0.007989473, 6.027689e-05, 0.004601391, -3.570581e-05, 0.0004110935, 
    0.0995264, 0.1260237, 0.1671625, 0.02017166, 0.02850299, 0.0001795885,
  7.858464e-05, 7.746468e-06, 2.037082e-06, 6.685274e-07, 1.527541e-06, 
    0.0005999933, 0.002620631, 0.06008932, 0.003751217, 0.06623248, 
    0.06436098, 0.0674202, 0.1178093, 0.04521747, 0.01296982, 0.001399052, 
    0.01535853, 0.03591232, 0.0288227, 0.06202899, 0.07280544, 0.02916609, 
    0.0003956749, 0.00412266, 0.0009377236, 1.819015e-07, 0.002530685, 
    0.0004544801, 0.1008439,
  0.1575584, 0.002843733, 0.0008368188, -4.226333e-07, 3.549101e-08, 0, 
    0.01849577, 0.02030777, 0.0595511, 0.008517009, 0.03639557, 0.01578193, 
    0.02294227, 0.002590511, -1.321466e-05, 9.509311e-05, 0.00078831, 
    0.05158991, 0.02870639, 0.1119935, 0.167148, 0.07391917, 0.0004309175, 
    0.0182463, 0.00831664, 0.004622436, 0.01575143, 0.02225661, 0.02997632,
  0.04096216, 0.07951738, 0.02937796, 0.03932369, 0.03616417, 0.0299755, 
    0.06730484, -0.000205172, 0.001182565, 0.05451606, 0.02655236, 
    0.03066062, 0.1327164, 0.08611132, 0.08879737, 0.08552159, 0.1270356, 
    0.185985, 0.2176432, 0.06783242, 0.02086389, 0.0668626, 0.03505445, 
    0.05852659, 0.1822202, 0.1956259, 0.1747139, 0.04302372, 0.04085006,
  0.09318119, 0.07279369, 0.06861106, 0.03368138, 0.01198087, 0.03871924, 
    0.002838254, 0.0004704174, 4.111493e-05, -8.60785e-10, 0, 0.0002501297, 
    0.03637302, 0.08124665, 0.1053157, 0.08298532, 0.1312245, 0.191535, 
    0.2079102, 0.1382584, 0.02088691, 0.04673568, 0.07825758, 0.1318817, 
    0.1549593, 0.2215153, 0.1864581, 0.1517099, 0.1530058,
  0.1185329, 0.05199175, 0.01703347, 0.007245821, 0.003748826, 0.001500549, 
    -4.838457e-06, 0, 0, 0, 0, 0, 0.001561517, 0.04728576, 0.01541158, 
    0.01807978, 0.03270311, 0.07504401, 0.09549496, 0.01303544, 0.00728212, 
    0.0143624, 0.007344335, -7.797888e-05, 0.04217207, 0.1070011, 0.1741962, 
    0.1576986, 0.1391322,
  0.05325194, 0.003371517, 0.0002039258, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.001047128, 0.005383277, 8.298047e-05, 0.0004833082, 0.0154397, 
    0.01560822, 0.01641091, 0.01301005, 0.0001486036, 0.0002394623, 
    0.0005348247, 0.006414944, 0.03783454, 0.0680419, 0.05992846, 0.04734464,
  0.0173113, 0.01289196, 0.002485129, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0002815416, -1.748529e-05, 0, 0, -4.735029e-05, 0, -2.061117e-05, 
    -1.068049e-05, -1.027113e-07, 0, 0.003306908, 0.004392277, -7.58029e-06, 
    0.02467484, 0.009384834,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001099813, 0.01445424, 0.01259656, 
    0.01062122, 0.01198137, 0.001901611, -4.585177e-06, -1.735027e-07, 
    -2.584241e-10, 0.0002966651, 0.007690875, 0.002754468, -0.00140737, 
    -0.0007232754, -0.0001027644, 0,
  0.07248737, 0.05136804, 0.01436824, 0.01555286, -0.0006362204, 0.01562331, 
    0.123424, 0.007269188, 0.003130623, -0.002481364, -9.894286e-06, 0, 
    0.01817732, 0.2075983, 0.1861272, 0.1213805, 0.1148305, 0.08107008, 
    0.05363712, 0.07194125, 0.06431992, 0.07168062, 0.06203262, 0.05965451, 
    0.08316776, 0.08704982, 0.02821475, 0.04650831, 0.08907621,
  0.1024832, 0.1466394, 0.1131817, 0.1115692, 0.1078449, 0.1190098, 
    0.1248832, 0.1312931, 0.04712952, 0.1725349, 0.1550831, 0.1288474, 
    0.1331611, 0.127436, 0.1053908, 0.2234028, 0.1378991, 0.1212733, 
    0.1121776, 0.09165332, 0.1206781, 0.1388669, 0.1920724, 0.1786861, 
    0.1662033, 0.2105012, 0.1725009, 0.1210395, 0.09741882,
  0.130261, 0.1489922, 0.1522757, 0.1903692, 0.1676403, 0.1656184, 0.1150208, 
    0.1454459, 0.1718854, 0.1179971, 0.1473399, 0.09286627, 0.0979191, 
    0.2129962, 0.1832237, 0.1240129, 0.09807997, 0.1398961, 0.1191628, 
    0.1097314, 0.1450017, 0.1918431, 0.1956896, 0.1359617, 0.1693544, 
    0.1701193, 0.1646755, 0.120857, 0.1453046,
  0.03158873, 0.03712245, 0.02565469, 0.06362619, 0.1028732, 0.1143756, 
    0.06400726, 0.04872185, 0.03073057, 0.03915324, 0.05004953, 0.1052576, 
    0.09482057, 0.1052427, 0.03068126, 0.03671233, 0.08109424, 0.09525473, 
    0.0754142, 0.1566918, 0.09395681, 0.0197745, 0.0247422, 0.008240219, 
    0.05991143, 0.1075012, 0.09332779, 0.1178403, 0.05241681,
  3.253199e-07, 1.545491e-09, 0.1223705, 0.07292605, 0.1316094, 0.04806081, 
    0.04592186, 0.009541579, 0.005823263, 0.06193326, 0.1138799, 0.0280152, 
    0.09468329, 0.102835, 0.05077467, 0.01040494, 0.1248914, 0.1399028, 
    0.08505755, 0.2262477, 0.0348432, 0.00277966, 3.638197e-08, 
    -6.453306e-06, 0.04394433, 0.1329888, 0.1210281, 0.01508946, 7.518342e-06,
  2.894153e-05, 0.04350193, 0.1211869, 0.03104757, 0.04900818, 0.02618057, 
    0.07930421, 0.003960156, 0.0001754675, 0.06101424, 0.0709266, 0.06212457, 
    0.1508229, 0.09148244, 0.009701177, 0.1195351, 0.1471767, 0.1096791, 
    0.09436476, 0.01172788, 0.003429303, -5.610123e-10, 0.01711984, 
    0.08200579, 0.1059538, 0.2185681, 0.04268573, 0.004472091, 1.147554e-06,
  6.384506e-06, 0.02481422, 0.2868088, 0.07590504, 0.05138726, 0.07164732, 
    0.1137685, 0.03729642, 0.03259282, 0.01266899, 0.02642588, 0.04201763, 
    0.03241858, 0.03284487, 0.03994516, 0.1132048, 0.07116508, 0.03131652, 
    0.0007440256, 8.746864e-07, -1.370042e-09, 1.429625e-07, 0.00188188, 
    0.2509793, 0.3589396, 0.145673, 0.0663665, 0.0007341441, 6.103888e-07,
  0.0008185209, 0.01317026, 0.004595545, 0.001979219, 0.04697962, 0.01596344, 
    0.1835987, 0.05859696, 0.05534884, 0.1569781, 0.005592797, 0.01560071, 
    0.07177354, 0.04941939, 0.08606442, 0.04282632, 0.0005057952, 
    -3.573315e-06, 0.0006721117, -1.816753e-05, 0.009436744, 0.0009541304, 
    0.0003493481, 0.05550541, 0.1256609, 0.1894213, 0.01530571, 0.02218435, 
    0.0002526358,
  1.494666e-05, 5.623043e-06, 8.588052e-07, 2.953922e-07, 1.383068e-06, 
    4.439146e-05, 0.005558326, 0.063692, 0.006550821, 0.0642002, 0.06993017, 
    0.081084, 0.1060524, 0.04126643, 0.009995863, 0.001168372, 0.01710781, 
    0.03815198, 0.03881002, 0.07470154, 0.06429198, 0.03211977, 0.0003564006, 
    0.001768097, 0.0008446287, 5.735175e-09, 0.007664109, 0.0002837702, 
    0.07461844,
  0.1043828, 0.0002778748, 6.022807e-05, -6.162446e-07, 4.274692e-09, 0, 
    0.02330017, 0.02048817, 0.07052886, 0.009365655, 0.07525111, 0.01834124, 
    0.02809067, 0.01695912, -9.717331e-05, -7.136539e-05, 0.002025203, 
    0.03779683, 0.02218709, 0.1126827, 0.1553165, 0.05535538, -4.987307e-05, 
    0.01523887, 0.003118954, 0.006282682, 0.007678187, 0.008079418, 0.01524445,
  0.03141628, 0.06383744, 0.04138937, 0.02787019, 0.0398622, 0.01073376, 
    0.0244052, 0.006530529, 0.009945821, 0.07218536, 0.03069145, 0.03658202, 
    0.1254905, 0.1028572, 0.09916374, 0.09890448, 0.1321511, 0.169221, 
    0.1874238, 0.03173798, 0.01993176, 0.06784227, 0.02727555, 0.04997112, 
    0.1782434, 0.1618815, 0.1181115, 0.03272432, 0.03939759,
  0.1208791, 0.1256378, 0.1443506, 0.08337086, 0.08727093, 0.1399065, 
    0.009085535, 0.04795751, 0.005903808, 1.750511e-05, 0.002302769, 
    0.01446764, 0.0599779, 0.09938206, 0.1330346, 0.1201124, 0.1935341, 
    0.2356919, 0.2306647, 0.235886, 0.0755351, 0.1041845, 0.1181593, 
    0.1297854, 0.1582365, 0.222761, 0.172239, 0.1167198, 0.1510904,
  0.18189, 0.1346746, 0.0807019, 0.08674503, 0.1084284, 0.09570998, 
    0.03446709, 0, -8.036515e-06, 0, 0, -2.16364e-09, 0.009283504, 
    0.07639845, 0.09381574, 0.04821621, 0.07087172, 0.1083544, 0.1672901, 
    0.04016086, 0.05090078, 0.07316324, 0.06366856, 0.02884008, 0.1176855, 
    0.1408294, 0.2022751, 0.2017446, 0.1928671,
  0.1028849, 0.06537935, 0.05323029, 0.01822644, -0.0003932117, 
    -1.692311e-05, 0.0003200885, 0, -0.0001213028, 0, 0, -8.679042e-08, 
    1.556587e-05, 0.05227868, 0.08732657, 0.05056315, 0.01246555, 0.06220113, 
    0.03708898, 0.05347804, 0.04273333, 0.02412507, 0.01321315, 0.03281754, 
    0.01267313, 0.04552528, 0.1371441, 0.1111576, 0.09177892,
  0.02784508, 0.03235491, 0.008051478, 0.0002604694, 0, 0, 0, 0, 0, 0, 0, 0, 
    -2.242412e-06, 0.003558525, 0.0223376, 0.01114349, -0.0001379554, 
    0.00114606, 0.003538645, 0.01701327, 0.02188704, 0.01462906, 0.008853889, 
    -0.000100286, 0.007073448, 0.007312764, -2.716394e-05, 0.03334449, 
    0.0138381,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.005050962, 0.01949537, 0.1197028, 
    0.1403229, 0.1009496, 0.02856351, 0.003399282, -0.0002509237, 
    -4.27968e-05, 0.0119129, 0.08657409, 0.06169285, 0.02224217, 0.03452748, 
    -0.0001122096, 0,
  0.1526136, 0.1517061, 0.08777229, 0.07909704, 0.0005056785, 0.05016379, 
    0.1488395, 0.02592694, 0.01816648, -0.00411931, -2.824797e-05, 
    -0.0004299633, 0.05635857, 0.3425734, 0.2551396, 0.2123336, 0.1596693, 
    0.1449056, 0.1255568, 0.1153652, 0.1115332, 0.1350249, 0.1793191, 
    0.1326883, 0.1643908, 0.1615259, 0.09542673, 0.1010389, 0.1976952,
  0.1510537, 0.2033711, 0.2106063, 0.1880565, 0.1643556, 0.1593395, 
    0.1338924, 0.1655967, 0.1479933, 0.2255113, 0.2156648, 0.2047288, 
    0.2309158, 0.1786928, 0.1232255, 0.2354384, 0.1802897, 0.1464992, 
    0.1248332, 0.1019706, 0.1687623, 0.2011804, 0.234494, 0.2097116, 
    0.2270362, 0.2511401, 0.2163953, 0.1754124, 0.166946,
  0.1431438, 0.1503208, 0.1437609, 0.188081, 0.1443507, 0.1633409, 0.127745, 
    0.1593623, 0.1968198, 0.1303471, 0.1456861, 0.08304837, 0.09106652, 
    0.20161, 0.1697354, 0.1150781, 0.1147956, 0.1407181, 0.09568056, 
    0.1043455, 0.1488001, 0.2002672, 0.224211, 0.1598766, 0.1588051, 
    0.1707171, 0.1547097, 0.1186948, 0.1426461,
  0.02887273, 0.03325192, 0.02606673, 0.0599153, 0.09469768, 0.09429917, 
    0.06698097, 0.04452645, 0.02235856, 0.04234326, 0.03798127, 0.08370123, 
    0.09108402, 0.09769314, 0.02593311, 0.03468214, 0.07637832, 0.08488797, 
    0.06779481, 0.1598949, 0.1225296, 0.01537135, 0.01456212, 0.007733481, 
    0.0545627, 0.08299555, 0.0908458, 0.1153699, 0.05218782,
  1.435593e-07, -1.246045e-08, 0.1084211, 0.05911712, 0.1023924, 0.03854237, 
    0.01604586, 0.002879271, 0.000142933, 0.0604561, 0.09499586, 0.02660158, 
    0.07886506, 0.07141977, 0.03882379, 0.01041245, 0.1172825, 0.1352065, 
    0.07715789, 0.2042813, 0.02641833, 0.0001101051, -7.297853e-10, 
    -5.217185e-06, 0.03969736, 0.1078308, 0.0978557, 0.0128893, 3.570969e-06,
  0.0007327988, 0.04299333, 0.1157384, 0.02905998, 0.04015746, 0.01799858, 
    0.06678224, 0.001341909, 0.0001947202, 0.07135325, 0.06219363, 
    0.04320408, 0.1140428, 0.06053865, 0.00645697, 0.09934297, 0.1438684, 
    0.09052087, 0.07188874, 0.006075489, 4.084209e-05, 0, 0.0153164, 
    0.06944234, 0.09155373, 0.1812246, 0.04652602, 0.0002862456, 0.0001963398,
  6.648257e-05, 0.01977646, 0.2683746, 0.0559434, 0.04546158, 0.05748262, 
    0.1006161, 0.02760664, 0.02719112, 0.01083023, 0.02168193, 0.03616774, 
    0.02601996, 0.02857271, 0.03601377, 0.1074835, 0.05723474, 0.03016635, 
    0.0007230752, 3.621912e-09, -2.976814e-10, 8.67178e-08, 0.0005184573, 
    0.1723049, 0.330457, 0.1315012, 0.06207963, 6.913655e-06, 1.422992e-06,
  0.005475344, 0.008846999, 0.004196061, 0.004352945, 0.04553221, 0.01183541, 
    0.1703422, 0.06851845, 0.0558017, 0.1295496, 0.004716547, 0.01030937, 
    0.05744482, 0.04099147, 0.07110017, 0.02922962, 0.001790095, 
    -1.180321e-05, -5.20706e-05, -4.422696e-05, 0.01289841, 0.001436026, 
    0.0006917354, 0.0272264, 0.1356466, 0.1899631, 0.01219793, 0.005787367, 
    0.0003417208,
  0.001356761, 3.455922e-06, 1.744077e-07, 8.903756e-07, 4.204597e-06, 
    -4.672729e-05, 0.01298588, 0.06813919, 0.004000566, 0.05933524, 
    0.0851507, 0.09578261, 0.09674276, 0.03384699, 0.007450025, 0.0008156045, 
    0.02047024, 0.04172399, 0.03026988, 0.07881235, 0.05623311, 0.03531357, 
    0.0003045663, 0.001191329, 0.001212591, 3.53164e-07, 0.02139368, 
    0.0008686686, 0.03014879,
  0.06792368, 2.558972e-05, 5.859701e-07, 1.651546e-05, -4.383323e-09, 
    -5.438428e-12, 0.03144702, 0.02129795, 0.0614513, 0.006652822, 
    0.08725926, 0.0377054, 0.0343128, 0.04004623, 0.005883718, 3.490575e-05, 
    0.005087804, 0.03107491, 0.00646169, 0.09482249, 0.1318637, 0.04982965, 
    0.0007190704, 0.01084573, 0.001028746, 0.0002930143, 0.00677592, 
    0.004376783, 0.009201162,
  0.01944811, 0.046073, 0.05224745, 0.02302139, 0.03562328, 0.00289518, 
    0.02774388, 0.01374914, 0.02992326, 0.08697242, 0.02832476, 0.04887203, 
    0.1043062, 0.1402687, 0.1386123, 0.09688902, 0.1245325, 0.1224275, 
    0.122745, 0.01318948, 0.0336929, 0.06325421, 0.04042932, 0.04789636, 
    0.1484471, 0.1298553, 0.1195959, 0.03876976, 0.03253172,
  0.1367248, 0.1436927, 0.2102242, 0.1638287, 0.1037379, 0.2258112, 
    0.04261816, 0.1008402, 0.03409506, 0.008411117, 0.01721843, 0.07459203, 
    0.08718101, 0.1310284, 0.1693335, 0.1639708, 0.2100389, 0.2496425, 
    0.2276031, 0.2244951, 0.1608415, 0.09159178, 0.1522702, 0.12866, 
    0.1687305, 0.2154623, 0.1529174, 0.09519034, 0.1525415,
  0.2106347, 0.1531511, 0.1147694, 0.1585324, 0.2229119, 0.2363807, 
    0.1303158, -0.0002398742, 0.0005669031, -0.0002920417, 0.009624463, 
    0.001331999, 0.05285726, 0.1304076, 0.1284279, 0.06236903, 0.0892472, 
    0.1329483, 0.1799207, 0.1230796, 0.09354767, 0.1333686, 0.1429231, 
    0.1088879, 0.1530448, 0.1529089, 0.2240039, 0.2267469, 0.1869733,
  0.1529579, 0.08340224, 0.107031, 0.08224573, 0.02090778, 0.09156495, 
    0.149507, 0.1242975, 0.02822505, 0.00164129, 2.592229e-06, -1.212439e-06, 
    0.003217133, 0.1085572, 0.1538796, 0.09199978, 0.04501791, 0.1247794, 
    0.08711237, 0.09232496, 0.07254543, 0.06179185, 0.05258206, 0.03942391, 
    0.02853801, 0.1402858, 0.220853, 0.2155388, 0.1645039,
  0.02902874, 0.04925116, 0.02471086, 0.01692184, 0.0129214, -3.684175e-07, 
    0, 8.723665e-05, -1.53559e-05, -7.897237e-06, 0.0002501126, 
    -9.773292e-05, 0.02245085, 0.02397555, 0.07004584, 0.06548745, 0.0702026, 
    0.03463543, 0.04669885, 0.07140167, 0.06535073, 0.03656851, 0.03864395, 
    0.008511829, 0.01847595, 0.01098384, -0.0003188165, 0.04437839, 0.01422191,
  -0.0001142998, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7.49361e-08, 7.227175e-08, 0, 0, 0, 0, -3.700158e-08, -3.599411e-05, 
    -0.0001582701,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  -1.903176e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.055668e-05, 0.04607869, 
    0.1370826, 0.2366671, 0.2530869, 0.1585735, 0.1052638, 0.0321125, 
    0.01709527, -0.0002049317, 0.04228267, 0.0971488, 0.08377275, 0.06897844, 
    0.1055911, 0.02981414, 0.001364371,
  0.1944479, 0.2252108, 0.0862438, 0.1474115, 0.009398163, 0.117357, 
    0.1731676, 0.06443431, 0.0959952, 0.01294194, -0.0001553939, 
    -0.002213643, 0.1507723, 0.3767981, 0.3298766, 0.2237698, 0.1275033, 
    0.1622297, 0.1309532, 0.1398931, 0.1445724, 0.1387373, 0.1826707, 
    0.1567717, 0.1621343, 0.1527849, 0.1080384, 0.1035459, 0.2693411,
  0.1645913, 0.2042028, 0.24753, 0.2198319, 0.1603436, 0.1709462, 0.1522488, 
    0.1808209, 0.16854, 0.2405051, 0.2229606, 0.2022378, 0.2414329, 
    0.1899176, 0.1573468, 0.2417516, 0.1784298, 0.1814887, 0.1457879, 
    0.1145953, 0.2095803, 0.2111745, 0.2430593, 0.1989509, 0.2332481, 
    0.2493245, 0.2141547, 0.1907047, 0.2140388,
  0.1451258, 0.1641929, 0.1523867, 0.1886526, 0.1324976, 0.1603602, 
    0.1272981, 0.1584011, 0.2047124, 0.140747, 0.1575416, 0.07589857, 
    0.09236718, 0.1887165, 0.1603348, 0.1000589, 0.1440794, 0.1240104, 
    0.09493785, 0.1195453, 0.1481785, 0.1896785, 0.1939916, 0.157034, 
    0.1464171, 0.1606503, 0.1394342, 0.1160686, 0.1507631,
  0.03218318, 0.03817274, 0.01861818, 0.06729776, 0.07944821, 0.07865333, 
    0.06293181, 0.03723996, 0.02870966, 0.02349606, 0.02015688, 0.06573679, 
    0.09263004, 0.07700575, 0.02380252, 0.02783678, 0.07286604, 0.0815311, 
    0.09109689, 0.1539232, 0.07916907, 0.01532823, 0.01422142, 0.008226475, 
    0.0569852, 0.06934026, 0.08414555, 0.09044829, 0.04989141,
  -5.637626e-07, 1.425767e-08, 0.09797886, 0.05092187, 0.08970978, 
    0.04124327, 0.02364695, 0.001883154, -4.734672e-05, 0.06709255, 
    0.07533195, 0.02639421, 0.07092034, 0.05453961, 0.03338362, 0.01262463, 
    0.08472255, 0.1422033, 0.07010496, 0.1714476, 0.01268424, 3.814484e-06, 
    -4.502756e-12, -2.59027e-05, 0.03893592, 0.08250288, 0.07697897, 
    0.003176299, 5.682381e-06,
  0.003973897, 0.04982936, 0.07845403, 0.02788414, 0.03318271, 0.0145516, 
    0.04802379, 0.0001593388, 0.0001872609, 0.07487684, 0.05388971, 
    0.03235186, 0.101956, 0.05589308, 0.0166712, 0.09506033, 0.1323451, 
    0.07615723, 0.05202926, 0.005406342, 5.577251e-06, 0, 0.0005416474, 
    0.04282045, 0.08433531, 0.1454538, 0.03619719, 1.340438e-05, 0.01670005,
  0.003529181, 0.02589602, 0.2481229, 0.05132698, 0.04295474, 0.04663796, 
    0.07951833, 0.02069402, 0.01745136, 0.0128165, 0.01958584, 0.0295838, 
    0.02130332, 0.02662919, 0.03567334, 0.08850719, 0.0558339, 0.0355593, 
    0.001258208, -2.076487e-08, -9.211675e-10, 3.981756e-08, 0.0001329954, 
    0.1251988, 0.3015924, 0.129624, 0.04167736, 4.199338e-06, 2.510177e-06,
  0.02546419, 0.007615761, 0.005655342, 0.0127449, 0.05938752, 0.00796358, 
    0.1567768, 0.07072879, 0.05311159, 0.1208567, 0.003818813, 0.006879613, 
    0.05194599, 0.03509301, 0.07552846, 0.01881223, 0.001827594, 0.006311337, 
    -2.393094e-05, -1.500134e-05, 0.01198565, 0.002277552, 0.0007747777, 
    0.01746462, 0.1764426, 0.1850805, 0.0133476, 0.003172577, 0.0008951339,
  0.007926437, 7.611438e-06, 3.27947e-07, 1.636951e-06, 5.163201e-06, 
    -2.649386e-05, 0.0370113, 0.06099409, 0.003970795, 0.07903542, 0.1204603, 
    0.1003604, 0.09182949, 0.03657851, 0.01174073, 0.0006883846, 0.0176612, 
    0.04343097, 0.02434514, 0.09568203, 0.05681465, 0.03521837, 0.000295497, 
    0.001038361, 0.001050131, 3.516417e-05, 0.02873384, 0.0007091755, 
    0.01548402,
  0.06645641, 7.892769e-06, 6.773697e-07, 6.137335e-06, 7.97272e-09, 
    1.712401e-09, 0.03113663, 0.02227144, 0.04830227, 0.01817361, 0.109466, 
    0.05998921, 0.04673296, 0.01329531, 0.000413529, -1.375715e-06, 
    0.0001137887, 0.02962616, 0.001055344, 0.07877617, 0.09886818, 0.0442906, 
    0.0007527801, 0.008487444, 0.0002247006, 0.0001107826, 0.009178122, 
    0.004972248, 0.01223475,
  0.01279455, 0.02860395, 0.03614814, 0.0274948, 0.03014347, 0.008339585, 
    0.03684278, 0.03567139, 0.03990546, 0.1014131, 0.02552122, 0.05099196, 
    0.07588753, 0.1440656, 0.1439898, 0.09335088, 0.1246448, 0.1041458, 
    0.09826841, 0.004568723, 0.02527489, 0.05758749, 0.05750397, 0.05153329, 
    0.1201377, 0.1301382, 0.09428947, 0.02875297, 0.02092219,
  0.1546298, 0.1410479, 0.2231086, 0.2128647, 0.1079447, 0.1986471, 
    0.0947448, 0.1316371, 0.05946753, 0.03766324, 0.03468704, 0.1066816, 
    0.111419, 0.140562, 0.174265, 0.2037053, 0.2162852, 0.2376417, 0.21487, 
    0.2097056, 0.1762199, 0.07661913, 0.1492729, 0.1114131, 0.174578, 
    0.1967407, 0.1471404, 0.07920422, 0.1585452,
  0.2061864, 0.2164836, 0.1332319, 0.1919127, 0.236147, 0.2749152, 0.1636023, 
    0.01858062, 0.006378496, 0.03761726, 0.05659078, 0.03582675, 0.08058901, 
    0.2568499, 0.1617362, 0.08103932, 0.1291516, 0.1648086, 0.1675772, 
    0.1533657, 0.1061675, 0.1786176, 0.1770015, 0.1921753, 0.2206734, 
    0.1666487, 0.2080933, 0.2057634, 0.1790718,
  0.1985082, 0.1512466, 0.1408568, 0.1198864, 0.07701552, 0.2511649, 
    0.3083136, 0.2872935, 0.217466, 0.09170378, 0.002809571, -0.0001851682, 
    0.04204453, 0.1522414, 0.1636532, 0.1016641, 0.09784758, 0.2024604, 
    0.1520214, 0.1152827, 0.1087073, 0.09514458, 0.055798, 0.04627994, 
    0.08680756, 0.229136, 0.2741416, 0.2528757, 0.168221,
  0.06163578, 0.08814752, 0.05118975, 0.05094939, 0.03946781, 0.01344404, 
    0.02992753, 0.0504044, 0.02446205, 0.03265555, 0.02034638, 0.03582387, 
    0.07830191, 0.06486776, 0.09235529, 0.07540183, 0.1124613, 0.1521331, 
    0.09553755, 0.1454391, 0.1078195, 0.05389488, 0.05225382, 0.03696382, 
    0.07051624, 0.01542285, -0.0003910362, 0.1049509, 0.06211895,
  0.03208523, 0.02781142, 0.0289249, 0.01096216, 0.001849172, 1.597334e-06, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, -2.872703e-05, 0, 0, -9.439057e-06, 
    8.807526e-05, 0.0001353369, 0.0004463632, -3.037216e-05, -2.160562e-06, 
    -3.973524e-08, 0, -4.59503e-06, -0.006860435, 0.04397248,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0.0121547, 0.008161363, 0.004756056, -9.977946e-05, 0, -0.0001761837, 0, 0, 
    0, 0, 0, 0, 6.066306e-05, 0.172928, 0.2252383, 0.351421, 0.3864838, 
    0.271392, 0.1745332, 0.1358318, 0.0954491, 0.02208991, 0.1291332, 
    0.09792241, 0.08842991, 0.07332444, 0.1164826, 0.1088875, 0.0332562,
  0.1915382, 0.2190218, 0.07534762, 0.1564371, 0.1034314, 0.2432549, 
    0.1814899, 0.1173679, 0.1317339, 0.0361456, 0.00170207, 0.01941195, 
    0.1808928, 0.3814788, 0.3336703, 0.2360748, 0.09351698, 0.1675185, 
    0.1598551, 0.1535057, 0.1479439, 0.0888322, 0.2112697, 0.1567599, 
    0.1710714, 0.1499865, 0.1090599, 0.1128111, 0.2673362,
  0.1668437, 0.1887194, 0.2721481, 0.2241686, 0.1540561, 0.1842724, 
    0.1517847, 0.1909175, 0.2000169, 0.2548541, 0.2387434, 0.2165486, 
    0.2266015, 0.214737, 0.1716975, 0.2370467, 0.1850522, 0.1803463, 
    0.1442348, 0.1506156, 0.2132971, 0.2212973, 0.2485472, 0.2164599, 
    0.2416807, 0.2399734, 0.2128787, 0.1991017, 0.2367083,
  0.1413515, 0.1663871, 0.1701232, 0.1905505, 0.1311613, 0.1666361, 
    0.1589416, 0.1670774, 0.1787123, 0.169271, 0.1542048, 0.07053168, 
    0.1001638, 0.1925712, 0.1697437, 0.1153092, 0.1558653, 0.1244761, 
    0.09273955, 0.1293595, 0.1430645, 0.2140048, 0.2137655, 0.1463823, 
    0.124222, 0.1563523, 0.1304589, 0.121883, 0.1484623,
  0.02541131, 0.04687662, 0.01775182, 0.06541728, 0.08108182, 0.06652089, 
    0.06370823, 0.03225126, 0.02391159, 0.01008668, 0.01832536, 0.06463627, 
    0.09441534, 0.06700306, 0.01999603, 0.02363931, 0.06888884, 0.08342698, 
    0.06629138, 0.1446256, 0.08405894, 0.01311251, 0.02130029, 0.006010946, 
    0.05736154, 0.06096529, 0.07773418, 0.09088551, 0.04779116,
  7.511949e-05, 5.168979e-07, 0.09135064, 0.04700458, 0.06789941, 0.03545142, 
    0.01325841, 0.0004556342, -7.530834e-06, 0.06953038, 0.06423673, 
    0.03201374, 0.06508966, 0.03150392, 0.04211126, 0.0125975, 0.06744365, 
    0.1287462, 0.04025695, 0.1773362, 0.002135112, 1.733033e-07, 0, 
    -1.908865e-05, 0.03490847, 0.06461211, 0.07182579, 0.00140604, 
    1.835157e-06,
  0.01011998, 0.04575177, 0.06469483, 0.02387339, 0.03235061, 0.01937591, 
    0.03358921, -0.0002645126, 0.0001358727, 0.06832153, 0.05407725, 
    0.02405479, 0.08462223, 0.04432142, 0.02079409, 0.1009734, 0.1326113, 
    0.06903892, 0.03840242, 0.006539264, -9.858633e-08, 0, -3.216419e-05, 
    0.01978906, 0.08771958, 0.1421485, 0.0328829, 0.001148993, 0.003985286,
  0.001032124, 0.06205954, 0.2583939, 0.0540652, 0.04890144, 0.04778831, 
    0.06198268, 0.02244697, 0.01262307, 0.01304545, 0.02004991, 0.02745419, 
    0.02471887, 0.02350186, 0.02995077, 0.08023418, 0.04516024, 0.03705786, 
    0.002088633, -1.681286e-08, 8.980439e-10, 1.155572e-07, 5.748116e-05, 
    0.08258442, 0.2803976, 0.1239896, 0.0336021, 1.993996e-05, 7.215858e-07,
  0.08367079, 0.05679219, 0.0138284, 0.02560558, 0.05329303, 0.007180819, 
    0.1455706, 0.06097224, 0.04112598, 0.1334412, 0.002658882, 0.004184659, 
    0.04698977, 0.0315909, 0.0654133, 0.01783001, 0.005921975, 0.009983154, 
    1.278043e-05, -3.019358e-05, 0.01089924, 0.02512512, 0.0008066956, 
    0.02227087, 0.1811446, 0.1746503, 0.01487624, 0.004124795, 0.002903499,
  0.004341155, 8.643346e-06, 1.904598e-07, 9.411563e-07, 1.706243e-06, 
    0.0003163643, 0.03252647, 0.05387868, 0.003202531, 0.06930201, 0.1235941, 
    0.1031002, 0.0771573, 0.03646514, 0.01201622, 0.001787209, 0.01776203, 
    0.04781849, 0.02500791, 0.08001646, 0.06709289, 0.03925177, 0.0002557346, 
    0.001066013, 0.006273127, 0.009882757, 0.03077315, 0.0001920182, 
    0.004591885,
  0.07458857, 1.330653e-05, 2.442819e-06, 2.573124e-06, 6.987729e-08, 
    7.728048e-08, 0.02032993, 0.01628543, 0.03912092, 0.01420293, 0.1057718, 
    0.08793227, 0.03899007, 0.01998458, -9.197515e-05, 6.019762e-06, 
    -7.141757e-05, 0.02772532, -2.034444e-05, 0.03290978, 0.06832745, 
    0.03591812, 0.0004851645, 0.001815251, -5.791565e-05, 9.091479e-05, 
    0.008252622, 0.005447824, 0.02640991,
  0.00520549, 0.01491819, 0.01689384, 0.03058877, 0.02878422, 0.006570073, 
    0.04103151, 0.04262447, 0.04814928, 0.1175094, 0.02602782, 0.04763076, 
    0.05927928, 0.1496565, 0.1281813, 0.08642156, 0.1401882, 0.1004834, 
    0.06727259, 0.004361178, 0.02174117, 0.05122452, 0.06445211, 0.05738768, 
    0.09970792, 0.119492, 0.08190392, 0.03286618, 0.01167523,
  0.1432895, 0.1198243, 0.2410197, 0.2534048, 0.09213973, 0.1679779, 
    0.2196946, 0.1074192, 0.08730496, 0.05859311, 0.04431983, 0.1200922, 
    0.1210709, 0.1420398, 0.1801256, 0.2093401, 0.2241074, 0.2361275, 
    0.1848756, 0.1905323, 0.170215, 0.06679335, 0.1505356, 0.1050508, 
    0.189141, 0.193499, 0.1515909, 0.060327, 0.1611638,
  0.2145505, 0.2374813, 0.1168429, 0.2265907, 0.2467839, 0.2609292, 
    0.1605369, 0.06596141, 0.05632335, 0.09554694, 0.07847619, 0.09106198, 
    0.1354476, 0.3066503, 0.1666386, 0.1052165, 0.1210218, 0.1586487, 
    0.1801232, 0.165265, 0.0945278, 0.1869588, 0.2113149, 0.2684649, 
    0.2262054, 0.1712252, 0.1886761, 0.2037858, 0.1860022,
  0.2322939, 0.1755366, 0.1955438, 0.1667766, 0.1160505, 0.309752, 0.3727993, 
    0.3156587, 0.2624283, 0.1915653, 0.08361954, 0.02900565, 0.09610108, 
    0.1681573, 0.1507571, 0.08395291, 0.1084371, 0.2285409, 0.2259757, 
    0.1092994, 0.1122488, 0.09736505, 0.08658041, 0.05739049, 0.136998, 
    0.253195, 0.2860114, 0.3272705, 0.2004219,
  0.1359365, 0.1107828, 0.1138324, 0.1214375, 0.1495439, 0.07199741, 
    0.1060526, 0.1574611, 0.122472, 0.1200812, 0.08591747, 0.08172613, 
    0.1319962, 0.1366445, 0.1051013, 0.07380981, 0.1273441, 0.2505704, 
    0.1975067, 0.2006631, 0.1786289, 0.1067679, 0.08383452, 0.05608053, 
    0.1167128, 0.01799093, 0.001402184, 0.1538478, 0.1129503,
  0.08448426, 0.1060433, 0.1103472, 0.04719431, 0.02228258, 0.002504176, 
    0.004864368, 0.008148154, 0.0212935, 0.0590229, 0.05678247, 0.03232923, 
    0.007763587, 0.01915436, 0.02406465, 0.01444897, 0.0003191155, 
    -0.0001162326, 9.614741e-05, 0.002069569, 0.01766732, 0.02849055, 
    0.005436833, 0.003526062, -0.0001359049, -1.541798e-05, -0.001041732, 
    0.05224138, 0.1137415,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -4.244298e-05, -4.244298e-05, 
    -4.244298e-05, -4.244298e-05, -4.244298e-05, -4.244298e-05, 
    -4.244298e-05, 0, 0, 0, 0, 0, 0, 0, 0,
  0.06501345, 0.02135089, 0.01394353, 0.004396476, 0.0003128976, 0.001102382, 
    -0.0004104373, -4.154364e-05, -1.385711e-08, 1.105676e-05, -3.885749e-06, 
    -2.047335e-06, 0.002826604, 0.2293585, 0.2305027, 0.3480542, 0.3944682, 
    0.2985877, 0.2207075, 0.202148, 0.1420017, 0.08617679, 0.1826533, 
    0.09161582, 0.09043242, 0.07248589, 0.1263793, 0.1295739, 0.09026657,
  0.2038738, 0.2061066, 0.07190622, 0.1530199, 0.2904222, 0.2912708, 
    0.166031, 0.1508258, 0.1274661, 0.06877178, 0.05552373, 0.07679199, 
    0.1959423, 0.3880225, 0.3493491, 0.2313509, 0.08130327, 0.2004559, 
    0.179031, 0.1616322, 0.1506329, 0.08200588, 0.3055553, 0.1846558, 
    0.1817647, 0.139156, 0.1223748, 0.1291498, 0.2709135,
  0.1718783, 0.1870699, 0.2838381, 0.210589, 0.1528965, 0.2195854, 0.1758773, 
    0.2187367, 0.2211276, 0.2743659, 0.2401702, 0.2334772, 0.2365569, 
    0.2449926, 0.1991747, 0.2201224, 0.1916523, 0.1884918, 0.1550136, 
    0.2050547, 0.2192625, 0.2578377, 0.258817, 0.2152429, 0.2354823, 
    0.2412867, 0.2103788, 0.2170239, 0.2459541,
  0.1399441, 0.1685823, 0.1661148, 0.189484, 0.1428579, 0.1587033, 0.1677811, 
    0.1724559, 0.1808969, 0.1781081, 0.1802961, 0.07466835, 0.1261155, 
    0.2145969, 0.1924015, 0.09999264, 0.1537596, 0.1162349, 0.08190954, 
    0.1417557, 0.1330303, 0.2149086, 0.1955424, 0.1422264, 0.1059184, 
    0.1574354, 0.1292703, 0.1200814, 0.1437224,
  0.03272336, 0.0360025, 0.01734927, 0.06680469, 0.08948362, 0.06158389, 
    0.0601653, 0.03782811, 0.0344721, 0.009495659, 0.02201091, 0.07454814, 
    0.09457522, 0.05526912, 0.0183709, 0.02034975, 0.09293333, 0.08918346, 
    0.0797432, 0.1363005, 0.08230205, 0.01717644, 0.01225576, 0.006097447, 
    0.06227457, 0.05715935, 0.0687267, 0.09438889, 0.04394099,
  0.0003040447, 7.460982e-07, 0.08692424, 0.05843069, 0.06424219, 0.02903178, 
    0.01085154, 0.0002779963, 1.817969e-06, 0.06203337, 0.06496409, 
    0.1041749, 0.07107327, 0.01702476, 0.03952422, 0.01642079, 0.06423892, 
    0.1045782, 0.02469322, 0.1722064, 0.0006676341, 1.317399e-08, 0, 
    0.0001363509, 0.0328977, 0.06271471, 0.08381116, 0.001659995, 8.365395e-07,
  0.002861937, 0.05303438, 0.06981669, 0.02073321, 0.03890284, 0.02644132, 
    0.02469402, -0.000818857, 0.001597096, 0.07653137, 0.0606498, 0.02472991, 
    0.07538597, 0.04630074, 0.02784764, 0.1115957, 0.1281796, 0.07147666, 
    0.02650862, 0.007204829, 1.426822e-08, 6.463718e-10, 1.006371e-05, 
    0.01214482, 0.096404, 0.153687, 0.03431756, 0.01219755, -0.0002505929,
  5.879281e-05, 0.06316858, 0.2739628, 0.05519857, 0.06257065, 0.04883833, 
    0.05656117, 0.02556284, 0.009798536, 0.0198947, 0.02212486, 0.02532414, 
    0.02368683, 0.02010735, 0.02626649, 0.09433174, 0.05205014, 0.03717363, 
    0.003368474, -3.177276e-08, 1.326626e-08, 2.584025e-07, 3.978513e-05, 
    0.07069885, 0.2978967, 0.1081628, 0.02670347, 0.0001047989, 1.646109e-05,
  0.07560529, 0.07418225, 0.03277747, 0.03436115, 0.04634599, 0.00704187, 
    0.1374985, 0.05541994, 0.04210867, 0.1538229, 0.002303377, 0.003388157, 
    0.04704392, 0.03616557, 0.06873484, 0.01732115, 0.008891455, 0.006560268, 
    0.0002060364, 0.0004080184, 0.01064876, 0.04661461, 0.006047443, 
    0.01879325, 0.1672693, 0.1581455, 0.01867754, 0.003381238, 0.02170531,
  -0.0003636097, 6.176894e-06, 3.507139e-07, -1.470534e-06, 9.599985e-06, 
    0.0003534406, 0.03372925, 0.04989995, 0.002243741, 0.07219829, 0.1373424, 
    0.1088281, 0.07006273, 0.03636449, 0.008315837, 0.01068658, 0.0219906, 
    0.05402786, 0.02529664, 0.0698474, 0.06622613, 0.03857896, 0.0003831797, 
    0.001171109, 0.006425676, 0.02384911, 0.008035381, -3.720138e-05, 
    0.007684969,
  0.05242121, -5.343452e-06, 2.008578e-06, 5.985491e-06, 3.018346e-07, 
    6.672651e-06, 0.009629606, 0.006924197, 0.03545184, 0.009090885, 
    0.09699713, 0.0986526, 0.0476563, 0.004721694, -2.483416e-06, 
    2.318751e-06, 0.002099182, 0.01992454, 1.340502e-05, 0.01222214, 
    0.05304892, 0.03059404, 0.02036238, 0.0006914125, 0.0003265886, 
    1.582591e-05, 0.00762952, 0.004264324, 0.03262253,
  0.001313947, 0.009039926, 0.01006074, 0.02280181, 0.0310408, 0.005094095, 
    0.03872767, 0.0449434, 0.0626818, 0.1099215, 0.03616282, 0.04351062, 
    0.04631758, 0.1390733, 0.114096, 0.08798792, 0.1461174, 0.09118491, 
    0.05238479, 0.0001697914, 0.01804943, 0.03633099, 0.06480636, 0.05316343, 
    0.09652878, 0.107651, 0.08180269, 0.04719839, 0.005722851,
  0.1296358, 0.1221175, 0.253843, 0.2612555, 0.08944117, 0.1317739, 
    0.2959383, 0.08533116, 0.07936972, 0.06499805, 0.05208731, 0.1190154, 
    0.1233989, 0.1549652, 0.1925499, 0.1926659, 0.2193825, 0.2149929, 
    0.1622391, 0.1742477, 0.1652862, 0.05587809, 0.1261404, 0.1044169, 
    0.1799206, 0.187226, 0.1406787, 0.05717254, 0.1511434,
  0.2208103, 0.2260567, 0.1269447, 0.2504239, 0.2712602, 0.2574631, 
    0.1547946, 0.1129654, 0.09648361, 0.1143174, 0.0786045, 0.1663398, 
    0.1393268, 0.2961699, 0.1608459, 0.1069338, 0.1221237, 0.1557605, 
    0.1664196, 0.1711432, 0.07984228, 0.2188494, 0.2363994, 0.2833869, 
    0.2425382, 0.1696431, 0.1731695, 0.180188, 0.1653958,
  0.2354116, 0.1986133, 0.2077262, 0.213349, 0.1656673, 0.3643479, 0.3948736, 
    0.3194309, 0.2634299, 0.2255, 0.1362688, 0.08551702, 0.123007, 0.2179118, 
    0.128992, 0.09516995, 0.1218179, 0.2312517, 0.2536319, 0.1073997, 
    0.1200823, 0.09249616, 0.09465051, 0.0672144, 0.1583515, 0.2849524, 
    0.2595688, 0.2740697, 0.1726635,
  0.154313, 0.1537641, 0.1747804, 0.2254578, 0.1774464, 0.1075, 0.2039449, 
    0.2258264, 0.1806646, 0.1929494, 0.1489155, 0.1358971, 0.1565983, 
    0.2003659, 0.1629405, 0.07382127, 0.1677601, 0.2936737, 0.3138196, 
    0.2219849, 0.168288, 0.1164226, 0.1130446, 0.1158636, 0.2294627, 
    0.03178971, 0.01209936, 0.1470373, 0.1008869,
  0.1464132, 0.20459, 0.1801621, 0.0632202, 0.04585875, 0.09898767, 
    0.06795635, 0.07891712, 0.1013774, 0.1036383, 0.0604211, 0.0495805, 
    0.0719739, 0.08503308, 0.0785462, 0.06595027, 0.04892068, 0.00755204, 
    0.0134404, 0.0292705, 0.03787166, 0.05703835, 0.0251621, 0.003922854, 
    0.0008168202, 0.0002935246, -0.009652924, 0.0712994, 0.1669507,
  8.785783e-09, 5.590953e-09, 2.396123e-09, -7.987075e-10, -3.993538e-09, 
    -7.188368e-09, -1.03832e-08, 0, 0, 0, 0, 0, 0, 0, -0.0006453824, 
    -0.0006453824, -0.0006453824, -0.0006453824, -0.0006453824, 
    -0.0006453824, -0.0006453824, -1.983732e-05, -1.983413e-05, 
    -1.983093e-05, -1.982774e-05, -1.982455e-05, -1.982135e-05, 
    -1.981816e-05, 1.134165e-08,
  0.1428165, 0.08510327, 0.02951694, 0.03259527, 0.02488438, 0.01459488, 
    0.01702001, 0.007052139, 0.004062629, 0.0009986293, 3.905739e-07, 
    -0.0002036023, 0.03192737, 0.2219287, 0.2319117, 0.3378726, 0.371248, 
    0.3123928, 0.1919854, 0.2922108, 0.2324097, 0.1678337, 0.1475224, 
    0.07487234, 0.07421789, 0.06464428, 0.1263756, 0.1175122, 0.2015869,
  0.2166261, 0.2063037, 0.06520765, 0.1525394, 0.3456756, 0.3278683, 0.16784, 
    0.1534915, 0.1354467, 0.1345644, 0.1539087, 0.1579499, 0.1915545, 
    0.3880159, 0.3513252, 0.2370692, 0.08612031, 0.2100583, 0.17971, 
    0.1760536, 0.1629108, 0.1114305, 0.3241489, 0.193421, 0.1960552, 
    0.1387337, 0.147415, 0.1446734, 0.2673106,
  0.195173, 0.2120637, 0.297201, 0.2422033, 0.1883111, 0.2688473, 0.232051, 
    0.2624793, 0.2525633, 0.285303, 0.2502697, 0.2359629, 0.2741333, 
    0.2432272, 0.2203488, 0.2192438, 0.1994839, 0.2279528, 0.2023881, 
    0.2105003, 0.2157473, 0.2703944, 0.2469339, 0.1987479, 0.2326568, 
    0.2343606, 0.1949925, 0.2333415, 0.2656083,
  0.1400001, 0.1665258, 0.1850753, 0.196371, 0.1691034, 0.1833896, 0.1808906, 
    0.1725022, 0.1934288, 0.1938023, 0.1820524, 0.09038328, 0.1517501, 
    0.2258327, 0.2208704, 0.116802, 0.154412, 0.1166571, 0.08943778, 
    0.122661, 0.1365853, 0.1959319, 0.2146525, 0.1344034, 0.1042062, 
    0.1680831, 0.1485094, 0.1254242, 0.1593525,
  0.04083007, 0.03181725, 0.01529808, 0.06964255, 0.09610409, 0.05977926, 
    0.0669585, 0.03613136, 0.02848946, 0.008865452, 0.01462382, 0.07451266, 
    0.09078206, 0.04838269, 0.02062436, 0.01861414, 0.05832604, 0.08109241, 
    0.08381841, 0.1329553, 0.06070952, 0.01551033, 0.0120441, 0.01011187, 
    0.06793686, 0.05233936, 0.06746527, 0.07929338, 0.04885508,
  0.0003027459, 1.025748e-05, 0.09410571, 0.07349957, 0.05950195, 0.02986032, 
    0.006438886, 0.0003524968, 1.596173e-06, 0.06978147, 0.06667127, 
    0.07067927, 0.08053165, 0.01065028, 0.03823036, 0.01366577, 0.06455735, 
    0.08729285, 0.02377456, 0.1755851, 0.001660102, 1.096863e-07, 
    2.143941e-12, 0.0005040742, 0.02979474, 0.06748989, 0.09012076, 
    0.002295065, 8.907352e-06,
  4.995487e-05, 0.06574718, 0.07774727, 0.01394311, 0.05311712, 0.03082023, 
    0.02309365, -0.0003797003, 0.009343017, 0.1026261, 0.1003673, 0.03581299, 
    0.08942834, 0.05879775, 0.03892231, 0.1462951, 0.1497814, 0.09395578, 
    0.02565913, 0.008732518, -3.952586e-07, -8.234938e-11, 3.05623e-05, 
    0.008788962, 0.1263451, 0.1618942, 0.03577362, 7.791859e-05, -4.722356e-05,
  0.0001330199, 0.08585954, 0.2909367, 0.08723143, 0.08478174, 0.06061868, 
    0.07090562, 0.03360559, 0.01197328, 0.03458942, 0.03142055, 0.03175876, 
    0.04076998, 0.01925231, 0.03944885, 0.1161851, 0.06352785, 0.03731699, 
    0.004245721, -1.468147e-07, 4.682402e-08, 8.674089e-07, 0.0001271181, 
    0.08047598, 0.3582172, 0.1091193, 0.02752658, 0.0002842635, 0.005874082,
  0.0781853, 0.05985181, 0.02482217, 0.03717026, 0.0403656, 0.01016225, 
    0.1318411, 0.05729916, 0.04868618, 0.1911419, 0.004057181, 0.004023626, 
    0.05164075, 0.04893016, 0.07420254, 0.01999279, 0.009779735, 0.0027488, 
    0.000197976, 0.002046749, 0.01687726, 0.09287202, 0.04329187, 0.03166062, 
    0.168744, 0.1639664, 0.02527141, 0.004112056, 0.03816252,
  -0.0001032334, 1.870523e-06, 7.421656e-07, 9.110511e-05, 1.470745e-06, 
    0.008371343, 0.03458477, 0.05788831, 0.001783859, 0.08546749, 0.1695178, 
    0.1213407, 0.07533976, 0.0433135, 0.005412167, 0.01085117, 0.02001684, 
    0.04412104, 0.0298265, 0.06666104, 0.07330513, 0.0426823, 0.0004673813, 
    0.001642794, 0.005004853, 0.007282684, -0.001310505, -4.431753e-05, 
    0.01995187,
  0.02929164, 1.533935e-06, 3.268999e-06, 3.413721e-05, 9.938583e-07, 
    0.0003051753, 0.0010237, 0.002859267, 0.03019934, 0.002847817, 
    0.09614558, 0.09344777, 0.04631377, 0.0004965581, 1.310319e-06, 
    1.00234e-06, 0.00666552, 0.01198989, 0.0009874309, 0.002271508, 
    0.04396185, 0.02845835, 0.05045336, 0.0008582352, 0.006337036, 
    0.0002239824, 0.00578607, 0.0019372, 0.04960458,
  0.001144066, 0.01568384, 0.01186716, 0.01346308, 0.03163612, 0.01220124, 
    0.03154692, 0.05624146, 0.08728712, 0.1058625, 0.06768702, 0.0500292, 
    0.05228502, 0.1334712, 0.1154645, 0.1135665, 0.1385357, 0.08818453, 
    0.04441152, -0.0002189018, 0.0143705, 0.02559578, 0.06493806, 0.05549339, 
    0.09496595, 0.1020088, 0.07556883, 0.03510936, 0.003727825,
  0.1150618, 0.132468, 0.250885, 0.2733125, 0.0889414, 0.09948932, 0.3325, 
    0.06082463, 0.07221123, 0.05532568, 0.06186703, 0.1155887, 0.1297369, 
    0.153667, 0.1938364, 0.200145, 0.2348726, 0.2066955, 0.1442158, 
    0.1635946, 0.1742481, 0.06007766, 0.1091463, 0.1114611, 0.1716452, 
    0.1659691, 0.1217475, 0.05354012, 0.1421703,
  0.2009059, 0.2228984, 0.1512437, 0.2665146, 0.2733917, 0.2316328, 
    0.1408015, 0.1149952, 0.1047572, 0.1005966, 0.07543814, 0.1953312, 
    0.1385858, 0.2830516, 0.1755471, 0.1030019, 0.09755768, 0.1469355, 
    0.161616, 0.1974771, 0.09875482, 0.2096756, 0.2024347, 0.3167044, 
    0.2434864, 0.1758216, 0.1687748, 0.1613382, 0.1730205,
  0.2107435, 0.2065298, 0.1999392, 0.254462, 0.2061434, 0.3777432, 0.3746559, 
    0.3389176, 0.2709655, 0.2274019, 0.1954193, 0.1172774, 0.1450127, 
    0.2182814, 0.1479549, 0.08663934, 0.142783, 0.2447578, 0.2664014, 
    0.1492744, 0.1334145, 0.1055484, 0.1068488, 0.1648037, 0.1671054, 
    0.2866861, 0.2444972, 0.2782509, 0.19447,
  0.1640449, 0.1586417, 0.2349187, 0.2778383, 0.2056701, 0.1929334, 
    0.2600307, 0.2876602, 0.200583, 0.209256, 0.2234971, 0.1653406, 
    0.1763415, 0.2417264, 0.2307779, 0.1143871, 0.22677, 0.3260788, 
    0.3785014, 0.2493417, 0.1818242, 0.1385238, 0.1182295, 0.1709882, 
    0.2778844, 0.06973193, 0.02729766, 0.1463314, 0.09925795,
  0.2376749, 0.2731006, 0.1976922, 0.1144807, 0.1129464, 0.1631703, 
    0.1647346, 0.1147928, 0.1114799, 0.1404686, 0.1256673, 0.1072913, 
    0.09484121, 0.1043637, 0.1116135, 0.09708848, 0.07111604, 0.06583745, 
    0.03796903, 0.05434741, 0.07457348, 0.1187536, 0.0531978, 0.03455959, 
    0.01399476, 0.001587591, 0.02333897, 0.1222212, 0.252665,
  0.002939393, 0.001987103, 0.001034814, 8.252418e-05, -0.0008697654, 
    -0.001822055, -0.002774345, -0.0002336047, 0.00164181, 0.003517225, 
    0.00539264, 0.007268055, 0.00914347, 0.01101888, 0.01331057, 0.01495553, 
    0.01660049, 0.01824545, 0.01989041, 0.02153537, 0.02318033, 0.007121198, 
    0.004553112, 0.001985026, -0.0005830606, -0.003151147, -0.005719233, 
    -0.008287319, 0.003701225,
  0.2557682, 0.1874608, 0.04252131, 0.03868494, 0.04245775, 0.03206955, 
    0.03012799, 0.02706428, 0.006992012, -5.24867e-05, -0.000590397, 
    0.007165307, 0.07628992, 0.2318533, 0.2513532, 0.3225276, 0.3828876, 
    0.2912799, 0.1730583, 0.314647, 0.2458526, 0.1925691, 0.1170579, 
    0.05701055, 0.06618941, 0.06445267, 0.1355296, 0.1111822, 0.1923922,
  0.2619868, 0.2400159, 0.09450962, 0.1473016, 0.3737861, 0.352385, 
    0.1601638, 0.1587377, 0.1792242, 0.2356036, 0.2857444, 0.1901959, 
    0.1994583, 0.3966737, 0.3305212, 0.2634673, 0.1266306, 0.1996767, 
    0.1537971, 0.176531, 0.1261743, 0.1596268, 0.2694212, 0.1855425, 
    0.2126732, 0.162993, 0.1794632, 0.13539, 0.2906297,
  0.2338101, 0.251722, 0.3056276, 0.325474, 0.2602569, 0.3183883, 0.2595633, 
    0.318667, 0.3127908, 0.3024224, 0.2327152, 0.2579809, 0.2509332, 
    0.1880404, 0.2297535, 0.2056321, 0.2131988, 0.2315501, 0.2219047, 
    0.1955425, 0.2477456, 0.264648, 0.2844574, 0.2657656, 0.2437879, 
    0.2311733, 0.2026251, 0.2449269, 0.2797915,
  0.1572738, 0.1918873, 0.1818475, 0.1954179, 0.1680271, 0.1906196, 
    0.1912493, 0.1843885, 0.2091915, 0.2076716, 0.1902246, 0.10347, 
    0.1756735, 0.2463975, 0.227174, 0.1329403, 0.1333318, 0.1210222, 
    0.09638622, 0.135339, 0.1465723, 0.2174786, 0.2031619, 0.1353329, 
    0.106021, 0.1470772, 0.1400933, 0.1420506, 0.1645939,
  0.04331438, 0.02985012, 0.01625542, 0.07089812, 0.09256153, 0.06032897, 
    0.0741709, 0.04237477, 0.03082267, 0.009950259, 0.01485321, 0.07013105, 
    0.08437167, 0.03891467, 0.02168056, 0.02143398, 0.05215487, 0.08120299, 
    0.09091223, 0.1325689, 0.06299181, 0.02379703, 0.01267072, 0.017092, 
    0.07473302, 0.05548179, 0.0660183, 0.07382692, 0.0521341,
  0.0002926122, 2.032987e-06, 0.1145824, 0.07156668, 0.0524032, 0.02832648, 
    0.005012807, 0.0005290338, -2.474318e-06, 0.08317378, 0.08258116, 
    0.08997179, 0.09128822, 0.009258487, 0.04329699, 0.001365972, 0.07226854, 
    0.103266, 0.02812756, 0.1750729, 0.003501951, 7.460692e-06, 4.411895e-08, 
    0.001237697, 0.02867794, 0.06996197, 0.09964442, 0.004921711, 5.246924e-05,
  1.847991e-05, 0.111965, 0.09596409, 0.01375919, 0.06995224, 0.03877165, 
    0.0268101, -0.0007351874, 0.01184362, 0.1114648, 0.1046139, 0.05430211, 
    0.09286746, 0.05833438, 0.03832558, 0.1664027, 0.1676083, 0.1442689, 
    0.03295098, 0.0151167, 9.526634e-06, 7.614196e-10, 1.980959e-05, 
    0.005072027, 0.1659487, 0.1903642, 0.03269553, 3.651415e-05, -1.148398e-05,
  0.0004708233, 0.04992448, 0.3500978, 0.1332857, 0.07974198, 0.07513612, 
    0.09135966, 0.04292205, 0.01668916, 0.04047307, 0.050483, 0.03817086, 
    0.06992374, 0.0195285, 0.04919377, 0.1471103, 0.06627758, 0.03058068, 
    0.003127997, -4.044456e-07, 6.892084e-08, 5.306894e-07, 0.0001059022, 
    0.1047115, 0.4469329, 0.1420116, 0.024869, 0.0001378558, 0.0007922583,
  0.1138871, 0.05929521, 0.01821693, 0.03329341, 0.03455711, 0.01212303, 
    0.1413, 0.06317664, 0.06606886, 0.2418685, 0.006788903, 0.004069885, 
    0.054408, 0.04813354, 0.08173338, 0.01898387, 0.01002697, 0.0009223594, 
    0.0001554366, 0.001913434, 0.009590381, 0.08805017, 0.0786244, 
    0.04876285, 0.1813864, 0.1676478, 0.02835337, 0.003456748, 0.04529035,
  -1.560852e-06, 1.028259e-05, 7.655725e-07, 0.003129956, -2.048047e-06, 
    0.01454691, 0.03216148, 0.06845709, 0.002455376, 0.08418757, 0.2044842, 
    0.1269164, 0.07951473, 0.05451339, 0.01007336, 0.008526591, 0.02997704, 
    0.04287133, 0.03647788, 0.06241528, 0.07071549, 0.04252798, 0.001265704, 
    0.003333521, 0.008961873, 0.0004527249, -0.0007924556, 0.0008903561, 
    0.01223535,
  0.009336205, 9.624398e-07, 2.308188e-06, 0.0001792411, 1.039511e-06, 
    0.004592853, -0.000100369, 0.004106907, 0.02307216, -0.0002475402, 
    0.1116558, 0.07992177, 0.04928265, 0.00177591, 7.979281e-07, 3.98712e-06, 
    0.01214322, 0.009478132, 0.002477461, 0.001410465, 0.03112166, 
    0.03370755, 0.05577229, 0.00373985, 0.01435658, 0.003586831, 0.003265691, 
    0.0003219362, 0.05179185,
  0.004429348, 0.03565004, 0.01757292, 0.01122432, 0.03668411, 0.01928413, 
    0.02477152, 0.04403765, 0.1125167, 0.1201319, 0.06021302, 0.05161414, 
    0.06005929, 0.138991, 0.1124994, 0.1240967, 0.1279285, 0.08572035, 
    0.04721481, 0.0004883315, 0.0122903, 0.03036485, 0.06564576, 0.05780622, 
    0.09210801, 0.1001757, 0.07273156, 0.02472158, 0.002743419,
  0.1009887, 0.1419174, 0.2419471, 0.2966229, 0.08689732, 0.07680572, 
    0.3419321, 0.03412467, 0.06781582, 0.042421, 0.0704709, 0.1009041, 
    0.1268543, 0.1441168, 0.1988074, 0.2033666, 0.2288365, 0.2071426, 
    0.1409352, 0.1660757, 0.1732522, 0.06458445, 0.09656224, 0.09289519, 
    0.1780648, 0.1524802, 0.1183083, 0.04667727, 0.1340423,
  0.2180285, 0.2267974, 0.122148, 0.2684949, 0.2637524, 0.2128632, 0.1284345, 
    0.1107334, 0.09304952, 0.08316696, 0.06551463, 0.1986999, 0.1312424, 
    0.2849231, 0.1851625, 0.0933103, 0.1053005, 0.1445316, 0.1558229, 
    0.2383535, 0.09365553, 0.1960559, 0.2007063, 0.3461184, 0.2491208, 
    0.1511696, 0.1786059, 0.1525736, 0.1769126,
  0.2069685, 0.1967626, 0.2033238, 0.2977465, 0.2332112, 0.3585589, 
    0.3586076, 0.3294325, 0.2619238, 0.2526036, 0.224554, 0.1640537, 
    0.176511, 0.2106954, 0.1393553, 0.08053803, 0.1283009, 0.2591492, 
    0.2655121, 0.172898, 0.158931, 0.11675, 0.1521793, 0.2143359, 0.1679424, 
    0.2871181, 0.2342026, 0.3152027, 0.1818433,
  0.1678563, 0.1628653, 0.2656201, 0.3204913, 0.3112827, 0.2852093, 
    0.2558533, 0.3271072, 0.2108519, 0.22082, 0.2363145, 0.2130022, 
    0.1968369, 0.2455983, 0.2381188, 0.1216827, 0.24038, 0.3477384, 0.39632, 
    0.3010626, 0.2216727, 0.1573349, 0.1688598, 0.2270614, 0.287601, 
    0.1855094, 0.04851608, 0.149783, 0.131218,
  0.2398305, 0.2874112, 0.2173205, 0.1389242, 0.1677187, 0.1882214, 
    0.2121256, 0.1652737, 0.1702679, 0.1867342, 0.1581023, 0.1393841, 
    0.1225635, 0.1289319, 0.1699747, 0.1836969, 0.1041352, 0.105437, 
    0.1028683, 0.1083314, 0.1417416, 0.1736762, 0.08556206, 0.04606305, 
    0.06326593, 0.004547732, 0.04352751, 0.1942991, 0.2667413,
  0.05468941, 0.05095281, 0.04721621, 0.0434796, 0.039743, 0.0360064, 
    0.0322698, 0.03199148, 0.03867174, 0.045352, 0.05203227, 0.05871253, 
    0.06539279, 0.07207306, 0.07411024, 0.07324464, 0.07237904, 0.07151344, 
    0.07064784, 0.06978225, 0.06891665, 0.0756513, 0.07357323, 0.07149517, 
    0.0694171, 0.06733904, 0.06526098, 0.06318291, 0.05767869,
  0.2539347, 0.2629735, 0.1416347, 0.0474176, 0.0575901, 0.05186553, 
    0.02660149, 0.02352542, 0.01098414, -9.99259e-06, -0.003720328, 
    0.0998875, 0.179478, 0.1949845, 0.2026486, 0.2618968, 0.3547908, 
    0.297543, 0.1503338, 0.3236479, 0.237551, 0.1966092, 0.1033061, 
    0.04063004, 0.09474317, 0.05587334, 0.1372223, 0.1012477, 0.2004278,
  0.2948124, 0.2842137, 0.1408406, 0.1646208, 0.401653, 0.3213618, 0.1796096, 
    0.1718374, 0.2130511, 0.2517143, 0.2775761, 0.176545, 0.2248289, 
    0.4041137, 0.3376143, 0.2394662, 0.2100229, 0.2665035, 0.2271232, 
    0.3131756, 0.1547527, 0.1369891, 0.2380105, 0.2123548, 0.2049699, 
    0.132575, 0.1581543, 0.1435553, 0.3191988,
  0.2534137, 0.3081811, 0.3563576, 0.2921126, 0.2461947, 0.2819603, 
    0.2909782, 0.3562482, 0.3318395, 0.3348682, 0.2999518, 0.2855109, 
    0.2455383, 0.2057985, 0.257203, 0.219429, 0.2658384, 0.2140183, 0.249178, 
    0.204105, 0.225301, 0.2662856, 0.280222, 0.2336365, 0.2349138, 0.2101099, 
    0.1777323, 0.2744493, 0.2849621,
  0.1821774, 0.1774102, 0.1865422, 0.194705, 0.176004, 0.2006721, 0.2198358, 
    0.2019465, 0.2164512, 0.1928145, 0.1854864, 0.1296307, 0.1866181, 
    0.245783, 0.2216724, 0.1530011, 0.1215484, 0.1162573, 0.1115212, 
    0.1191993, 0.1519376, 0.2131034, 0.2059717, 0.1359046, 0.1158693, 
    0.1404807, 0.1469294, 0.1528949, 0.1722713,
  0.04637339, 0.02924107, 0.01900031, 0.05228952, 0.103055, 0.06514028, 
    0.0762791, 0.04537741, 0.03708437, 0.01327532, 0.017631, 0.05963806, 
    0.073954, 0.03957172, 0.03843167, 0.02020743, 0.06573386, 0.07826795, 
    0.1112931, 0.132854, 0.06713431, 0.02303423, 0.01205714, 0.02697566, 
    0.05759057, 0.04838707, 0.07778285, 0.09867956, 0.05979321,
  0.0002093069, -4.863718e-06, 0.1259312, 0.05376435, 0.04245657, 0.02842961, 
    0.006420062, 0.001496752, -1.946901e-05, 0.06136178, 0.05066349, 
    0.04651612, 0.1077742, 0.005675423, 0.04822297, 0.0002433905, 0.1011942, 
    0.1184691, 0.04330438, 0.1789191, 0.005966464, 0.0001262444, 
    1.507128e-07, 0.001436908, 0.02497408, 0.0807628, 0.1155333, 0.007515823, 
    5.674696e-05,
  1.796026e-05, 0.1582915, 0.1276952, 0.01121041, 0.08793937, 0.03330711, 
    0.0332538, -0.0002943907, 0.002445224, 0.08073087, 0.08726464, 
    0.06066807, 0.07408836, 0.03797469, 0.03489473, 0.1615181, 0.1022306, 
    0.1374572, 0.03767518, 0.0165041, 0.00131954, 8.863823e-09, 2.469093e-06, 
    0.002540564, 0.1460117, 0.1906722, 0.02875892, 0.0004968675, -8.300624e-06,
  0.000177549, 0.01664206, 0.3901995, 0.1459407, 0.07715938, 0.07001971, 
    0.08578745, 0.04352956, 0.0113234, 0.03183049, 0.04960852, 0.02909606, 
    0.06339501, 0.01823539, 0.03665861, 0.1315456, 0.06784116, 0.03129828, 
    0.005861125, -1.014906e-06, 8.170392e-08, -7.590857e-07, 3.388509e-05, 
    0.1021434, 0.4102653, 0.1566526, 0.02788545, 0.0003105912, 0.0001663104,
  0.05330837, 0.05729457, 0.02406094, 0.025865, 0.03720862, 0.02116501, 
    0.1366394, 0.04890799, 0.08541902, 0.2774361, 0.005831827, 0.004456319, 
    0.04428484, 0.0378022, 0.07751754, 0.01463237, 0.002477031, 0.000617242, 
    0.0006981019, 0.004473968, 0.003910162, 0.0804903, 0.09250271, 
    0.05536911, 0.1615114, 0.1702249, 0.03478317, 0.007225591, 0.01697079,
  -1.858244e-06, 6.631683e-06, 2.437765e-06, 0.02978329, 1.51962e-05, 
    0.02105353, 0.01928596, 0.0835288, 0.004229483, 0.08702549, 0.2180181, 
    0.1217673, 0.06376614, 0.04893833, 0.01268699, 0.01940935, 0.04119109, 
    0.03757399, 0.04062388, 0.06186579, 0.0632733, 0.04013497, 0.006166412, 
    0.005036352, 0.01008118, 0.007650412, -0.0003841125, 0.0004745547, 
    0.004371565,
  0.0001333463, 4.956072e-06, 1.288288e-06, 0.0001026613, 2.903739e-06, 
    0.006688063, 1.564023e-05, 0.005457271, 0.01549278, -0.0002502972, 
    0.1346684, 0.0834057, 0.05020671, 0.0004572954, -3.984662e-07, 
    -4.377497e-06, 0.01392484, 0.01087426, 0.002207616, 0.001838512, 
    0.02631531, 0.05082104, 0.0658915, 0.01532643, 0.01616274, 0.005044589, 
    0.004587386, 0.01130523, 0.03406239,
  0.007073888, 0.03789158, 0.01605265, 0.007783851, 0.04598033, 0.02600111, 
    0.01956336, 0.03186655, 0.1301328, 0.1492252, 0.06408689, 0.04912154, 
    0.0733994, 0.1445449, 0.1026328, 0.135339, 0.1165837, 0.08572562, 
    0.05181303, 0.008089569, 0.01535913, 0.03757297, 0.06846919, 0.05979282, 
    0.09493488, 0.09808658, 0.08075827, 0.02131749, 0.00293629,
  0.08800994, 0.1361721, 0.2140637, 0.3175672, 0.09901529, 0.05616292, 
    0.3523974, 0.02067502, 0.05352925, 0.03054138, 0.08371644, 0.0972937, 
    0.1409906, 0.1589988, 0.1978507, 0.2150378, 0.2142421, 0.197658, 0.1359, 
    0.1763251, 0.1640527, 0.07094587, 0.1062963, 0.1043349, 0.1731246, 
    0.1481615, 0.1156216, 0.04502214, 0.1269194,
  0.2041505, 0.21919, 0.1847979, 0.2630713, 0.249262, 0.2103969, 0.112894, 
    0.1075379, 0.0858572, 0.08089561, 0.06193547, 0.1883399, 0.1361445, 
    0.2843679, 0.1779849, 0.096343, 0.09484749, 0.1394661, 0.144485, 
    0.2246247, 0.1059973, 0.1785824, 0.2040565, 0.3129365, 0.2685905, 
    0.1628466, 0.1718872, 0.1549254, 0.1814786,
  0.2030305, 0.2010772, 0.209386, 0.3175585, 0.239408, 0.3565283, 0.3518959, 
    0.3252398, 0.2451093, 0.2222538, 0.238215, 0.1992059, 0.1833111, 
    0.1975057, 0.1379808, 0.08777644, 0.1506281, 0.2673501, 0.2772774, 
    0.1575499, 0.1636726, 0.128256, 0.1953308, 0.256822, 0.1740976, 
    0.3078324, 0.2394705, 0.3347917, 0.1834314,
  0.1610522, 0.1565399, 0.2839798, 0.3319641, 0.3230737, 0.3091026, 
    0.2799943, 0.3812483, 0.2253685, 0.2444068, 0.2613569, 0.2511376, 
    0.2788279, 0.2297329, 0.2470399, 0.1359613, 0.266747, 0.3646972, 
    0.4051102, 0.3629017, 0.2512009, 0.1822125, 0.1786713, 0.2327875, 
    0.2815318, 0.2966022, 0.102914, 0.153959, 0.1404151,
  0.225641, 0.2526156, 0.2272813, 0.1489414, 0.1691718, 0.2067081, 0.1933488, 
    0.1664824, 0.2059061, 0.1958364, 0.1989047, 0.1725618, 0.1723011, 
    0.1863235, 0.2068845, 0.2274069, 0.1813151, 0.1596057, 0.1461899, 
    0.1279191, 0.1998637, 0.1729535, 0.1205254, 0.06423213, 0.1242223, 
    0.01496612, 0.04785366, 0.2168736, 0.2642549,
  0.07082365, 0.06972443, 0.06862522, 0.06752601, 0.0664268, 0.06532758, 
    0.06422837, 0.04802161, 0.05191779, 0.05581397, 0.05971016, 0.06360634, 
    0.06750252, 0.0713987, 0.09945761, 0.09912524, 0.09879287, 0.09846051, 
    0.09812815, 0.09779578, 0.09746341, 0.1033577, 0.1008931, 0.09842849, 
    0.09596389, 0.09349928, 0.09103467, 0.08857007, 0.07170302,
  0.2560496, 0.269366, 0.237291, 0.145137, 0.09962125, 0.07562226, 
    0.06229747, 0.03800704, 0.01383411, 0.01582247, 0.136904, 0.1244114, 
    0.1939612, 0.2475553, 0.1945606, 0.2929043, 0.3243831, 0.3023002, 
    0.1359079, 0.3116316, 0.2651066, 0.2115086, 0.1158029, 0.05730011, 
    0.07372011, 0.0612432, 0.1105439, 0.107712, 0.1825913,
  0.230407, 0.1836414, 0.1019916, 0.1893559, 0.3708786, 0.288459, 0.1594685, 
    0.1745805, 0.2149334, 0.2691946, 0.2486261, 0.1733562, 0.2814307, 
    0.3850233, 0.3142743, 0.2414707, 0.1892194, 0.2806998, 0.2479731, 
    0.2159989, 0.2472581, 0.254735, 0.3077984, 0.2349256, 0.2151255, 
    0.1277999, 0.2347215, 0.256994, 0.2713107,
  0.2681254, 0.3578939, 0.3683714, 0.3311998, 0.2768773, 0.3811679, 
    0.4144224, 0.2829394, 0.4035628, 0.3259031, 0.2758598, 0.2902638, 
    0.2704806, 0.2358575, 0.2421957, 0.2486176, 0.2420785, 0.1971324, 
    0.2286261, 0.2273501, 0.2290936, 0.2738029, 0.2493603, 0.2319627, 
    0.2543204, 0.226017, 0.1937381, 0.2299739, 0.2680541,
  0.2282313, 0.2393432, 0.1976598, 0.2027849, 0.1648803, 0.2150331, 
    0.1941177, 0.2038936, 0.1968358, 0.2036017, 0.1759014, 0.1658189, 
    0.1980739, 0.2520825, 0.215416, 0.1398806, 0.1235221, 0.1209868, 
    0.1116935, 0.1177873, 0.1734181, 0.1996796, 0.2056496, 0.1503636, 
    0.125868, 0.1219672, 0.1626659, 0.1587371, 0.1651955,
  0.04886576, 0.03385666, 0.02066593, 0.03800271, 0.1213497, 0.06816658, 
    0.07305216, 0.05989119, 0.0500681, 0.01571461, 0.0213969, 0.04513681, 
    0.05564159, 0.04228401, 0.05225025, 0.02513973, 0.07552913, 0.09585167, 
    0.1241815, 0.1268163, 0.07574337, 0.03305254, 0.02941421, 0.05333555, 
    0.04193857, 0.04757771, 0.08971315, 0.1071971, 0.07902362,
  0.0004347435, -1.23376e-06, 0.1390344, 0.04489859, 0.02215649, 0.01494063, 
    0.009415258, 0.003305702, -2.935098e-06, 0.03438746, 0.01954071, 
    0.008807246, 0.1028232, 0.002220035, 0.04032629, 0.0007444072, 
    0.07928029, 0.1142969, 0.05532498, 0.164939, 0.007409559, 0.0004735848, 
    -4.025051e-07, 0.001253862, 0.02581813, 0.05607658, 0.1115791, 
    0.01333684, 0.0001340138,
  1.21474e-05, 0.1394617, 0.1280005, 0.01253395, 0.08490399, 0.03105243, 
    0.02948761, 6.458414e-05, 0.001178376, 0.07525889, 0.07305545, 
    0.05422845, 0.07360627, 0.0234382, 0.03230206, 0.157543, 0.07792502, 
    0.09307258, 0.04187465, 0.02228362, 0.006197341, 2.43765e-08, 
    4.292835e-07, 0.0005376737, 0.1483494, 0.2011998, 0.02551598, 
    0.001915101, -4.76676e-07,
  -3.959209e-05, 0.001503919, 0.4154265, 0.09593888, 0.07316441, 0.05143213, 
    0.06118971, 0.04408418, 0.01323208, 0.02794047, 0.04196041, 0.02107527, 
    0.05793063, 0.01696087, 0.03431261, 0.1196383, 0.0700987, 0.03244393, 
    0.01095775, 0.000469076, 1.453586e-07, 7.899455e-07, 5.33916e-06, 
    0.04916294, 0.2689543, 0.1142331, 0.02872993, 0.0008798721, -7.734298e-05,
  0.01575661, 0.03762015, 0.02016619, 0.02566126, 0.03094468, 0.03269488, 
    0.1024049, 0.04719842, 0.08679359, 0.2304993, 0.007795207, 0.004698551, 
    0.03933126, 0.02843125, 0.05712165, 0.01528079, 0.003272464, 
    0.0006319863, 0.004485239, 0.008508406, 0.00728749, 0.0397576, 0.1052366, 
    0.04129898, 0.130655, 0.165648, 0.0469257, 0.006638904, 0.006711297,
  5.10312e-07, 3.001816e-06, -6.833224e-06, 0.05472543, 0.0001979298, 
    0.03724004, 0.007591269, 0.08116972, 0.009949182, 0.06311152, 0.2300052, 
    0.1070598, 0.05085561, 0.03116633, 0.01812094, 0.03352745, 0.04294411, 
    0.0321479, 0.02267279, 0.0573706, 0.05759345, 0.03468182, 0.01464841, 
    0.006317837, 0.0124349, 0.001949669, 0.0004655478, 2.882879e-06, 
    0.005776663,
  1.170994e-05, 1.895477e-06, 4.767505e-07, 9.457072e-05, 0.02338325, 
    0.01003696, 1.132176e-05, 0.009248141, 0.01950925, -0.0001592604, 
    0.1275062, 0.05492618, 0.05818107, -1.201794e-05, 5.496902e-07, 
    9.625751e-05, 0.005449235, 0.01066918, 0.001972333, 0.004700982, 
    0.02410758, 0.05896178, 0.06468518, 0.03723942, 0.01594042, 0.01329314, 
    0.004475, 0.003468202, 0.003836676,
  0.01562901, 0.03298365, 0.01114091, 0.007405342, 0.05506731, 0.03098714, 
    0.01692673, 0.03061341, 0.1406233, 0.172327, 0.05114786, 0.05141501, 
    0.1019179, 0.1524363, 0.104755, 0.1484891, 0.1139926, 0.08369146, 
    0.0588336, 0.002879033, 0.008397533, 0.04776764, 0.06903221, 0.06851372, 
    0.1078506, 0.1117047, 0.08529349, 0.02174496, 0.005584827,
  0.08124594, 0.1219036, 0.2042026, 0.3400542, 0.1252073, 0.04736295, 
    0.3516619, 0.01408997, 0.03615505, 0.02356222, 0.07968407, 0.09722187, 
    0.1661711, 0.1570828, 0.2020065, 0.2213025, 0.1948316, 0.2010905, 
    0.1386381, 0.181171, 0.1639373, 0.06338289, 0.1120305, 0.121086, 
    0.190275, 0.1463527, 0.1296891, 0.05554046, 0.1182252,
  0.1994633, 0.2245175, 0.217746, 0.2830497, 0.2343232, 0.1877075, 
    0.09871579, 0.1054912, 0.08399647, 0.0808056, 0.06901786, 0.1730131, 
    0.1405578, 0.2864921, 0.2254582, 0.1119599, 0.1051463, 0.1459135, 
    0.1502409, 0.2313726, 0.1229727, 0.1742563, 0.2044806, 0.3555659, 
    0.2765242, 0.1723243, 0.1972902, 0.1663111, 0.1939689,
  0.2175259, 0.2007672, 0.2329118, 0.3646733, 0.2641326, 0.3427913, 0.36285, 
    0.32212, 0.2404164, 0.2193995, 0.2430482, 0.2057932, 0.1931053, 
    0.2039916, 0.1417022, 0.1088791, 0.1659, 0.283646, 0.3018921, 0.1546172, 
    0.1612424, 0.1563786, 0.1948794, 0.250279, 0.1817401, 0.3128943, 
    0.2636601, 0.3462334, 0.1983045,
  0.174685, 0.1828386, 0.3007276, 0.3482092, 0.3385208, 0.321917, 0.3099622, 
    0.3980577, 0.2370445, 0.2306696, 0.2552628, 0.3001685, 0.3247839, 
    0.2303494, 0.2543841, 0.1626957, 0.2931461, 0.3633702, 0.4089831, 
    0.3734288, 0.2402062, 0.1809181, 0.231738, 0.3072093, 0.268241, 
    0.3575844, 0.1299058, 0.1597492, 0.1612235,
  0.2211671, 0.2385217, 0.2118593, 0.1445686, 0.1661389, 0.1977114, 0.187826, 
    0.1737542, 0.2134693, 0.1850557, 0.2280674, 0.2120852, 0.219421, 
    0.3168217, 0.3527227, 0.360522, 0.304317, 0.2062082, 0.1812213, 
    0.1587543, 0.2404853, 0.1960386, 0.1174293, 0.1019437, 0.1465813, 
    0.03632773, 0.08903243, 0.1987186, 0.2664195,
  0.07199486, 0.06983482, 0.06767479, 0.06551475, 0.06335472, 0.06119468, 
    0.05903465, 0.05727842, 0.06073736, 0.06419629, 0.06765523, 0.07111416, 
    0.0745731, 0.07803203, 0.108493, 0.1098127, 0.1111324, 0.1124521, 
    0.1137718, 0.1150915, 0.1164112, 0.1199275, 0.1173089, 0.1146903, 
    0.1120717, 0.1094531, 0.1068345, 0.1042159, 0.07372288,
  0.228195, 0.2628424, 0.2521629, 0.240318, 0.1478631, 0.1131822, 0.130764, 
    0.09690775, 0.01517622, 0.1723459, 0.1557173, 0.1244672, 0.2076006, 
    0.1991893, 0.1536932, 0.3241965, 0.3531649, 0.2637236, 0.1713631, 
    0.3484079, 0.2820216, 0.2382639, 0.1080707, 0.05841375, 0.07764569, 
    0.06083959, 0.08775719, 0.1262838, 0.1502497,
  0.270108, 0.2387877, 0.1350628, 0.198345, 0.347638, 0.2861773, 0.1380807, 
    0.1706176, 0.2074856, 0.2636341, 0.2596637, 0.1690375, 0.281513, 
    0.3535795, 0.3367543, 0.2676538, 0.1545981, 0.2176529, 0.2260134, 
    0.212613, 0.2489927, 0.26494, 0.3821166, 0.262346, 0.2426507, 0.1804286, 
    0.2227816, 0.3162321, 0.3180916,
  0.2611543, 0.4450341, 0.392908, 0.3345445, 0.3871278, 0.3910132, 0.3460116, 
    0.3814792, 0.375568, 0.3299104, 0.3174753, 0.2660842, 0.2857648, 
    0.2327133, 0.3180896, 0.2472998, 0.293895, 0.2170787, 0.2783349, 
    0.2463422, 0.2503344, 0.3037593, 0.3057067, 0.2663527, 0.2770685, 
    0.2333819, 0.2507578, 0.3010311, 0.302221,
  0.2571795, 0.2097327, 0.2060699, 0.217209, 0.1860886, 0.2396459, 0.2175048, 
    0.1941815, 0.2082431, 0.2233552, 0.1773721, 0.1694252, 0.2109236, 
    0.2479316, 0.2201708, 0.1734468, 0.1384996, 0.1415154, 0.1608042, 
    0.1234063, 0.202708, 0.2078774, 0.2201784, 0.1570703, 0.11664, 0.1078512, 
    0.164765, 0.1703393, 0.1981431,
  0.04889676, 0.04083532, 0.03169136, 0.04011914, 0.1108514, 0.06731309, 
    0.07744316, 0.06822808, 0.05673156, 0.02323286, 0.02846439, 0.01949821, 
    0.04592812, 0.0322613, 0.06280452, 0.0564301, 0.08516289, 0.0947319, 
    0.1045045, 0.1343019, 0.07011172, 0.03188455, 0.03610918, 0.04818671, 
    0.03287484, 0.04854752, 0.09660629, 0.1040338, 0.07664641,
  0.001409864, 1.616108e-06, 0.1503063, 0.03785196, 0.02830968, 0.01100271, 
    0.009790001, 0.004707304, -6.396414e-06, 0.01482588, 0.007413333, 
    0.0004789728, 0.08680578, 0.00201064, 0.04516071, 0.002087409, 
    0.07428198, 0.1144231, 0.05480909, 0.1051678, 0.009500365, 0.001053836, 
    -5.266025e-06, 0.0008188599, 0.02953684, 0.04880996, 0.1063418, 
    0.02055896, 0.0007128951,
  6.335358e-06, 0.1148673, 0.1086227, 0.01915611, 0.08032241, 0.03074351, 
    0.0273192, 0.0008839878, 0.0004439061, 0.06469061, 0.06911885, 
    0.06029827, 0.08519986, 0.02282293, 0.03417525, 0.1594832, 0.07213641, 
    0.06611988, 0.04603948, 0.05337785, 0.0186887, 2.044767e-07, 
    7.762132e-08, -0.0002165576, 0.167193, 0.1641789, 0.02562855, 
    0.004796945, -1.47153e-06,
  -7.537949e-06, -0.0006504453, 0.3319691, 0.07754162, 0.06658107, 
    0.04475877, 0.05154025, 0.05207692, 0.01688693, 0.0265632, 0.03551993, 
    0.01716327, 0.04907827, 0.01602857, 0.03384237, 0.1148555, 0.07129967, 
    0.05067128, 0.0251982, 0.007084599, 1.306046e-05, 4.603271e-07, 
    2.615043e-06, 0.04216827, 0.2154536, 0.0956594, 0.03658399, 0.001644086, 
    7.396179e-06,
  0.009351894, 0.01380571, 0.01673059, 0.0418974, 0.03176435, 0.02681591, 
    0.08959347, 0.03876681, 0.1056966, 0.2215835, 0.009162713, 0.005178744, 
    0.03753501, 0.02106696, 0.0420894, 0.02015407, 0.005326188, 0.0005469896, 
    0.0106537, 0.0125013, 0.008768024, 0.0171733, 0.08021167, 0.0471127, 
    0.113665, 0.1626428, 0.05229629, 0.01053347, 0.003217568,
  2.648058e-07, 1.895962e-06, 6.613247e-07, 0.06412885, 0.001166927, 
    0.05104107, 0.006358335, 0.0769105, 0.0201103, 0.08065904, 0.2334942, 
    0.1017883, 0.05017926, 0.02654924, 0.01912335, 0.03613083, 0.03951168, 
    0.02501042, 0.01786105, 0.05107901, 0.05408942, 0.03274602, 0.03259502, 
    0.01180658, 0.01889176, 0.001039664, 0.0003151395, 2.701251e-07, 
    0.001411658,
  6.628799e-06, 9.199727e-07, 2.1599e-07, 0.0002845734, 0.007259917, 
    0.009986018, 2.012666e-05, 0.01424042, 0.02302553, -0.0003982745, 
    0.1073365, 0.03395258, 0.06134881, 0.0003115107, 0.001008593, 
    0.0006013514, 0.00794222, 0.00812665, 0.001163271, 0.00264823, 
    0.02203299, 0.07499731, 0.06092751, 0.06734734, 0.02161157, 0.02073617, 
    0.004587964, 8.651125e-05, 2.778238e-05,
  0.02261413, 0.03650177, 0.007161949, 0.0123349, 0.05899869, 0.03553602, 
    0.01100131, 0.03348808, 0.1213335, 0.1645377, 0.04157173, 0.06747968, 
    0.1188529, 0.1451746, 0.1041709, 0.1678905, 0.1183009, 0.08121929, 
    0.0688252, 0.002048464, 0.00570543, 0.05888697, 0.0762265, 0.08740283, 
    0.1186416, 0.1190576, 0.09257898, 0.03127305, 0.006888893,
  0.0779694, 0.1129995, 0.188703, 0.3568318, 0.1387434, 0.03855019, 
    0.3544337, 0.01023374, 0.01867228, 0.01953205, 0.08053403, 0.1149049, 
    0.1741925, 0.1676442, 0.2113215, 0.2357225, 0.1989898, 0.2123944, 
    0.1579541, 0.1942725, 0.1738921, 0.07326061, 0.1479577, 0.1409327, 
    0.2041634, 0.1540004, 0.1454933, 0.08557045, 0.1275881,
  0.199875, 0.195116, 0.1776047, 0.2373798, 0.2313626, 0.1771546, 0.09503631, 
    0.1014528, 0.08791455, 0.06801422, 0.07072058, 0.1659834, 0.1592567, 
    0.3008272, 0.2481041, 0.1513108, 0.1372868, 0.1397298, 0.1514752, 
    0.2426073, 0.106974, 0.1704792, 0.2003703, 0.3151264, 0.2500141, 
    0.1989007, 0.1813876, 0.1694283, 0.1850937,
  0.2086017, 0.2013288, 0.2172003, 0.3770013, 0.2924255, 0.3049914, 
    0.4128187, 0.3280397, 0.2556009, 0.2416139, 0.2478531, 0.2023237, 
    0.2065315, 0.2080107, 0.1724263, 0.1003463, 0.1871977, 0.3136394, 
    0.3135282, 0.1589825, 0.1925555, 0.1299993, 0.1961785, 0.2164431, 
    0.2084167, 0.329877, 0.277371, 0.3358914, 0.2045781,
  0.2158468, 0.2502865, 0.3145017, 0.3054282, 0.3237877, 0.3706982, 
    0.3141899, 0.4387285, 0.2392507, 0.2212462, 0.2380756, 0.3594863, 
    0.3153784, 0.229116, 0.2652295, 0.1802847, 0.2839377, 0.3746017, 
    0.3609786, 0.3358147, 0.3020908, 0.2084924, 0.2618453, 0.3003063, 
    0.2379314, 0.3866895, 0.1346715, 0.1713622, 0.2144724,
  0.2146259, 0.2437685, 0.2131707, 0.1554883, 0.1666251, 0.2016201, 
    0.1865087, 0.1680383, 0.2048256, 0.2146861, 0.2726348, 0.2334885, 
    0.2582422, 0.3181087, 0.4129278, 0.4373316, 0.3412019, 0.1858174, 
    0.1998141, 0.1564015, 0.2579356, 0.2142557, 0.124252, 0.09804947, 
    0.1579337, 0.05973439, 0.1490173, 0.1933227, 0.2810833,
  0.09812149, 0.09578804, 0.09345459, 0.09112114, 0.0887877, 0.08645425, 
    0.0841208, 0.0792889, 0.08119854, 0.08310816, 0.0850178, 0.08692744, 
    0.08883707, 0.09074671, 0.1163413, 0.118908, 0.1214747, 0.1240414, 
    0.1266081, 0.1291748, 0.1317415, 0.1398999, 0.137757, 0.1356141, 
    0.1334712, 0.1313284, 0.1291855, 0.1270426, 0.09998824,
  0.2298899, 0.2502919, 0.2584889, 0.2604323, 0.1913023, 0.1313418, 
    0.1822803, 0.1626195, 0.1050613, 0.242863, 0.152464, 0.134285, 0.2335278, 
    0.1671988, 0.167303, 0.2667588, 0.2857472, 0.2090181, 0.2400911, 
    0.3210686, 0.2517062, 0.2506117, 0.1083818, 0.04788801, 0.06489641, 
    0.04415599, 0.07425418, 0.1146566, 0.1598505,
  0.2165564, 0.1903808, 0.1163136, 0.1767427, 0.3013662, 0.2980725, 
    0.1405174, 0.1658481, 0.18831, 0.2150116, 0.2595209, 0.16105, 0.2666838, 
    0.3360998, 0.2969834, 0.2745115, 0.1390808, 0.2144546, 0.3199214, 
    0.1801464, 0.1293133, 0.2177044, 0.3008061, 0.2990615, 0.2426103, 
    0.1304595, 0.1747134, 0.3023573, 0.2740983,
  0.3241018, 0.3582062, 0.3542485, 0.383353, 0.4280885, 0.4748853, 0.3375246, 
    0.3419767, 0.4231944, 0.3330669, 0.3294964, 0.3540594, 0.2916991, 
    0.2473483, 0.2861181, 0.288253, 0.2984816, 0.2568073, 0.2613443, 
    0.2301719, 0.2254473, 0.2718096, 0.2788645, 0.2646459, 0.2474395, 
    0.2266562, 0.2043568, 0.3082276, 0.3486141,
  0.2491677, 0.2306693, 0.1965518, 0.2060937, 0.213729, 0.2416357, 0.2153621, 
    0.2427581, 0.2328305, 0.2107062, 0.207053, 0.2083987, 0.2413312, 
    0.2621765, 0.2445477, 0.1929277, 0.1499246, 0.1416963, 0.1908426, 
    0.1330317, 0.2087043, 0.2453658, 0.2565088, 0.1683422, 0.1120855, 
    0.09595462, 0.1596717, 0.1797943, 0.2206349,
  0.05036892, 0.04908193, 0.04558811, 0.04305314, 0.1099815, 0.06892207, 
    0.08053297, 0.08668758, 0.07088318, 0.02933395, 0.02158638, 0.008152676, 
    0.04688577, 0.037593, 0.06864041, 0.058967, 0.1046572, 0.09112279, 
    0.094249, 0.1252008, 0.07196525, 0.02666439, 0.04630549, 0.04899792, 
    0.02335779, 0.04552903, 0.1095902, 0.09536713, 0.08744273,
  0.001997468, 0.0001437554, 0.1141877, 0.03843388, 0.04490617, 0.01639008, 
    0.01377621, 0.009488993, 0.0002287854, 0.01078422, 0.002054063, 
    3.920129e-05, 0.07060387, 0.004878112, 0.05030135, 0.004359683, 
    0.07348023, 0.1086976, 0.04603855, 0.07986576, 0.01790111, 0.004882047, 
    3.393724e-05, 0.0003917792, 0.04813349, 0.04338513, 0.107187, 0.03238055, 
    0.005163881,
  1.980466e-06, 0.08696243, 0.1254798, 0.02533213, 0.07536222, 0.04252784, 
    0.04043089, 0.005794254, 0.0004128437, 0.05376682, 0.0620072, 0.05547073, 
    0.09088372, 0.02556143, 0.03714646, 0.1620924, 0.05519023, 0.05601168, 
    0.03618865, 0.04875742, 0.07234468, 0.001023152, 2.905904e-07, 
    -0.0002352337, 0.1889448, 0.1552035, 0.04881797, 0.02753241, 0.000453522,
  8.042815e-07, -0.0005213716, 0.2998961, 0.06432801, 0.05794522, 0.0424945, 
    0.0518663, 0.05678084, 0.0233735, 0.02853129, 0.03593056, 0.01654423, 
    0.04516453, 0.01522006, 0.03374154, 0.09064081, 0.07276789, 0.04954731, 
    0.02998897, 0.007579671, 0.0007676855, 2.364033e-05, 3.579483e-05, 
    0.04300436, 0.170853, 0.08949922, 0.04517509, 0.003161702, 0.0001479137,
  0.007680495, 0.006111559, 0.01686104, 0.04133179, 0.03455013, 0.03060817, 
    0.07967158, 0.03634018, 0.1388365, 0.2128513, 0.01131273, 0.006588823, 
    0.0350628, 0.02189076, 0.03495071, 0.02186756, 0.008087662, 0.004555598, 
    0.0185652, 0.02352897, 0.01235368, 0.01905029, 0.07602542, 0.04797771, 
    0.09692094, 0.1512461, 0.05189653, 0.02514509, 0.005725517,
  1.028779e-07, 8.209698e-07, 2.799177e-07, 0.05175591, 0.003602726, 
    0.05756529, 0.01416204, 0.0759335, 0.02976224, 0.1050237, 0.2531599, 
    0.1011707, 0.04988028, 0.02918695, 0.022881, 0.04036097, 0.02995924, 
    0.02000863, 0.0241994, 0.04854591, 0.05412919, 0.03988922, 0.06065439, 
    0.01919974, 0.03466611, 0.001578951, 0.0003140115, -2.991072e-07, 
    -2.096253e-05,
  4.115275e-06, 5.128563e-07, 1.032235e-07, 0.001016198, 0.0002075605, 
    0.007723037, 0.0004059713, 0.02805934, 0.02794411, -0.0004336204, 
    0.07203772, 0.04184286, 0.07624301, 0.0003570642, 0.002093281, 
    0.003765143, 0.01814831, 0.01006973, 0.000663762, 0.003850868, 
    0.01809908, 0.1098782, 0.05798162, 0.09657307, 0.02572421, 0.02112379, 
    0.01123061, -3.459246e-06, 2.759694e-06,
  0.0114355, 0.006943634, 0.008719128, 0.01350451, 0.05531874, 0.03505479, 
    0.008571824, 0.03107358, 0.1127452, 0.1189481, 0.03739258, 0.10763, 
    0.1321688, 0.1451797, 0.1066566, 0.1654217, 0.1139174, 0.07790143, 
    0.06739824, 0.01429033, 0.01552261, 0.06302462, 0.07369169, 0.08752206, 
    0.1172863, 0.1226512, 0.08855715, 0.03720403, 0.006943122,
  0.07485463, 0.1189931, 0.1791356, 0.364123, 0.1474063, 0.04794673, 
    0.3504911, 0.01126602, 0.01147346, 0.01505933, 0.07389951, 0.1592678, 
    0.1746494, 0.1865187, 0.2453209, 0.25151, 0.2270882, 0.2188457, 
    0.1700532, 0.216867, 0.167812, 0.05438943, 0.1347617, 0.1314145, 
    0.2448986, 0.1587798, 0.1600604, 0.08425831, 0.1416546,
  0.2040566, 0.1923495, 0.2000016, 0.2011412, 0.2134887, 0.1786516, 
    0.08585417, 0.1028331, 0.08889586, 0.05307551, 0.07060014, 0.169999, 
    0.1715956, 0.3185094, 0.2869745, 0.1855482, 0.1432101, 0.1593613, 
    0.1510779, 0.2379638, 0.09515446, 0.1775601, 0.2380868, 0.2650197, 
    0.2351244, 0.1917589, 0.2120912, 0.1875547, 0.1899423,
  0.2562014, 0.2323956, 0.185122, 0.3708671, 0.2849815, 0.34445, 0.4024571, 
    0.3254688, 0.2698889, 0.2676663, 0.2608416, 0.1917276, 0.2114758, 
    0.2180766, 0.1936726, 0.09310359, 0.1994836, 0.3426034, 0.3014426, 
    0.153755, 0.2002099, 0.1247334, 0.1746821, 0.2146348, 0.1719923, 
    0.3428917, 0.3031012, 0.3416546, 0.2675149,
  0.2296666, 0.3059205, 0.310178, 0.3459743, 0.2941398, 0.365979, 0.3798456, 
    0.460112, 0.2446018, 0.2314576, 0.2694528, 0.3989337, 0.3390227, 
    0.2449603, 0.2955417, 0.1845615, 0.2508661, 0.4095096, 0.3154249, 
    0.2922751, 0.3123659, 0.2068596, 0.2574733, 0.2215325, 0.2325782, 
    0.4243263, 0.1212835, 0.1681082, 0.2257389,
  0.2320511, 0.2653683, 0.2101011, 0.1503262, 0.1949159, 0.2410375, 
    0.1972779, 0.1789749, 0.1847216, 0.2301775, 0.2760635, 0.2497641, 
    0.2736025, 0.323177, 0.3945145, 0.4493248, 0.3295735, 0.1668403, 
    0.2280553, 0.1813233, 0.2591712, 0.2222986, 0.1391127, 0.1061608, 
    0.1558623, 0.0839877, 0.1232728, 0.1975699, 0.2921595,
  0.1267387, 0.1250323, 0.1233259, 0.1216195, 0.1199132, 0.1182068, 
    0.1165004, 0.119056, 0.118644, 0.118232, 0.11782, 0.1174081, 0.1169961, 
    0.1165841, 0.1180754, 0.1196239, 0.1211725, 0.122721, 0.1242695, 
    0.125818, 0.1273666, 0.1450854, 0.1456552, 0.1462251, 0.1467949, 
    0.1473647, 0.1479345, 0.1485044, 0.1281038,
  0.2373341, 0.2178164, 0.2850004, 0.2633871, 0.1809406, 0.1588729, 0.237067, 
    0.2990479, 0.0873994, 0.23242, 0.1585751, 0.129557, 0.2837545, 0.113776, 
    0.1248824, 0.2029339, 0.2536363, 0.1602911, 0.233447, 0.2647225, 
    0.2452144, 0.2541555, 0.07767094, 0.08132558, 0.01117913, 0.08167906, 
    0.1123798, 0.0989681, 0.1978717,
  0.2214868, 0.1883933, 0.1888925, 0.1581721, 0.2798815, 0.3121749, 
    0.1382909, 0.1712617, 0.1606979, 0.1808588, 0.2406571, 0.1678378, 
    0.2824696, 0.2972034, 0.2580721, 0.1873766, 0.1325506, 0.1869366, 
    0.2648646, 0.2884347, 0.08059277, 0.1177379, 0.2316505, 0.2644808, 
    0.1800828, 0.1513083, 0.1664297, 0.3242827, 0.2392855,
  0.3175586, 0.3809126, 0.3531239, 0.3700925, 0.3977169, 0.3992243, 
    0.3169098, 0.267904, 0.4095755, 0.3615281, 0.3470644, 0.3048765, 
    0.2369356, 0.2309198, 0.23821, 0.277328, 0.2803371, 0.2425911, 0.2250843, 
    0.229424, 0.2063428, 0.2534007, 0.2640943, 0.2608802, 0.2335624, 
    0.2157148, 0.1952039, 0.2626678, 0.3224214,
  0.2385697, 0.2171837, 0.1995593, 0.2041727, 0.2311235, 0.2241599, 
    0.2288242, 0.2741814, 0.2741034, 0.208926, 0.2219843, 0.2307948, 
    0.2728103, 0.2717508, 0.2435595, 0.193872, 0.1550391, 0.1472659, 
    0.1676916, 0.1412704, 0.2119431, 0.2491559, 0.2750903, 0.1778799, 
    0.102478, 0.1004233, 0.1585222, 0.16273, 0.207741,
  0.05848797, 0.06782576, 0.07467506, 0.06448202, 0.1346917, 0.07195735, 
    0.09368165, 0.09955665, 0.09753286, 0.03340801, 0.01694792, 0.005752006, 
    0.05315796, 0.04054216, 0.07525748, 0.06247455, 0.1416913, 0.08220871, 
    0.09392673, 0.127123, 0.09924645, 0.03852177, 0.06914625, 0.05745037, 
    0.01376022, 0.04222668, 0.1340818, 0.08836763, 0.09083366,
  0.007780862, 0.008336442, 0.1002604, 0.05691117, 0.03344075, 0.03298097, 
    0.02362495, 0.02564972, 0.001485275, 0.008472157, 0.000498027, 
    2.299804e-06, 0.0597741, 0.009486417, 0.05684638, 0.0211427, 0.07304071, 
    0.108389, 0.04339248, 0.07710439, 0.0253025, 0.01571872, 0.001260093, 
    0.0001586048, 0.05756566, 0.0439472, 0.09970853, 0.03767064, 0.01178364,
  0.0001421599, 0.05679596, 0.1338936, 0.02627104, 0.05718897, 0.04112827, 
    0.04264905, 0.02591437, 0.001500915, 0.04976068, 0.04482277, 0.05310275, 
    0.09194088, 0.02807778, 0.03880347, 0.1647644, 0.04634077, 0.04494421, 
    0.02649009, 0.03148, 0.08633427, 0.04855671, 2.115208e-06, -4.679476e-05, 
    0.202521, 0.1370269, 0.04382078, 0.0901759, 0.008260047,
  -4.211903e-06, -0.0007283363, 0.2771317, 0.05528478, 0.0494577, 0.03911525, 
    0.05043299, 0.06015977, 0.02667129, 0.02916943, 0.04522968, 0.01583361, 
    0.04327498, 0.01832644, 0.02911687, 0.07139684, 0.06723896, 0.04018364, 
    0.02857724, 0.01264658, 0.002995372, 0.0004822866, 0.0001653952, 
    0.04776086, 0.1395101, 0.07828011, 0.04567778, 0.006522676, 0.004317832,
  0.006332991, 0.004880682, 0.01221811, 0.0301642, 0.0417003, 0.03558252, 
    0.06737297, 0.02430011, 0.19078, 0.2086815, 0.01388099, 0.009501141, 
    0.03131709, 0.0214562, 0.02924204, 0.02255961, 0.0170769, 0.01023107, 
    0.02237833, 0.02817751, 0.02435454, 0.02980213, 0.06096218, 0.0448706, 
    0.1077352, 0.1353157, 0.04663302, 0.02639457, 0.004872195,
  3.759855e-08, 1.551248e-07, 1.430164e-07, 0.01368901, 0.01803458, 
    0.08733496, 0.01634187, 0.07047705, 0.03908084, 0.1150449, 0.2694783, 
    0.09731986, 0.05484786, 0.04181345, 0.02702902, 0.04135961, 0.027992, 
    0.02040317, 0.0319064, 0.04984652, 0.05422145, 0.03631212, 0.08209515, 
    0.02715402, 0.03248917, 0.002378591, 0.0007226223, -8.314589e-07, 
    -2.036266e-05,
  2.40621e-06, 3.88552e-07, 5.640755e-08, 0.01644387, 1.084467e-05, 
    0.009513328, 0.02039642, 0.03913593, 0.02817575, 0.02708789, 0.05333598, 
    0.04568519, 0.07373923, 0.003195951, 0.01993499, 0.01112584, 0.02461, 
    0.02418137, 0.0008932253, 0.005284851, 0.01111784, 0.1601889, 0.06401887, 
    0.1176284, 0.02761544, 0.04699533, 0.02773507, 0.0001791668, 1.249788e-06,
  0.02226583, 0.01053636, 0.01731959, 0.01852603, 0.05189772, 0.02807305, 
    0.00912373, 0.02187042, 0.1024486, 0.06362742, 0.05052066, 0.1796602, 
    0.1313923, 0.144619, 0.1160499, 0.166541, 0.1105043, 0.08484703, 
    0.0716813, 0.01553981, 0.01675997, 0.07949863, 0.05872276, 0.1136638, 
    0.119853, 0.1195255, 0.09012584, 0.05036157, 0.009114992,
  0.06441274, 0.1291702, 0.1805741, 0.3743854, 0.1627304, 0.04078829, 
    0.3343402, 0.01155502, 0.005004951, 0.01135059, 0.06683245, 0.2029007, 
    0.2106549, 0.2258206, 0.2555124, 0.2722916, 0.2406399, 0.2310246, 
    0.1923427, 0.2250698, 0.1617733, 0.05199807, 0.1442494, 0.1339039, 
    0.2320676, 0.1690468, 0.1590096, 0.09011475, 0.1709057,
  0.2193098, 0.2228283, 0.1992892, 0.2077666, 0.184582, 0.1935767, 
    0.08006436, 0.1090179, 0.08511852, 0.03745291, 0.06954658, 0.1880044, 
    0.2077563, 0.3365152, 0.3188883, 0.1706173, 0.1378565, 0.1793521, 
    0.1575422, 0.2372486, 0.08747976, 0.1884078, 0.2597627, 0.2441292, 
    0.2539336, 0.1894117, 0.2455828, 0.2188038, 0.1854477,
  0.3072751, 0.211402, 0.1927468, 0.3635921, 0.3670721, 0.3652014, 0.3879783, 
    0.3163702, 0.287548, 0.2947325, 0.2853163, 0.1725142, 0.2105033, 
    0.2302249, 0.2086989, 0.07118397, 0.166413, 0.3597967, 0.3046926, 
    0.1406387, 0.1744971, 0.1394603, 0.1791667, 0.1845822, 0.1609966, 
    0.3559485, 0.3075174, 0.3604655, 0.2681212,
  0.2696948, 0.3523493, 0.3245989, 0.3600355, 0.286824, 0.4135352, 0.3920092, 
    0.4883317, 0.2754633, 0.2566983, 0.2991201, 0.390192, 0.3735701, 
    0.2548559, 0.3570318, 0.1716896, 0.2510634, 0.4606549, 0.3039207, 
    0.294843, 0.3210998, 0.2225163, 0.3124824, 0.1493931, 0.2283441, 
    0.5084056, 0.1171582, 0.1776997, 0.2036234,
  0.2486571, 0.2271812, 0.2486868, 0.1365547, 0.2162237, 0.2593516, 
    0.2065339, 0.1790071, 0.1918554, 0.2284798, 0.2597321, 0.271371, 
    0.2976811, 0.3283517, 0.400268, 0.4429399, 0.3346428, 0.178652, 
    0.2206397, 0.23385, 0.252023, 0.2482471, 0.1739817, 0.1208564, 0.1424779, 
    0.1061263, 0.1156242, 0.2200361, 0.3427826,
  0.1310529, 0.1308487, 0.1306445, 0.1304403, 0.1302361, 0.1300319, 
    0.1298277, 0.1308679, 0.1285792, 0.1262905, 0.1240018, 0.121713, 
    0.1194243, 0.1171356, 0.1362837, 0.1375724, 0.1388611, 0.1401498, 
    0.1414385, 0.1427272, 0.144016, 0.1503088, 0.1515131, 0.1527173, 
    0.1539215, 0.1551257, 0.1563299, 0.1575341, 0.1312163,
  0.2460021, 0.2085861, 0.2690362, 0.2810227, 0.1819723, 0.1634298, 0.301962, 
    0.3009206, 0.08786773, 0.1966633, 0.1875734, 0.1508344, 0.294888, 
    0.1002036, 0.101874, 0.2319968, 0.2221416, 0.1605268, 0.2441931, 
    0.282184, 0.3277703, 0.2160326, 0.1017661, 0.04778757, 0.04369852, 
    0.04549122, 0.05058902, 0.07420711, 0.1877344,
  0.1875151, 0.2100673, 0.1619253, 0.1267122, 0.2514237, 0.3296548, 
    0.1003696, 0.1663229, 0.1462205, 0.1995394, 0.2199916, 0.1646573, 
    0.2602389, 0.3020382, 0.2652367, 0.2174295, 0.2059786, 0.2803045, 
    0.3405438, 0.2815526, 0.1928925, 0.1440001, 0.2780828, 0.2473156, 
    0.2059061, 0.2321879, 0.2866766, 0.3074911, 0.2259366,
  0.3619404, 0.3609481, 0.3892934, 0.35711, 0.3758633, 0.4555425, 0.3492899, 
    0.3358404, 0.436995, 0.3823101, 0.4370606, 0.3301649, 0.2447374, 
    0.2550844, 0.2493668, 0.3180465, 0.3012486, 0.2797775, 0.2579541, 
    0.2517374, 0.2845407, 0.3429684, 0.3184243, 0.2979689, 0.251505, 
    0.2339467, 0.2152859, 0.2809868, 0.3417706,
  0.2609493, 0.2277685, 0.2391277, 0.2282597, 0.2771439, 0.2568834, 
    0.2623994, 0.3394413, 0.2773866, 0.2559825, 0.2351547, 0.2594872, 
    0.2865249, 0.284651, 0.2372888, 0.1828423, 0.1756741, 0.1605552, 
    0.1768014, 0.1825623, 0.2238032, 0.2797329, 0.312027, 0.1849412, 
    0.1101932, 0.1069298, 0.1808668, 0.1831805, 0.2304135,
  0.07745003, 0.1023381, 0.1276748, 0.1048781, 0.1449788, 0.08370881, 
    0.1356002, 0.119109, 0.1445866, 0.05968766, 0.02939973, 0.009329961, 
    0.06805503, 0.04936933, 0.0981294, 0.0984447, 0.1580049, 0.09567139, 
    0.1231246, 0.1563338, 0.112135, 0.07078043, 0.1060831, 0.06990676, 
    0.01186582, 0.04854891, 0.1669726, 0.09410837, 0.09820535,
  0.02284521, 0.0528959, 0.09830191, 0.08364065, 0.02994076, 0.05869976, 
    0.0395895, 0.02457421, 0.005315172, 0.005203024, 0.0002125866, 
    4.289359e-07, 0.0466246, 0.01681109, 0.06467014, 0.0465357, 0.09343684, 
    0.1108958, 0.04125516, 0.07073643, 0.02575544, 0.05345071, 0.02052855, 
    6.646105e-05, 0.06991421, 0.07112034, 0.08586653, 0.03282912, 0.03278213,
  0.007105337, 0.0394016, 0.1321707, 0.02767964, 0.04563616, 0.03624431, 
    0.04072789, 0.03771627, 0.002187595, 0.05748207, 0.03688154, 0.0534563, 
    0.09004236, 0.02562107, 0.04471911, 0.1652417, 0.04190202, 0.03454655, 
    0.02222386, 0.0256338, 0.04746164, 0.1584684, 0.001812647, 0.0002576082, 
    0.2170575, 0.1298034, 0.03206086, 0.08655613, 0.07484657,
  -9.004741e-05, -0.0005025662, 0.2404401, 0.04947473, 0.04208925, 
    0.03484713, 0.04593901, 0.05767897, 0.03059311, 0.02665978, 0.06627182, 
    0.01538702, 0.04408855, 0.01863809, 0.02496295, 0.05197892, 0.05638541, 
    0.03394806, 0.03044934, 0.03399865, 0.01976602, 0.003165436, 
    0.0004489346, 0.05074095, 0.1125129, 0.06858118, 0.05113796, 0.01514331, 
    0.01830506,
  0.00539513, 0.006889487, 0.0141087, 0.01853496, 0.0428468, 0.03504593, 
    0.05190741, 0.0187997, 0.2113511, 0.2291917, 0.01737369, 0.01163253, 
    0.02659081, 0.01993563, 0.02810486, 0.02456346, 0.02064952, 0.01082584, 
    0.02264673, 0.03715491, 0.04016249, 0.04763138, 0.05127601, 0.04017159, 
    0.1136614, 0.1139984, 0.03807551, 0.02302193, 0.003656972,
  1.484937e-08, 4.498743e-08, 6.602752e-08, 0.002197226, 0.05162653, 
    0.08427268, 0.02269361, 0.05829631, 0.04758082, 0.1196967, 0.2672401, 
    0.08251856, 0.06090849, 0.0485153, 0.03682892, 0.04027856, 0.02674074, 
    0.02650524, 0.03770233, 0.04704285, 0.05411785, 0.03349467, 0.1159063, 
    0.03546577, 0.03008124, 0.007914863, 0.001392515, -8.21799e-07, 
    -1.321854e-05,
  1.421697e-06, 3.208953e-07, 2.790843e-08, 0.02226071, 2.6271e-07, 
    0.07252191, 0.04588786, 0.02996309, 0.06914799, 0.1292797, 0.08291174, 
    0.1011164, 0.08855025, 0.0335312, 0.04506121, 0.02642088, 0.03163001, 
    0.0276104, 0.01280034, 0.01021601, 0.006750012, 0.1764825, 0.06971647, 
    0.1482198, 0.02454213, 0.04190267, 0.06461685, 0.005260674, 1.468375e-06,
  0.005154419, 0.01137745, 0.04170678, 0.01319764, 0.05117275, 0.02190455, 
    0.02702668, 0.01479044, 0.08497546, 0.04491535, 0.2134188, 0.2447195, 
    0.1675903, 0.1609526, 0.1512438, 0.1766336, 0.1338115, 0.1032702, 
    0.07160679, 0.02109098, 0.01424347, 0.1026012, 0.05466356, 0.1569555, 
    0.1459688, 0.1159206, 0.09414771, 0.0647196, 0.01068871,
  0.05913744, 0.1413503, 0.1809293, 0.383317, 0.1621432, 0.03682877, 
    0.2829729, 0.01082232, 0.002192563, 0.009656967, 0.06029705, 0.283741, 
    0.2500641, 0.2666047, 0.2692404, 0.2856017, 0.2574417, 0.2463323, 
    0.2417173, 0.2644973, 0.1613331, 0.07090151, 0.1759755, 0.1470078, 
    0.2325132, 0.1752395, 0.1772654, 0.1214388, 0.2004051,
  0.2912845, 0.2723061, 0.1772375, 0.2179951, 0.1809047, 0.2292076, 
    0.09612434, 0.1314127, 0.08346041, 0.02948251, 0.0753231, 0.2106043, 
    0.2314288, 0.4297281, 0.3722624, 0.2771827, 0.2162032, 0.2473006, 
    0.2315814, 0.2392157, 0.09474282, 0.2055095, 0.2715696, 0.2745574, 
    0.2487632, 0.2616085, 0.3151134, 0.2319929, 0.2201003,
  0.3363743, 0.189413, 0.2148678, 0.3328251, 0.380845, 0.3483649, 0.4436247, 
    0.3614317, 0.2981115, 0.3152677, 0.3106051, 0.1569728, 0.2090092, 
    0.2487538, 0.2280023, 0.05960211, 0.1722601, 0.3668022, 0.2989102, 
    0.1419258, 0.1899688, 0.1777531, 0.1828778, 0.1559703, 0.2197829, 
    0.3324255, 0.2866092, 0.3847631, 0.2827188,
  0.4025725, 0.3164278, 0.3331999, 0.3462135, 0.3234758, 0.432528, 0.4386351, 
    0.5281458, 0.31554, 0.2914191, 0.3061859, 0.386903, 0.354624, 0.2831423, 
    0.4064571, 0.1911178, 0.3203191, 0.5103765, 0.3282816, 0.2636147, 
    0.3082736, 0.2372774, 0.3088672, 0.1169151, 0.219733, 0.5560444, 
    0.1185386, 0.1621686, 0.3371703,
  0.2562349, 0.2072667, 0.3019622, 0.2013153, 0.2236411, 0.2843014, 
    0.2479368, 0.2402373, 0.2471581, 0.2310235, 0.2591391, 0.2977021, 
    0.3207761, 0.3504846, 0.4271715, 0.4260789, 0.3573124, 0.1774852, 
    0.255657, 0.2922522, 0.2611153, 0.2520796, 0.1916311, 0.1246198, 
    0.1359864, 0.1465274, 0.1162359, 0.2617254, 0.405911,
  0.1995048, 0.2002687, 0.2010326, 0.2017965, 0.2025604, 0.2033243, 
    0.2040882, 0.2046532, 0.1986643, 0.1926755, 0.1866866, 0.1806977, 
    0.1747088, 0.1687199, 0.140226, 0.1404159, 0.1406058, 0.1407957, 
    0.1409857, 0.1411756, 0.1413655, 0.1552067, 0.1602418, 0.1652768, 
    0.1703119, 0.175347, 0.1803821, 0.1854172, 0.1988937,
  0.2216481, 0.2018702, 0.2308922, 0.2634928, 0.1878555, 0.1879734, 
    0.3026508, 0.2915793, 0.09667979, 0.1810428, 0.2313359, 0.1555051, 
    0.2966634, 0.1039944, 0.1306864, 0.2574723, 0.2678067, 0.2400794, 
    0.2287855, 0.2679854, 0.3223388, 0.2742341, 0.1415672, 0.1194799, 
    0.1809281, 0.0763047, 0.171791, 0.1532283, 0.193707,
  0.1875753, 0.2028724, 0.1536219, 0.1110265, 0.239708, 0.3677318, 
    0.06892183, 0.173371, 0.1624527, 0.2029787, 0.1982952, 0.1786337, 
    0.2437088, 0.2911052, 0.291094, 0.2294358, 0.32029, 0.4348457, 0.3280671, 
    0.2812092, 0.1838794, 0.1967467, 0.3786414, 0.2850615, 0.2622093, 
    0.30099, 0.336396, 0.4293032, 0.3030625,
  0.4336515, 0.3842433, 0.4095671, 0.4278751, 0.4042864, 0.485449, 0.4439571, 
    0.3691804, 0.4696276, 0.3877984, 0.4597009, 0.4334136, 0.3769597, 
    0.3666399, 0.3471365, 0.3571632, 0.367207, 0.3485362, 0.3281073, 
    0.3728098, 0.3620183, 0.407628, 0.4417522, 0.3852984, 0.3591371, 
    0.3434372, 0.2888699, 0.3608395, 0.4493523,
  0.3086489, 0.2787368, 0.2839527, 0.2810853, 0.339397, 0.2859019, 0.3064543, 
    0.382822, 0.2885398, 0.305873, 0.2886828, 0.3249811, 0.3309109, 
    0.3284157, 0.2200003, 0.1766986, 0.1966223, 0.1870978, 0.1908649, 
    0.2064243, 0.2626712, 0.2998138, 0.3394822, 0.1798871, 0.09402486, 
    0.1065629, 0.228617, 0.2454199, 0.2599654,
  0.11826, 0.1470281, 0.2219453, 0.182639, 0.1739335, 0.1366484, 0.1924449, 
    0.1566104, 0.1838885, 0.08998088, 0.07666086, 0.05856391, 0.08733992, 
    0.101294, 0.1263844, 0.09182199, 0.1920207, 0.1423481, 0.200241, 
    0.1839546, 0.149359, 0.1459471, 0.1496772, 0.09839984, 0.0168581, 
    0.08945667, 0.218832, 0.1431641, 0.1278486,
  0.1282176, 0.04147675, 0.1049786, 0.1185676, 0.03175991, 0.08462676, 
    0.06809225, 0.07465226, 0.0594814, 0.00530202, 6.625086e-05, 
    -1.958702e-08, 0.03986695, 0.0281673, 0.1073204, 0.09153199, 0.1448416, 
    0.1209634, 0.05734888, 0.06098973, 0.0270406, 0.09585252, 0.08280768, 
    2.952625e-05, 0.09422668, 0.07089272, 0.08794278, 0.03274884, 0.08280883,
  0.1388806, 0.0233215, 0.1178137, 0.03083032, 0.04141149, 0.03862963, 
    0.04628284, 0.05962095, 0.02993659, 0.05946019, 0.04576477, 0.04499035, 
    0.08699474, 0.02397315, 0.04764671, 0.1617091, 0.03917208, 0.02754298, 
    0.02330585, 0.03053606, 0.03345357, 0.1258153, 0.0737633, 0.0003509829, 
    0.2494459, 0.1376983, 0.03177191, 0.08014005, 0.152821,
  0.004638018, 0.0006858617, 0.2056427, 0.04999726, 0.03385993, 0.03374796, 
    0.04313644, 0.04960829, 0.03561407, 0.03117814, 0.06844512, 0.02056284, 
    0.04551873, 0.02224243, 0.02357462, 0.04657171, 0.05206561, 0.03190214, 
    0.02921336, 0.03002452, 0.03488157, 0.01610037, 0.009075479, 0.04823405, 
    0.09136482, 0.0665382, 0.05566537, 0.03551273, 0.03409361,
  0.005689632, 0.01777516, 0.007316018, 0.0158849, 0.04392878, 0.03328026, 
    0.04302459, 0.02031094, 0.1978713, 0.2173119, 0.02559004, 0.0132936, 
    0.02379707, 0.02064005, 0.03092805, 0.02793503, 0.0213544, 0.01322296, 
    0.0246885, 0.03302836, 0.0397049, 0.0427833, 0.04359015, 0.04323416, 
    0.1217997, 0.09303566, 0.03319357, 0.02498094, 0.004570853,
  9.307811e-09, 1.866843e-08, 2.28949e-08, 6.136048e-05, 0.1060214, 
    0.08582816, 0.02930011, 0.06552796, 0.08630162, 0.1083793, 0.2407449, 
    0.07147458, 0.05531473, 0.04574302, 0.03827086, 0.04124858, 0.02586532, 
    0.03448992, 0.04668284, 0.04353217, 0.05276118, 0.03775206, 0.1283722, 
    0.05237851, 0.03758062, 0.02210968, 0.008297832, -5.841642e-07, 
    -6.637466e-06,
  7.260832e-07, 1.464096e-07, 1.368544e-08, 0.01499341, -1.745971e-07, 
    0.08922529, 0.05602962, 0.08432768, 0.04295143, 0.1565669, 0.2264773, 
    0.1992551, 0.1461416, 0.1005842, 0.1512077, 0.125199, 0.04783497, 
    0.02550605, 0.03659205, 0.04359204, 0.0100876, 0.2154824, 0.122401, 
    0.1390667, 0.05748865, 0.07979356, 0.09854215, 0.01746788, 7.134017e-07,
  0.007629942, 0.0247012, 0.07772559, 0.01477306, 0.06357982, 0.01778468, 
    0.02474836, 0.008660826, 0.06011481, 0.05528627, 0.4495324, 0.1468237, 
    0.1157176, 0.1743468, 0.1405679, 0.1590812, 0.1507621, 0.1625582, 
    0.1121744, 0.04671226, 0.01349287, 0.1137262, 0.05212423, 0.1097797, 
    0.1262941, 0.1667676, 0.1003303, 0.093133, 0.01247944,
  0.05145815, 0.1501566, 0.2050445, 0.3853393, 0.1649804, 0.05637053, 
    0.2430568, 0.01103295, 0.0009519162, 0.008382203, 0.07165598, 0.4090267, 
    0.3114821, 0.258456, 0.2547193, 0.2819381, 0.2758375, 0.2668624, 
    0.285782, 0.309413, 0.1664424, 0.07025734, 0.2121549, 0.1787701, 
    0.2713383, 0.1811258, 0.189675, 0.1902675, 0.2425585,
  0.3194087, 0.3271007, 0.2079431, 0.293083, 0.2284231, 0.3263941, 
    0.07851982, 0.1398188, 0.07810724, 0.02253738, 0.08426299, 0.234262, 
    0.3565286, 0.4693539, 0.3592363, 0.2955433, 0.3253807, 0.3307567, 
    0.2596527, 0.2653035, 0.1138231, 0.2479513, 0.2944427, 0.2863562, 
    0.2720791, 0.3339297, 0.3615846, 0.2507426, 0.2543002,
  0.3549249, 0.200889, 0.2029994, 0.3225562, 0.3747414, 0.3419793, 0.4826836, 
    0.418251, 0.3376652, 0.368281, 0.3278761, 0.1593769, 0.2135024, 
    0.2651991, 0.3863358, 0.08504308, 0.2406662, 0.3872575, 0.3151807, 
    0.1512228, 0.2144085, 0.1761227, 0.1765448, 0.1319795, 0.3219536, 
    0.3129217, 0.3052698, 0.3609359, 0.3239771,
  0.3828876, 0.2601709, 0.3586147, 0.376907, 0.3649846, 0.4498712, 0.4625722, 
    0.5616986, 0.3516575, 0.3398775, 0.327141, 0.3845271, 0.3396532, 
    0.3012413, 0.4431954, 0.2052606, 0.3760836, 0.5739313, 0.3343596, 
    0.2804588, 0.3120451, 0.2462378, 0.2897617, 0.1147704, 0.2156683, 
    0.5616366, 0.1222026, 0.136911, 0.4379399,
  0.2660161, 0.2121129, 0.340012, 0.2179483, 0.2498117, 0.3279023, 0.2940344, 
    0.2790894, 0.3055176, 0.2842199, 0.2901028, 0.337524, 0.3523771, 
    0.3998347, 0.4944645, 0.4546115, 0.3578491, 0.1806231, 0.2458719, 
    0.3682429, 0.283845, 0.2826722, 0.1931631, 0.1306992, 0.139603, 
    0.1784032, 0.1243482, 0.2862576, 0.4171298,
  0.2625196, 0.2618038, 0.261088, 0.2603721, 0.2596563, 0.2589405, 0.2582246, 
    0.2521561, 0.2463469, 0.2405377, 0.2347285, 0.2289193, 0.2231101, 
    0.2173009, 0.1863643, 0.1867068, 0.1870493, 0.1873918, 0.1877343, 
    0.1880769, 0.1884194, 0.1804279, 0.1866104, 0.1927929, 0.1989754, 
    0.2051579, 0.2113404, 0.2175229, 0.2630922,
  0.2523988, 0.2091967, 0.2381832, 0.25733, 0.1606745, 0.1886688, 0.2644289, 
    0.2559236, 0.1149759, 0.2223846, 0.2485604, 0.182742, 0.3266189, 
    0.08964215, 0.1866874, 0.280392, 0.2468593, 0.2163713, 0.2353761, 
    0.2559859, 0.3213358, 0.2978739, 0.1910852, 0.1175157, 0.2330979, 
    0.1612967, 0.1483033, 0.2309715, 0.2698172,
  0.2589997, 0.2101701, 0.1501796, 0.09657989, 0.2324667, 0.4289099, 
    0.03963409, 0.1735557, 0.1824073, 0.2003998, 0.2123661, 0.2198727, 
    0.2063552, 0.2804565, 0.3599419, 0.3604015, 0.4057179, 0.466009, 
    0.3163113, 0.3677478, 0.312644, 0.3571192, 0.4740551, 0.2977772, 
    0.3080544, 0.4141665, 0.5309566, 0.4611161, 0.3953823,
  0.4551875, 0.3913895, 0.4634894, 0.5235822, 0.4806491, 0.5318726, 
    0.4792022, 0.4674684, 0.5143766, 0.3873864, 0.4899859, 0.5096467, 
    0.4641837, 0.4865096, 0.4023675, 0.4000113, 0.4069861, 0.4012025, 
    0.4221686, 0.4089468, 0.4466256, 0.4601866, 0.4915329, 0.4328077, 
    0.4373053, 0.4597723, 0.3429427, 0.4148513, 0.4708834,
  0.3695188, 0.3449558, 0.3924462, 0.3428927, 0.3589343, 0.3204493, 
    0.3569766, 0.3834415, 0.3216559, 0.3975204, 0.3877639, 0.3202251, 
    0.3372384, 0.2891459, 0.1579197, 0.1421571, 0.2036764, 0.2273645, 
    0.2693425, 0.2609936, 0.3178709, 0.332584, 0.3494479, 0.1719729, 
    0.06704259, 0.1279251, 0.2832686, 0.3170666, 0.2844431,
  0.1680663, 0.2161856, 0.2536867, 0.2387963, 0.2200974, 0.2526653, 
    0.2069113, 0.18197, 0.2900761, 0.1636783, 0.2133748, 0.1178705, 
    0.09911139, 0.1283782, 0.1509322, 0.1556178, 0.2880684, 0.2681296, 
    0.2279395, 0.2499959, 0.1407569, 0.1950143, 0.1917011, 0.1280906, 
    0.0327929, 0.1059138, 0.2866665, 0.2013575, 0.2160484,
  0.1731411, 0.04268733, 0.1041873, 0.1293735, 0.0344722, 0.08170981, 
    0.151758, 0.215579, 0.2744507, 0.01536164, -2.372679e-05, 1.15022e-07, 
    0.03102423, 0.04533226, 0.1860203, 0.1339517, 0.2453328, 0.1817056, 
    0.1238367, 0.07088318, 0.03674026, 0.1079149, 0.211522, 6.264533e-05, 
    0.08382221, 0.1247408, 0.09756672, 0.03826113, 0.1383593,
  0.2960837, 0.01940953, 0.0893859, 0.04197602, 0.04679263, 0.05043763, 
    0.05884515, 0.06606643, 0.1351711, 0.06885564, 0.04168356, 0.03072766, 
    0.0976343, 0.0512916, 0.07352769, 0.145426, 0.04510574, 0.03099389, 
    0.03096764, 0.04291625, 0.04283357, 0.1260256, 0.5146338, 0.001419058, 
    0.2410083, 0.1471069, 0.04493601, 0.06431413, 0.1467575,
  0.032865, 0.005896134, 0.1708391, 0.06073595, 0.03323831, 0.03552391, 
    0.04280319, 0.04720191, 0.04392818, 0.03894596, 0.05374117, 0.03481106, 
    0.04452226, 0.03114675, 0.02928992, 0.04977841, 0.08669493, 0.03876654, 
    0.03871289, 0.04963943, 0.06572095, 0.05879017, 0.04418593, 0.03988478, 
    0.0736696, 0.04563664, 0.09977623, 0.07149292, 0.07000779,
  0.008831084, 0.006048754, 0.001979727, 0.01130238, 0.05353843, 0.03894222, 
    0.04503448, 0.02461113, 0.1786188, 0.1766517, 0.02844291, 0.01723172, 
    0.02816069, 0.02629413, 0.04191, 0.03997657, 0.02923547, 0.024111, 
    0.02511233, 0.03385018, 0.04233634, 0.03543313, 0.04427146, 0.03601632, 
    0.110238, 0.07859974, 0.03643094, 0.0321708, 0.02495668,
  6.937231e-09, 9.659462e-09, 6.881985e-09, -0.0007893678, 0.1365093, 
    0.1477126, 0.01145778, 0.1387632, 0.1336518, 0.09475777, 0.22176, 
    0.06910458, 0.0503541, 0.06321144, 0.06111987, 0.08286534, 0.06388951, 
    0.04730874, 0.05672761, 0.05232568, 0.05431683, 0.06388703, 0.1691549, 
    0.05949688, 0.06700171, 0.07062572, 0.1641359, -1.16946e-07, -4.223918e-06,
  3.166984e-07, 3.96409e-08, -1.900611e-08, 0.02125677, 4.276432e-08, 
    0.07934602, 0.03340694, 0.0776595, 0.04889382, 0.2308746, 0.2140636, 
    0.2198969, 0.2016553, 0.1764665, 0.1258636, 0.1254717, 0.1463975, 
    0.04668238, 0.0781177, 0.1142811, 0.02325128, 0.2538729, 0.1871466, 
    0.1499919, 0.110022, 0.0779586, 0.08482887, 0.01563088, 3.901585e-07,
  0.00840342, 0.03909434, 0.03235152, 0.03115461, 0.07652684, 0.01567067, 
    0.01053951, 0.006011958, 0.04245511, 0.07016809, 0.2479982, 0.06043729, 
    0.06518253, 0.1168218, 0.1042754, 0.1324016, 0.1031139, 0.1646439, 
    0.1241172, 0.09119352, 0.01807759, 0.1161107, 0.06498989, 0.06176715, 
    0.0836316, 0.1410825, 0.1366237, 0.114869, 0.01470691,
  0.03699039, 0.1530041, 0.2149206, 0.3872949, 0.1583387, 0.05530138, 
    0.2087221, 0.01039267, 0.0009547694, 0.01009879, 0.08784256, 0.3447546, 
    0.2474699, 0.191888, 0.22307, 0.2609859, 0.2780896, 0.3115685, 0.2678473, 
    0.3524918, 0.1733821, 0.09458601, 0.2481678, 0.2254453, 0.3044326, 
    0.2043596, 0.150753, 0.2305691, 0.2592864,
  0.3494912, 0.3426641, 0.2549901, 0.3113468, 0.2577687, 0.3814569, 
    0.1086209, 0.1366291, 0.07043118, 0.02053882, 0.08913594, 0.2766395, 
    0.4708861, 0.4220438, 0.3381466, 0.2560202, 0.3443203, 0.2902449, 
    0.2195646, 0.294288, 0.1220804, 0.2821752, 0.308603, 0.3035246, 
    0.2971759, 0.3383284, 0.3065118, 0.2757098, 0.3230333,
  0.2866969, 0.1463301, 0.2437181, 0.4175604, 0.440059, 0.3362184, 0.4805897, 
    0.4365402, 0.3732276, 0.4162011, 0.4033056, 0.1675427, 0.2158112, 
    0.2545813, 0.5405907, 0.1992242, 0.3028055, 0.3897968, 0.3582526, 
    0.1919764, 0.2223623, 0.1648252, 0.1822775, 0.1130974, 0.5268399, 
    0.2241086, 0.2982176, 0.3038398, 0.2492719,
  0.2801118, 0.1534043, 0.3048783, 0.327723, 0.3943841, 0.4896518, 0.4805968, 
    0.5826818, 0.3657389, 0.4125363, 0.3729678, 0.3959574, 0.3675935, 
    0.325161, 0.4469154, 0.2163048, 0.4202483, 0.6071155, 0.3303706, 
    0.3637745, 0.3310622, 0.2495559, 0.2842754, 0.1198129, 0.20143, 0.585701, 
    0.1242769, 0.1079452, 0.4533389,
  0.2463699, 0.2252677, 0.3443794, 0.2123538, 0.2527085, 0.3467361, 
    0.3679762, 0.3686228, 0.3418585, 0.3392485, 0.3339962, 0.3720763, 
    0.377695, 0.482765, 0.5262405, 0.4848337, 0.3679845, 0.2003698, 
    0.2789097, 0.3864576, 0.3433209, 0.2898632, 0.2179433, 0.1399217, 
    0.1464671, 0.2133223, 0.1260678, 0.2879007, 0.3948085,
  0.255346, 0.2593552, 0.2633644, 0.2673737, 0.2713829, 0.2753921, 0.2794014, 
    0.289465, 0.2814697, 0.2734745, 0.2654792, 0.257484, 0.2494887, 
    0.2414934, 0.2239514, 0.2229218, 0.2218921, 0.2208625, 0.2198328, 
    0.2188032, 0.2177735, 0.1967918, 0.2018075, 0.2068231, 0.2118388, 
    0.2168545, 0.2218701, 0.2268858, 0.2521386,
  0.2741496, 0.2189191, 0.2742016, 0.244502, 0.1331853, 0.1848973, 0.239039, 
    0.2016865, 0.1114881, 0.3063394, 0.2991833, 0.2514887, 0.3785217, 
    0.05811419, 0.1879088, 0.3118738, 0.2740824, 0.3031078, 0.2518331, 
    0.2757216, 0.3614895, 0.3449896, 0.1696657, 0.08233459, 0.1151562, 
    0.3543113, 0.1600054, 0.1582858, 0.2358488,
  0.2618141, 0.3482399, 0.1991889, 0.1240926, 0.1813735, 0.45998, 0.03242227, 
    0.1571543, 0.1675165, 0.2086913, 0.2606503, 0.2523552, 0.1620665, 
    0.3436438, 0.5239218, 0.5634452, 0.5040992, 0.5043615, 0.3715831, 
    0.3668555, 0.3833048, 0.3674154, 0.4247718, 0.318158, 0.2982216, 
    0.4624692, 0.5172659, 0.4602084, 0.3727222,
  0.4709201, 0.4139944, 0.4761175, 0.5433463, 0.589334, 0.6127769, 0.4798857, 
    0.4897821, 0.5612097, 0.4207302, 0.4645746, 0.5489247, 0.4978903, 
    0.4410179, 0.4167241, 0.4879982, 0.4879194, 0.4756784, 0.5231514, 
    0.4758236, 0.4440089, 0.443245, 0.4022975, 0.3930329, 0.4701847, 
    0.516596, 0.4621259, 0.4971608, 0.5647114,
  0.3953996, 0.3750406, 0.4737258, 0.3585928, 0.4281541, 0.373004, 0.3704463, 
    0.3530533, 0.3402242, 0.3873705, 0.3853695, 0.3304664, 0.2596729, 
    0.241556, 0.138997, 0.109154, 0.2529507, 0.2810826, 0.3078259, 0.2784826, 
    0.4284177, 0.3798611, 0.3307175, 0.1708809, 0.05194467, 0.1247114, 
    0.2919227, 0.3249674, 0.3035058,
  0.2491103, 0.2497704, 0.1824108, 0.2704461, 0.2996509, 0.2699105, 
    0.2100184, 0.2012169, 0.3203167, 0.3361924, 0.3098328, 0.1378798, 
    0.128437, 0.1742902, 0.1752951, 0.1613646, 0.3082659, 0.3731997, 
    0.2527254, 0.3313313, 0.3148164, 0.2478953, 0.1997131, 0.1542292, 
    0.01212528, 0.1557081, 0.2894055, 0.2842253, 0.2494525,
  0.1299684, 0.1369815, 0.07584456, 0.1331479, 0.04940619, 0.09737863, 
    0.1942196, 0.1966713, 0.3625839, 0.02235877, 3.598947e-05, 1.125947e-07, 
    0.03097731, 0.1533428, 0.2143146, 0.08143123, 0.3159508, 0.2884681, 
    0.1971593, 0.1052473, 0.109408, 0.1154512, 0.2572824, 0.0006936262, 
    0.08540919, 0.09023876, 0.08541154, 0.1103697, 0.1295509,
  0.3622233, 0.01830067, 0.06791759, 0.07530416, 0.07066273, 0.04872159, 
    0.04549556, 0.07109073, 0.3768092, 0.1005689, 0.03870437, 0.02148612, 
    0.1018691, 0.08455151, 0.05950824, 0.1409141, 0.09113917, 0.04073515, 
    0.0318372, 0.0259286, 0.03289342, 0.07874142, 0.4875641, 0.008420843, 
    0.2000074, 0.1308204, 0.07238556, 0.03928172, 0.08356227,
  0.1522999, 0.03806369, 0.1284689, 0.06750031, 0.04254419, 0.06157638, 
    0.08825804, 0.07755715, 0.1012186, 0.04714601, 0.03373257, 0.03252931, 
    0.05596132, 0.1257347, 0.1019522, 0.1031012, 0.05269909, 0.05250122, 
    0.05878676, 0.06316877, 0.1158966, 0.2555059, 0.1768139, 0.02441154, 
    0.05875709, 0.02864597, 0.09512226, 0.1342367, 0.1740679,
  0.01491868, 0.002787143, 0.0009732535, 0.008957098, 0.08946723, 0.1227737, 
    0.101644, 0.06532492, 0.1882592, 0.1283326, 0.058982, 0.1252398, 
    0.04571793, 0.05887957, 0.07450037, 0.08221575, 0.04473236, 0.05430382, 
    0.05369313, 0.0769887, 0.1085959, 0.0767796, 0.05071664, 0.01481452, 
    0.07119204, 0.07880663, 0.05628582, 0.09626075, 0.05419208,
  6.00633e-09, 5.777896e-09, 2.208202e-09, -0.001932591, 0.1551285, 
    0.1413161, 0.005289394, 0.09146494, 0.06644434, 0.09567514, 0.1993382, 
    0.08609781, 0.06892154, 0.06488311, 0.0818547, 0.1039482, 0.1011031, 
    0.07888202, 0.09756245, 0.06388746, 0.08165191, 0.08246394, 0.2355358, 
    0.075746, 0.04088221, 0.07475036, 0.1845925, -0.000264908, -1.842266e-06,
  1.234262e-07, 7.226938e-09, -2.647975e-09, 0.01919788, 4.471275e-08, 
    0.01624432, 0.01546984, 0.04644031, 0.02560152, 0.2519119, 0.1016253, 
    0.1315293, 0.1499347, 0.1510027, 0.1117926, 0.0805423, 0.09069397, 
    0.07361802, 0.08320266, 0.2563309, 0.02748483, 0.2548133, 0.1127351, 
    0.1008738, 0.09214814, 0.1070934, 0.08695874, 0.00420795, 1.491416e-07,
  0.001423617, 0.03854327, 0.0106786, 0.03401677, 0.09106094, 0.01047245, 
    0.01426289, 0.006851979, 0.03030161, 0.06544176, 0.1052244, 0.02863875, 
    0.04453665, 0.09311236, 0.07685471, 0.1088602, 0.08398268, 0.1383787, 
    0.1957502, 0.1504186, 0.01880995, 0.1304941, 0.09450222, 0.0400329, 
    0.05422795, 0.1195319, 0.1383078, 0.1616018, 0.01931176,
  0.02282001, 0.1072856, 0.1985568, 0.3834973, 0.1050264, 0.05555611, 
    0.1844288, 0.01070954, 0.0005765, 0.0123208, 0.09347083, 0.1579844, 
    0.1653819, 0.1469125, 0.1833221, 0.2082198, 0.20637, 0.2472782, 
    0.2460154, 0.3713001, 0.1735281, 0.1033174, 0.3001491, 0.2701826, 
    0.2581148, 0.21072, 0.1410263, 0.2057976, 0.2819531,
  0.3367765, 0.3114871, 0.2734732, 0.3121609, 0.289567, 0.3822334, 0.1319125, 
    0.1317423, 0.06216134, 0.03376511, 0.1034878, 0.287757, 0.4279613, 
    0.3504435, 0.3401094, 0.2906224, 0.3552687, 0.2589311, 0.1885286, 
    0.3077173, 0.1411229, 0.321127, 0.3032826, 0.3285531, 0.3336685, 
    0.2667013, 0.3062175, 0.235015, 0.2774768,
  0.2219694, 0.1514359, 0.2421367, 0.4619996, 0.5399821, 0.4007511, 
    0.5407946, 0.4989622, 0.4170618, 0.4599204, 0.4711511, 0.1811972, 
    0.2172213, 0.2423234, 0.5351969, 0.3357097, 0.3324626, 0.4042369, 
    0.4203845, 0.2153635, 0.2715955, 0.2287798, 0.1703551, 0.1027702, 
    0.649685, 0.1520993, 0.2512214, 0.2516448, 0.2079685,
  0.1831849, 0.09917734, 0.2372598, 0.2633487, 0.4239074, 0.4564626, 
    0.5222291, 0.6101581, 0.3625007, 0.4815046, 0.425895, 0.3830083, 
    0.4088071, 0.3589463, 0.4670954, 0.2276067, 0.4513908, 0.618574, 
    0.320729, 0.4416946, 0.3650979, 0.227976, 0.2963223, 0.1305841, 
    0.1825442, 0.5758297, 0.139784, 0.1048002, 0.3168103,
  0.2217967, 0.273375, 0.3452997, 0.2677854, 0.2814087, 0.3963366, 0.4194437, 
    0.394675, 0.3576686, 0.3686048, 0.3687896, 0.4223517, 0.4441392, 
    0.5650255, 0.5294794, 0.5366043, 0.4183416, 0.250537, 0.3157219, 
    0.4390325, 0.4123977, 0.3149433, 0.1973611, 0.1430136, 0.1539441, 
    0.2316247, 0.1366742, 0.2854776, 0.4061148,
  0.2551941, 0.2605655, 0.2659368, 0.2713082, 0.2766795, 0.2820508, 
    0.2874222, 0.3321361, 0.3244289, 0.3167216, 0.3090143, 0.3013071, 
    0.2935998, 0.2858925, 0.2561615, 0.2562808, 0.2564001, 0.2565194, 
    0.2566387, 0.2567579, 0.2568772, 0.2569425, 0.2591591, 0.2613757, 
    0.2635924, 0.265809, 0.2680256, 0.2702422, 0.250897,
  0.2815016, 0.2265071, 0.295856, 0.2965772, 0.1188235, 0.1536029, 0.1963754, 
    0.181691, 0.133719, 0.3074466, 0.387976, 0.2581261, 0.3716767, 
    0.06349557, 0.208549, 0.2871356, 0.2270754, 0.2081237, 0.2402116, 
    0.1684249, 0.2861705, 0.3862461, 0.153684, 0.0588212, 0.1104776, 
    0.2484111, 0.2296383, 0.1088974, 0.1924638,
  0.2379006, 0.3026634, 0.2675447, 0.1164611, 0.1224446, 0.3962608, 
    0.0297077, 0.1009693, 0.1115295, 0.1658609, 0.2570006, 0.2648924, 
    0.1028499, 0.3132188, 0.5821581, 0.5314795, 0.4635668, 0.4994892, 
    0.405643, 0.4748991, 0.3877406, 0.4640248, 0.5275506, 0.3349102, 
    0.3089278, 0.3785092, 0.4566244, 0.3517823, 0.3107212,
  0.5271766, 0.4438048, 0.4389647, 0.4711809, 0.5736684, 0.6216266, 0.469186, 
    0.4220151, 0.5380893, 0.4214417, 0.4554735, 0.5071119, 0.4770258, 
    0.384515, 0.3970254, 0.5064864, 0.5823851, 0.5339032, 0.5610372, 
    0.4987693, 0.3931015, 0.4107128, 0.3313428, 0.3600154, 0.4635561, 
    0.4895949, 0.4992781, 0.4755083, 0.5203054,
  0.4040743, 0.3527558, 0.4423089, 0.3560558, 0.4629834, 0.3660648, 
    0.3606634, 0.3067915, 0.3510368, 0.3676181, 0.3451355, 0.2875794, 
    0.2304644, 0.2301376, 0.1412753, 0.1251276, 0.2926124, 0.3614657, 
    0.3709431, 0.363633, 0.4614191, 0.3646491, 0.3015755, 0.1750925, 
    0.04320293, 0.1343778, 0.3018459, 0.3280457, 0.3706479,
  0.1797268, 0.1576868, 0.1206802, 0.1869677, 0.2859562, 0.2624135, 0.229794, 
    0.1879299, 0.2298424, 0.2336976, 0.2494345, 0.08885959, 0.08435747, 
    0.1383213, 0.1905229, 0.1871686, 0.2591366, 0.2985209, 0.2946378, 
    0.287564, 0.3074779, 0.2302863, 0.1403653, 0.1876559, 0.008450813, 
    0.1940094, 0.2902223, 0.3067389, 0.207703,
  0.06161965, 0.06421979, 0.06152366, 0.1170319, 0.0952957, 0.07653882, 
    0.06933057, 0.08211511, 0.1617539, 0.02426521, -1.721944e-05, 
    4.871661e-08, 0.03126129, 0.1502842, 0.1219314, 0.05457298, 0.2391544, 
    0.3034111, 0.1572962, 0.08527321, 0.09772532, 0.02748834, 0.08945979, 
    0.02483547, 0.08018114, 0.06550501, 0.09643263, 0.07249856, 0.07225145,
  0.1506696, 0.03569414, 0.0438962, 0.07799407, 0.02720403, 0.01213431, 
    0.01466631, 0.01865058, 0.1577531, 0.1150998, 0.03756054, 0.01453416, 
    0.07593863, 0.0339271, 0.05533104, 0.1000932, 0.05830571, 0.03185456, 
    0.0115119, 0.003068706, 0.004355724, 0.01861754, 0.1774524, 0.2020815, 
    0.1788334, 0.108525, 0.01730832, 0.007627664, 0.02517182,
  0.4714819, 0.2063862, 0.1036665, 0.07483757, 0.05229317, 0.0548322, 
    0.0412382, 0.04178703, 0.03741582, 0.03388334, 0.01716864, 0.03787274, 
    0.03664718, 0.02546196, 0.03047504, 0.02263238, 0.02266264, 0.01364285, 
    0.01513806, 0.01123193, 0.02045063, 0.06959517, 0.2387962, 0.01266025, 
    0.04085729, 0.01967436, 0.0254829, 0.03590105, 0.1482747,
  0.03643867, 0.001026716, 0.0005277722, 0.00680114, 0.05907815, 0.1122352, 
    0.06988411, 0.08863281, 0.1268086, 0.09067017, 0.1086318, 0.1838418, 
    0.03151608, 0.02349411, 0.03231192, 0.0429244, 0.02806123, 0.02341074, 
    0.03087967, 0.06606349, 0.1441115, 0.1584483, 0.09039444, 0.003875381, 
    0.03906036, 0.06719634, 0.02563299, 0.06895523, 0.05890113,
  5.471426e-09, 4.542217e-09, 1.115274e-09, -0.00298285, 0.09663334, 
    0.04080191, -0.002573817, 0.07037732, 0.02222245, 0.04725251, 0.1542346, 
    0.0792513, 0.04004497, 0.02289485, 0.02673807, 0.03831148, 0.05762068, 
    0.03339902, 0.05687628, 0.05527548, 0.06352875, 0.0321939, 0.3505829, 
    0.1206741, 0.007590373, 0.03039568, 0.05355852, -5.262938e-05, 
    -1.286009e-06,
  3.456347e-08, 2.314541e-09, 7.054954e-10, 0.003337769, 2.212765e-08, 
    0.004972306, 0.00172492, 0.02412038, 0.01620284, 0.1997541, 0.04565313, 
    0.05533008, 0.08365232, 0.09035827, 0.0762258, 0.0325217, 0.05669857, 
    0.05091344, 0.0831112, 0.1115213, 0.04273847, 0.2123991, 0.02653116, 
    0.04939089, 0.05673822, 0.03127711, 0.02821486, 0.0006284356, 3.384065e-08,
  0.0002161835, 0.02949617, 0.009030622, 0.03158682, 0.09183934, 0.004783132, 
    0.007700851, 0.009656745, 0.02283442, 0.051648, 0.05231591, 0.01847533, 
    0.03284028, 0.08008357, 0.06653672, 0.09166677, 0.05901386, 0.1204176, 
    0.1480709, 0.1204877, 0.02156809, 0.1152148, 0.09855603, 0.03181517, 
    0.04961557, 0.09468643, 0.08279003, 0.1601408, 0.02763685,
  0.01729936, 0.05318953, 0.1497395, 0.3716173, 0.0515751, 0.06128447, 
    0.1624098, 0.01419562, 0.0005149317, 0.01375704, 0.08430605, 0.07549363, 
    0.1099486, 0.1226721, 0.1409802, 0.1636835, 0.1489455, 0.2038287, 
    0.2372644, 0.3778902, 0.161903, 0.09011425, 0.3425949, 0.2327019, 
    0.1876617, 0.1945829, 0.1845017, 0.1720436, 0.2896393,
  0.3067803, 0.3650764, 0.2839574, 0.3478104, 0.3469, 0.4043746, 0.1116647, 
    0.1219035, 0.05650702, 0.05675282, 0.1151772, 0.305732, 0.3438632, 
    0.2904779, 0.3211196, 0.2579648, 0.2779231, 0.19639, 0.2075063, 
    0.3325213, 0.1569146, 0.3418391, 0.3054048, 0.3683325, 0.387145, 
    0.2238823, 0.2713717, 0.1964232, 0.1926546,
  0.1679294, 0.1853291, 0.2482727, 0.5408015, 0.640243, 0.397236, 0.6145945, 
    0.523301, 0.4432611, 0.5041767, 0.5124056, 0.2128868, 0.2124791, 
    0.2265977, 0.41387, 0.3144041, 0.3509143, 0.3909312, 0.4656986, 
    0.2339291, 0.3548904, 0.2677846, 0.1904455, 0.1094741, 0.6054901, 
    0.1135523, 0.2254236, 0.1999744, 0.1808065,
  0.1013496, 0.06989624, 0.2118005, 0.2032022, 0.5037847, 0.5106124, 
    0.6224787, 0.6129884, 0.3342286, 0.4899983, 0.4942856, 0.3697604, 
    0.4366136, 0.4059531, 0.5133402, 0.2556018, 0.5196752, 0.632899, 
    0.3283457, 0.4806539, 0.3812051, 0.2195427, 0.3151262, 0.1340993, 
    0.1549967, 0.5643258, 0.1541241, 0.1098185, 0.2298739,
  0.2545707, 0.3444769, 0.4040787, 0.3151406, 0.3317782, 0.4485909, 
    0.4726231, 0.4539118, 0.4184242, 0.4321176, 0.4242695, 0.4521697, 
    0.5112625, 0.5698227, 0.5452654, 0.5492264, 0.4227606, 0.2899612, 
    0.3611756, 0.4604598, 0.4523572, 0.3178052, 0.1912451, 0.1622324, 
    0.1835458, 0.2396416, 0.1386124, 0.2632405, 0.4633456,
  0.2703033, 0.2749571, 0.279611, 0.2842648, 0.2889187, 0.2935725, 0.2982264, 
    0.3185563, 0.3111595, 0.3037626, 0.2963657, 0.2889689, 0.281572, 
    0.2741752, 0.3070595, 0.3072574, 0.3074555, 0.3076534, 0.3078514, 
    0.3080494, 0.3082474, 0.3127391, 0.3152841, 0.3178291, 0.3203741, 
    0.3229191, 0.3254642, 0.3280092, 0.2665802,
  0.229144, 0.2730744, 0.3108729, 0.3154697, 0.1372461, 0.1239211, 0.1494556, 
    0.1599912, 0.1354214, 0.2815374, 0.3270128, 0.2187504, 0.2961664, 
    0.04739109, 0.2138294, 0.2282733, 0.1282836, 0.1645068, 0.1836793, 
    0.1187209, 0.2139455, 0.3005202, 0.1522904, 0.04963164, 0.1485722, 
    0.1852511, 0.1833978, 0.0773446, 0.1533161,
  0.2336854, 0.211866, 0.2824288, 0.1216605, 0.06941417, 0.3191116, 
    0.02482055, 0.06298694, 0.07174672, 0.1133969, 0.1917779, 0.2057207, 
    0.06505381, 0.3099023, 0.4468115, 0.4091842, 0.4163618, 0.4154219, 
    0.4298839, 0.5274133, 0.4296102, 0.4702141, 0.5788945, 0.3274591, 
    0.3402011, 0.3259471, 0.3558352, 0.2753344, 0.2450367,
  0.4734031, 0.4994401, 0.4007769, 0.3897384, 0.4819414, 0.5822116, 
    0.4616177, 0.343408, 0.5043896, 0.4291252, 0.4579582, 0.4587049, 
    0.4299093, 0.3532313, 0.3372943, 0.4235853, 0.558199, 0.4922811, 
    0.4933888, 0.4496998, 0.3280429, 0.3753822, 0.2870956, 0.3463975, 
    0.3757999, 0.4487882, 0.4189634, 0.3922915, 0.4697577,
  0.4105104, 0.3720998, 0.4120248, 0.3390059, 0.4391142, 0.3314841, 
    0.3317378, 0.263721, 0.2982803, 0.3482225, 0.3051088, 0.2448984, 
    0.1991981, 0.2329154, 0.1064139, 0.1946121, 0.2856227, 0.3406963, 
    0.4073211, 0.4331455, 0.4283605, 0.314842, 0.2762689, 0.1490069, 
    0.04128028, 0.1674245, 0.3486317, 0.3887881, 0.3880184,
  0.1396899, 0.1022959, 0.1058377, 0.1486781, 0.2819594, 0.2193502, 
    0.1867768, 0.1396511, 0.1897044, 0.120818, 0.1467431, 0.04822324, 
    0.06987421, 0.1166351, 0.1859508, 0.1298293, 0.2005779, 0.2013165, 
    0.2562322, 0.2586725, 0.235595, 0.1405445, 0.09633899, 0.1888256, 
    0.01159712, 0.1665724, 0.2854895, 0.3325987, 0.2229558,
  0.03520789, 0.02370118, 0.0512959, 0.09481534, 0.08690671, 0.0593513, 
    0.02495456, 0.02868463, 0.04485812, 0.03225543, 3.346627e-05, 
    -3.142054e-10, 0.02844979, 0.07111169, 0.0799267, 0.0251886, 0.1970708, 
    0.3629017, 0.09752852, 0.04888855, 0.02149145, 0.007548975, 0.02572864, 
    0.05970703, 0.06861006, 0.06745325, 0.06688095, 0.01936033, 0.02444481,
  0.04380786, 0.08087825, 0.03300524, 0.02009732, 0.000633658, 0.002501398, 
    0.003429299, 0.003726533, 0.04621173, 0.08449119, 0.03060771, 
    0.009389579, 0.03903378, 0.01065582, 0.01941614, 0.0565339, 0.02551579, 
    0.01192341, 0.0008360025, 8.074158e-05, 5.503179e-05, 0.002258245, 
    0.04929929, 0.1921865, 0.1470129, 0.1028307, 0.004517326, 0.0003302449, 
    0.00393753,
  0.136985, 0.1070554, 0.09520793, 0.06765584, 0.01755302, 0.01382122, 
    0.0167245, 0.0195197, 0.0110136, 0.005926427, 0.008459367, 0.003662039, 
    0.01272442, 0.005351186, 0.005102965, 0.007850461, 0.01214893, 
    0.004728004, 0.002593141, 0.002152669, 0.004579757, 0.01941137, 
    0.04711889, 0.00551731, 0.03339955, 0.01208113, 0.004703417, 0.008204662, 
    0.03805853,
  0.004144323, 0.0003940702, 0.0002829301, 0.005127691, 0.02126266, 
    0.01508152, 0.03456506, 0.01717507, 0.07910489, 0.05687614, 0.02477962, 
    0.02142423, 0.01260694, 0.003315854, 0.008333306, 0.01313557, 0.01057109, 
    0.007888949, 0.01147834, 0.02337175, 0.07012707, 0.1956011, 0.2738048, 
    0.00113741, 0.02247315, 0.05038624, 0.004676843, 0.007649272, 0.01113821,
  5.230068e-09, 4.160622e-09, 8.50029e-10, -0.003289833, 0.04361998, 
    0.01031775, -0.002658783, 0.01342443, 0.003554858, 0.01427826, 
    0.08087259, 0.04513792, 0.02416806, 0.01036358, 0.004308217, 0.01079999, 
    0.01701213, 0.01477158, 0.02310469, 0.03054461, 0.02716469, 0.01351658, 
    0.3844523, 0.1267815, 0.0009976866, 0.006495613, 0.01596811, 
    -6.637179e-06, -4.824167e-07,
  5.542955e-09, 1.568449e-09, 2.089601e-10, -0.000329938, 9.630432e-09, 
    0.002144116, 0.001189108, 0.01183062, 0.02063544, 0.1490623, 0.01704398, 
    0.02699942, 0.03868291, 0.0297653, 0.01752857, 0.006648968, 0.01203986, 
    0.01048338, 0.05390496, 0.0497588, 0.04268579, 0.147134, 0.01147403, 
    0.01680081, 0.01194159, 0.005782969, 0.00696829, 0.0002406651, 
    6.680235e-09,
  -0.0001559285, 0.02227332, 0.005749016, 0.02437697, 0.0875859, 0.000388967, 
    0.004245539, 0.008982624, 0.01942508, 0.0475736, 0.03204492, 0.01317527, 
    0.02302668, 0.06342797, 0.05214078, 0.06751952, 0.03803948, 0.1061386, 
    0.1118464, 0.138699, 0.02381778, 0.1114408, 0.06994728, 0.02273129, 
    0.0387395, 0.08067971, 0.0434255, 0.08263863, 0.02790155,
  0.006568849, 0.03456019, 0.09517477, 0.3384269, 0.02198869, 0.08372337, 
    0.1419884, 0.01351534, 0.0001146026, 0.01001174, 0.06234247, 0.04482745, 
    0.07547202, 0.1009588, 0.1055149, 0.1386621, 0.1173511, 0.1803255, 
    0.2295996, 0.3658152, 0.1384884, 0.07277464, 0.3064766, 0.1812508, 
    0.143064, 0.1471247, 0.1749047, 0.1769408, 0.2513472,
  0.2463057, 0.3439196, 0.3000794, 0.3477772, 0.3319065, 0.388924, 0.0682809, 
    0.1134256, 0.05749705, 0.06839833, 0.1076996, 0.3461656, 0.2611369, 
    0.2388071, 0.2624733, 0.1764118, 0.2332928, 0.160721, 0.2149573, 
    0.3515467, 0.1629816, 0.3563052, 0.3490078, 0.4237696, 0.366896, 
    0.1843522, 0.2229459, 0.155786, 0.1543345,
  0.1310015, 0.2071688, 0.2645233, 0.6298556, 0.6936072, 0.4416884, 0.638874, 
    0.5654522, 0.4731975, 0.5537083, 0.5505485, 0.2715102, 0.2094727, 
    0.2106149, 0.3336068, 0.2180376, 0.3922642, 0.3444217, 0.4759686, 
    0.2832009, 0.4660413, 0.2802431, 0.2640544, 0.1512648, 0.5075324, 
    0.08886223, 0.1935003, 0.1585524, 0.1346596,
  0.05909876, 0.05227132, 0.1713356, 0.1640253, 0.5186672, 0.5668151, 
    0.6560461, 0.5931057, 0.312592, 0.4547115, 0.5546018, 0.3765176, 
    0.436761, 0.4142902, 0.5273237, 0.2869083, 0.5615875, 0.6289989, 0.36293, 
    0.5364577, 0.4099294, 0.2497868, 0.3816839, 0.1380804, 0.1444676, 
    0.5432483, 0.1712068, 0.105137, 0.1801732,
  0.3519327, 0.3937253, 0.4967637, 0.3562616, 0.3914448, 0.5315636, 
    0.5380915, 0.4912551, 0.4681976, 0.5379437, 0.5102604, 0.4916638, 
    0.5350986, 0.5849479, 0.5711217, 0.5503855, 0.4349643, 0.3131498, 
    0.402801, 0.5277842, 0.5177391, 0.3145117, 0.2075762, 0.2111027, 
    0.2080038, 0.2437078, 0.129497, 0.2483048, 0.5339603,
  0.2689278, 0.2741974, 0.279467, 0.2847366, 0.2900062, 0.2952757, 0.3005453, 
    0.3102272, 0.3052164, 0.3002056, 0.2951948, 0.290184, 0.2851732, 
    0.2801624, 0.3034653, 0.30046, 0.2974547, 0.2944494, 0.2914441, 
    0.2884387, 0.2854334, 0.339519, 0.3422655, 0.345012, 0.3477586, 
    0.3505051, 0.3532516, 0.3559981, 0.2647122,
  0.1832122, 0.2486309, 0.2516188, 0.2507927, 0.1411708, 0.09651097, 
    0.111502, 0.1273663, 0.1072624, 0.2212859, 0.2119697, 0.1327743, 
    0.2203036, 0.03639461, 0.1694294, 0.167854, 0.07749775, 0.1144412, 
    0.1217199, 0.08434123, 0.1536938, 0.213037, 0.1003782, 0.0530333, 
    0.1414998, 0.156589, 0.108032, 0.05393597, 0.1160135,
  0.162192, 0.1667591, 0.1811729, 0.09456396, 0.03396088, 0.2560957, 
    0.03100165, 0.03205426, 0.04484883, 0.06991011, 0.1341797, 0.1584291, 
    0.05876352, 0.2424921, 0.3271889, 0.3240542, 0.3518291, 0.3522427, 
    0.369952, 0.4628789, 0.4350152, 0.4086343, 0.5228142, 0.3080776, 
    0.3506608, 0.2870371, 0.3105047, 0.2117802, 0.1733336,
  0.437313, 0.4558392, 0.3350127, 0.3193647, 0.3996775, 0.513648, 0.4435991, 
    0.2705971, 0.4383462, 0.3896061, 0.4547388, 0.4379019, 0.4297126, 
    0.315293, 0.296122, 0.3577064, 0.4918809, 0.4850647, 0.4373839, 
    0.3718562, 0.2677381, 0.3196891, 0.2334698, 0.2930934, 0.3061048, 
    0.3930309, 0.3532451, 0.3077681, 0.4282275,
  0.3800457, 0.3453952, 0.3791461, 0.3473623, 0.4118185, 0.3113205, 
    0.3007256, 0.2136918, 0.2366092, 0.2995811, 0.2518193, 0.2170166, 
    0.1653623, 0.2131754, 0.07311895, 0.2003098, 0.2621857, 0.2782056, 
    0.363102, 0.4240197, 0.371293, 0.2698639, 0.2509797, 0.11914, 0.04878436, 
    0.195571, 0.4017416, 0.3976333, 0.3841486,
  0.1085596, 0.06283565, 0.0706342, 0.128453, 0.2921013, 0.1733919, 
    0.1359178, 0.08922492, 0.1591014, 0.07277793, 0.06789482, 0.02361186, 
    0.05387837, 0.1079002, 0.1654026, 0.07269181, 0.1803673, 0.164495, 
    0.1509181, 0.2461129, 0.1723442, 0.07053913, 0.04981101, 0.1862897, 
    0.03494879, 0.1312624, 0.2902566, 0.3125913, 0.1881762,
  0.00735328, 0.006447796, 0.0365287, 0.05944719, 0.07289607, 0.01568969, 
    0.009451655, 0.009963682, 0.01950246, 0.009617614, -4.724384e-05, 
    2.372237e-08, 0.02394261, 0.02701987, 0.04578146, 0.01244855, 0.1394187, 
    0.25061, 0.05898992, 0.01310165, 0.0070247, 0.003407166, 0.01154922, 
    0.06789978, 0.05787888, 0.07888185, 0.04149936, 0.004237229, 0.006929375,
  0.01301052, 0.09567783, 0.02148147, 0.003997888, -0.004319078, 
    0.0002894392, 0.00100381, 0.001573278, 0.0164536, 0.03064157, 0.02485043, 
    0.005566856, 0.01277056, 0.002651017, 0.003155425, 0.03368341, 
    0.004957023, 0.002362774, 3.459708e-05, 1.510796e-05, 9.572285e-06, 
    0.0006634707, 0.01708322, 0.07537889, 0.1195493, 0.1001548, 0.00147558, 
    8.520995e-05, 0.0006400055,
  0.05343185, 0.03233116, 0.09147637, 0.04436963, 0.005350724, 0.001689545, 
    0.004373736, 0.003131995, 0.002302665, 0.0009391147, 0.003237803, 
    0.0004583008, 0.001622556, 0.001448131, 0.0005084504, 0.002906738, 
    0.007866402, 0.002064266, 0.000607761, 0.001051354, 0.002157828, 
    0.008522779, 0.01905769, 0.003067289, 0.03700707, 0.01049864, 
    0.001176729, 0.003398389, 0.01357706,
  0.0007003684, 0.0002248066, 0.000158446, 0.005460195, 0.008938201, 
    0.002596124, 0.01129908, 0.002219256, 0.05456821, 0.03748981, 
    0.005444372, 0.006000965, 0.005798672, 0.000354723, 0.003197186, 
    0.002297957, 0.0009055699, 0.002063165, 0.003122927, 0.004882974, 
    0.01664136, 0.04190581, 0.06725631, 0.0003645723, 0.01462194, 0.04331521, 
    0.0006227779, 0.002149204, 0.002107233,
  5.08285e-09, 4.029074e-09, 7.7583e-10, -0.002501811, 0.01726874, 
    0.002761068, -0.001756769, 0.003865888, 0.001230379, 0.003166043, 
    0.03288983, 0.0152663, 0.01146669, 0.004126945, 0.0006776942, 
    0.002525534, 0.005743562, 0.005221463, 0.008178595, 0.0109723, 
    0.01722212, 0.009779434, 0.3027794, 0.1072537, 0.0003003429, 0.002690538, 
    0.006800178, -1.795611e-06, -4.285262e-07,
  -1.066647e-09, 1.504054e-09, 2.370767e-10, -0.0004039216, 7.000431e-09, 
    0.001251539, 0.00110015, 0.00403628, 0.02761229, 0.07774459, 0.006340726, 
    0.01521893, 0.01910108, 0.007328744, 0.005027631, 0.002730778, 
    0.004228372, 0.00407459, 0.02117218, 0.02268327, 0.0218776, 0.1208113, 
    0.005411223, 0.003522365, 0.003319819, 0.002057007, 0.00313576, 
    0.0001282509, 3.728474e-09,
  -0.000179897, 0.01369494, 0.001130831, 0.01670109, 0.08122931, 
    -0.001137679, 0.002958112, 0.009608601, 0.0164539, 0.05067149, 
    0.02301629, 0.008025425, 0.01521202, 0.04563642, 0.03186805, 0.04594684, 
    0.02273057, 0.06998666, 0.07524614, 0.07514388, 0.02931115, 0.108006, 
    0.05655431, 0.01666437, 0.02725029, 0.06589172, 0.02264605, 0.02933786, 
    0.02012523,
  0.002385471, 0.02341854, 0.06476495, 0.3099637, 0.009781418, 0.08494645, 
    0.1280224, 0.01071645, -5.890915e-05, 0.006634629, 0.04385829, 
    0.02863649, 0.05721725, 0.0879679, 0.07800627, 0.1168195, 0.102922, 
    0.1452716, 0.1772509, 0.3454194, 0.1205297, 0.0585011, 0.2472055, 
    0.1528271, 0.09479187, 0.1263257, 0.1390233, 0.1165393, 0.2077635,
  0.1802553, 0.3014211, 0.2785322, 0.3393691, 0.286316, 0.3381565, 
    0.03892827, 0.1029036, 0.05392679, 0.07132579, 0.09293502, 0.3791293, 
    0.2086445, 0.1850169, 0.2192786, 0.1460632, 0.2027106, 0.1323405, 
    0.1866661, 0.3786363, 0.1598841, 0.3157432, 0.3636766, 0.4161154, 
    0.278088, 0.1448086, 0.1857697, 0.11466, 0.1309984,
  0.1039079, 0.1973284, 0.3347509, 0.6778048, 0.7198774, 0.5016139, 
    0.5815119, 0.5395504, 0.5159763, 0.5769837, 0.5773445, 0.3588218, 
    0.202625, 0.2060406, 0.2727374, 0.226263, 0.4521058, 0.3164295, 
    0.4746844, 0.3210306, 0.5868077, 0.2332734, 0.3113029, 0.2072405, 
    0.4354019, 0.06914837, 0.1606381, 0.1181673, 0.1044699,
  0.04041301, 0.03978024, 0.1406767, 0.1190144, 0.4389452, 0.6279389, 
    0.8006266, 0.5348891, 0.3015583, 0.4099596, 0.56573, 0.4417549, 
    0.4878452, 0.4120587, 0.5234673, 0.3210206, 0.6387644, 0.6458958, 
    0.4466632, 0.5773792, 0.3594835, 0.3048458, 0.4571706, 0.1553575, 
    0.1397871, 0.4870054, 0.1939166, 0.1, 0.142781,
  0.5027321, 0.4970677, 0.5552808, 0.4826445, 0.4836788, 0.6177313, 
    0.5787752, 0.5671626, 0.6104237, 0.6170743, 0.549014, 0.5408875, 
    0.6310064, 0.61027, 0.5751505, 0.5419362, 0.4612156, 0.3639987, 
    0.4785304, 0.592352, 0.5779119, 0.2879075, 0.2757252, 0.2614703, 
    0.1773051, 0.2229736, 0.1207351, 0.2459332, 0.6102465,
  0.2748757, 0.2809682, 0.2870606, 0.293153, 0.2992454, 0.3053379, 0.3114303, 
    0.2842204, 0.2814619, 0.2787034, 0.2759449, 0.2731864, 0.2704278, 
    0.2676693, 0.3063928, 0.2999921, 0.2935914, 0.2871906, 0.2807899, 
    0.2743891, 0.2679884, 0.3172679, 0.3203347, 0.3234015, 0.3264684, 
    0.3295352, 0.3326021, 0.3356689, 0.2700018,
  0.1385254, 0.198225, 0.1832338, 0.1873788, 0.11788, 0.07099578, 0.08427884, 
    0.09808168, 0.07923149, 0.1508718, 0.1315664, 0.08176906, 0.1350155, 
    0.03505892, 0.1447435, 0.1220741, 0.05593548, 0.07643699, 0.08418173, 
    0.05472568, 0.1167708, 0.1527823, 0.05785425, 0.04395968, 0.1671344, 
    0.134144, 0.094005, 0.0341715, 0.07099399,
  0.1099081, 0.1213306, 0.1263517, 0.07109819, 0.01502489, 0.2129574, 
    0.04181542, 0.01699309, 0.02730461, 0.04650136, 0.09340197, 0.1212582, 
    0.04470645, 0.1844974, 0.2447763, 0.2532496, 0.2845194, 0.2662364, 
    0.3028363, 0.3780916, 0.3822989, 0.4027493, 0.4902173, 0.2799897, 
    0.3036725, 0.2794012, 0.2736608, 0.1532028, 0.10815,
  0.3800749, 0.3687563, 0.2516226, 0.2402417, 0.3092896, 0.4281842, 
    0.3705407, 0.2050139, 0.3373695, 0.3424377, 0.4293195, 0.4054043, 
    0.4058428, 0.2663332, 0.2467552, 0.3027785, 0.4264084, 0.4586388, 
    0.4035028, 0.3063515, 0.2150909, 0.2458315, 0.1791236, 0.2429151, 
    0.280236, 0.3333322, 0.2968527, 0.2336915, 0.3611696,
  0.3220631, 0.2680014, 0.3073061, 0.3288087, 0.3645693, 0.2800028, 
    0.2537545, 0.1617707, 0.1851614, 0.2358922, 0.1935637, 0.1651351, 
    0.1305801, 0.1685937, 0.05255734, 0.1522402, 0.2103476, 0.2295253, 
    0.285648, 0.3576304, 0.3012002, 0.2031144, 0.2001138, 0.09124607, 
    0.03888317, 0.2369705, 0.3795387, 0.3608975, 0.3426853,
  0.07401668, 0.03739735, 0.04970834, 0.1063411, 0.2515562, 0.1283749, 
    0.09716932, 0.05970429, 0.1207041, 0.04535978, 0.04135869, 0.01506073, 
    0.03772105, 0.08021768, 0.1474578, 0.04911172, 0.1439382, 0.12036, 
    0.1050439, 0.2123571, 0.1265174, 0.04399217, 0.02552419, 0.1752796, 
    0.03018807, 0.09349009, 0.2801627, 0.2642561, 0.148117,
  0.003340182, 0.003357865, 0.02244925, 0.02649974, 0.04037492, 0.002336997, 
    0.003512136, 0.005349116, 0.01145363, 0.004555539, -2.28196e-05, 
    4.910679e-08, 0.01978302, 0.00937293, 0.0275795, 0.005050666, 0.09832091, 
    0.1426754, 0.0522392, 0.004214021, 0.003898924, 0.001970431, 0.006901759, 
    0.04455282, 0.04359846, 0.05807791, 0.0216538, 0.002145284, 0.003540838,
  0.005636486, 0.07800407, 0.01293061, 0.001459474, -0.003816657, 
    6.97139e-05, 0.0004219489, 0.0009130831, 0.008509316, 0.0103731, 
    0.0157785, 0.003477823, 0.004487413, 0.0009449201, 0.001054479, 
    0.01711015, 0.0009974859, 0.0004629718, 1.053153e-05, 3.88493e-06, 
    2.500119e-06, 0.0003188647, 0.008059315, 0.04042022, 0.09686363, 
    0.08344308, 0.0005127484, 3.586978e-05, 0.0002647571,
  0.02860148, 0.01488213, 0.08850822, 0.02327652, 0.002049054, 0.0003801134, 
    0.00144884, 0.0006921973, 0.001050372, 0.000282062, 0.001295475, 
    0.0001672888, -8.379747e-05, 0.0005204533, 0.0001818363, 0.001072088, 
    0.004688137, 0.0009845522, 0.0003272958, 0.0006287181, 0.001278816, 
    0.004907736, 0.01064846, 0.002900469, 0.05233315, 0.006745348, 
    0.000493886, 0.001974576, 0.00711665,
  0.0002846616, 0.0001781361, 7.557352e-05, 0.01002356, 0.001553391, 
    0.00124373, 0.004317003, 0.0007027817, 0.04845758, 0.0394198, 
    0.002422927, 0.002953632, 0.002963799, 0.000108169, 0.001536249, 
    0.000767481, 0.0002826238, 0.0009853889, 0.0009149562, 0.00153398, 
    0.004153755, 0.01384115, 0.02771601, 0.0002018045, 0.01034849, 
    0.02678697, 0.000211135, 0.001023239, 0.00104545,
  5.065919e-09, 3.982892e-09, 7.62282e-10, 0.0002271204, 0.008823743, 
    0.001254239, -0.001320376, 0.001945087, 0.0008256526, 0.0006330055, 
    0.0116816, 0.004485949, 0.004476083, 0.001876619, 0.000368574, 
    0.0009043511, 0.002561115, 0.002252101, 0.003494575, 0.004974838, 
    0.01056711, 0.007119074, 0.216837, 0.08679994, 0.0001385791, 0.001501397, 
    0.003826022, -7.460375e-07, -1.232012e-05,
  -3.483442e-09, 1.501403e-09, 5.947403e-10, -0.0002228919, 6.522319e-09, 
    0.0008540183, 0.000479575, 0.001884901, 0.04623203, 0.04152117, 
    0.002986081, 0.008547066, 0.009327595, 0.003314941, 0.002494811, 
    0.001735663, 0.002033088, 0.001244568, 0.01022131, 0.01332409, 
    0.01300175, 0.09368774, 0.003109641, -0.0002989036, 0.001715256, 
    0.001181151, 0.001849188, 8.195142e-05, 3.209763e-09,
  -0.0001203373, 0.008221732, 0.0006441388, 0.01037809, 0.07146072, 
    -0.001322442, 0.001769073, 0.01288437, 0.01291995, 0.03906394, 
    0.01799522, 0.004855774, 0.008525149, 0.03170785, 0.02006586, 0.02710399, 
    0.01140328, 0.04137775, 0.04347518, 0.04470508, 0.02715706, 0.1080009, 
    0.05291446, 0.01107155, 0.01671669, 0.04150242, 0.009502027, 0.01531549, 
    0.01355606,
  0.0004927504, 0.01156943, 0.04684824, 0.2818773, 0.005039095, 0.0656336, 
    0.1139834, 0.008412693, -8.442642e-05, 0.004967248, 0.02950137, 
    0.02107595, 0.04565554, 0.07615451, 0.05336815, 0.08999436, 0.08562409, 
    0.1034823, 0.116613, 0.321964, 0.1072535, 0.04850387, 0.1959974, 
    0.1294333, 0.06022992, 0.09836175, 0.09647228, 0.0668587, 0.1587323,
  0.1267421, 0.2583197, 0.2089096, 0.3345522, 0.2489069, 0.2855029, 
    0.02409755, 0.09226938, 0.04385176, 0.07179382, 0.06650875, 0.4178136, 
    0.1710852, 0.1452446, 0.1862457, 0.1262194, 0.1792147, 0.09637622, 
    0.1363514, 0.4099755, 0.1628561, 0.2364664, 0.3212105, 0.4186459, 
    0.2089451, 0.1123948, 0.147445, 0.08882017, 0.1066689,
  0.07167259, 0.2222928, 0.3110894, 0.6538901, 0.7241043, 0.4925706, 
    0.5041357, 0.4485811, 0.516211, 0.5385397, 0.5869897, 0.4366581, 
    0.1921777, 0.2451671, 0.2185672, 0.2506826, 0.4906528, 0.2745728, 
    0.4195103, 0.3765384, 0.6357248, 0.2193844, 0.2830917, 0.2067234, 
    0.3839111, 0.05136073, 0.1340209, 0.08554281, 0.07189675,
  0.03049611, 0.03023781, 0.156156, 0.08647119, 0.4050899, 0.6605142, 
    0.8210875, 0.4909984, 0.2816097, 0.4644193, 0.5716761, 0.4661126, 
    0.6829699, 0.4181119, 0.5040287, 0.3563053, 0.5793397, 0.5951602, 
    0.4180583, 0.531175, 0.3556165, 0.3686534, 0.5018503, 0.1982058, 
    0.2144553, 0.4331278, 0.2128271, 0.1049979, 0.1102943,
  0.584953, 0.5689881, 0.5932758, 0.5594079, 0.5500134, 0.6396872, 0.5456101, 
    0.5888736, 0.6553225, 0.6687621, 0.5428129, 0.5836306, 0.666252, 
    0.5780604, 0.5090459, 0.5163209, 0.5349583, 0.429725, 0.5551785, 
    0.5872219, 0.5466553, 0.280636, 0.3120445, 0.3179775, 0.139068, 
    0.2127081, 0.1130293, 0.2101626, 0.6392059,
  0.216422, 0.2239572, 0.2314923, 0.2390275, 0.2465626, 0.2540978, 0.2616329, 
    0.2157476, 0.2148561, 0.2139647, 0.2130733, 0.2121819, 0.2112905, 
    0.210399, 0.2837183, 0.2770138, 0.2703094, 0.263605, 0.2569006, 
    0.2501962, 0.2434917, 0.264695, 0.2647557, 0.2648164, 0.2648771, 
    0.2649378, 0.2649985, 0.2650591, 0.2103939,
  0.1053532, 0.1415415, 0.135984, 0.1556303, 0.1094943, 0.05325291, 
    0.06176831, 0.07138228, 0.06214998, 0.09945782, 0.0899852, 0.04778848, 
    0.07888185, 0.03404015, 0.112083, 0.0781533, 0.03628513, 0.0470045, 
    0.0630115, 0.03429186, 0.09304159, 0.1210008, 0.03934442, 0.03756535, 
    0.1414358, 0.114764, 0.08533641, 0.02427911, 0.04689875,
  0.07284372, 0.08466832, 0.09576013, 0.05441547, 0.007136996, 0.1735501, 
    0.03029625, 0.009781817, 0.01617762, 0.0352202, 0.06199824, 0.09652767, 
    0.03369631, 0.1350188, 0.1806618, 0.1984024, 0.2222505, 0.1989721, 
    0.2291184, 0.2826992, 0.3319843, 0.3642726, 0.4509876, 0.2278492, 
    0.2543813, 0.2496275, 0.229866, 0.1055497, 0.07046727,
  0.2975492, 0.2724094, 0.1697643, 0.1742689, 0.2200754, 0.3251838, 
    0.2875072, 0.1492301, 0.2564217, 0.2918428, 0.3584725, 0.332225, 
    0.3574607, 0.199233, 0.1787952, 0.2398255, 0.3403529, 0.405803, 
    0.3367969, 0.2333881, 0.1633744, 0.1736832, 0.1277763, 0.1764276, 
    0.241038, 0.276329, 0.2276117, 0.1740728, 0.2725138,
  0.2520767, 0.1985581, 0.2325063, 0.2712688, 0.2963803, 0.2327579, 
    0.2059242, 0.1219234, 0.1346812, 0.1665602, 0.1237232, 0.103445, 
    0.08899709, 0.11456, 0.03309148, 0.1113689, 0.1469423, 0.1786417, 
    0.217738, 0.2629319, 0.2077254, 0.1398997, 0.1304471, 0.07111551, 
    0.02758587, 0.2079625, 0.3265675, 0.3029595, 0.2857529,
  0.04812164, 0.02178377, 0.03394932, 0.07716336, 0.1839294, 0.07999422, 
    0.06444254, 0.03243572, 0.0820049, 0.02877604, 0.02797041, 0.009619007, 
    0.02821566, 0.05076392, 0.128635, 0.03105243, 0.09690346, 0.0830472, 
    0.0694133, 0.1629819, 0.0888728, 0.025635, 0.01414338, 0.1572816, 
    0.02241517, 0.06513516, 0.2302572, 0.1897075, 0.1042368,
  0.002090455, 0.002205104, 0.01382934, 0.01090976, 0.01933784, 0.00103961, 
    0.00226133, 0.003775283, 0.007840021, 0.002212929, -1.560881e-05, 
    4.265839e-08, 0.01479812, 0.004184233, 0.01611809, 0.003014037, 
    0.06302001, 0.08806217, 0.02257707, 0.002069867, 0.002621958, 
    0.001327937, 0.004765389, 0.02893785, 0.02920471, 0.02761301, 
    0.006254899, 0.001390818, 0.002346217,
  0.003208189, 0.04899814, 0.00732309, 0.0007921431, -0.002856236, 
    3.890798e-05, 0.0002010339, 0.0006158353, 0.005402497, 0.005338081, 
    0.01073475, 0.000947126, 0.001971334, 0.0005791153, 0.0006472598, 
    0.006790624, 0.0005158094, 0.0001891305, 5.808005e-06, 2.475285e-06, 
    1.410859e-06, 0.0001906623, 0.004802762, 0.02645482, 0.07224624, 
    0.06621864, 0.0002467727, 1.943806e-05, 0.0001492917,
  0.01886582, 0.009148893, 0.08093786, 0.01245635, 0.000691565, 0.0002067175, 
    0.0007298119, 0.0002214272, 0.0006843169, 0.0001837284, 0.0004982182, 
    8.949461e-05, -7.708877e-05, 0.0002881328, 0.000102271, 0.0005238691, 
    0.002193118, 0.0005474054, 0.0002099832, 0.0004286386, 0.0008732981, 
    0.003287372, 0.007100545, 0.002864277, 0.0444099, 0.004047381, 
    0.0002453636, 0.001332975, 0.004599586,
  0.0001495239, 0.0006056053, 5.196197e-05, 0.009701422, 0.00059461, 
    0.0007769832, 0.00171329, 0.0004207421, 0.05371304, 0.03743201, 
    0.001477296, 0.001814559, 0.001330789, 6.287575e-05, 0.0007859955, 
    0.0004305311, 0.0001604977, 0.000636122, 0.0004951871, 0.0007827985, 
    0.002209943, 0.007346779, 0.01611362, 0.0001288718, 0.007442195, 
    0.01358849, 0.0001136872, 0.0006148616, 0.000669062,
  5.244676e-09, 3.989099e-09, 7.661018e-10, 0.001411016, 0.004605449, 
    0.0007813726, -0.0008268402, 0.001176389, 0.0006044915, 0.0001758895, 
    0.004022918, 0.001653692, 0.001628534, 0.0007330917, 0.0002625902, 
    0.0005561205, 0.001275142, 0.0007390382, 0.001674292, 0.00192092, 
    0.00508684, 0.003733815, 0.1620786, 0.07061815, 0.0001073103, 
    0.0009836463, 0.002530011, -3.955706e-07, -6.20439e-05,
  -1.858039e-09, 1.586669e-09, 7.188553e-10, -0.000113976, 6.38563e-09, 
    0.0006429981, 0.0004612936, 0.001243367, 0.04837319, 0.02584759, 
    0.001953921, 0.00491379, 0.004441758, 0.002180443, 0.001612287, 
    0.001266257, 0.001184761, 0.0006620353, 0.006092595, 0.009280063, 
    0.009243381, 0.07796965, 0.00217797, -0.0009372335, 0.00125141, 
    0.0008119419, 0.001269641, 5.915025e-05, 3.096592e-09,
  -6.725131e-05, 0.005294065, 0.0004491387, 0.004648038, 0.06114404, 
    -0.001264133, 0.003310474, 0.02093105, 0.01152078, 0.02639006, 0.0149108, 
    0.00313012, 0.004600987, 0.01815244, 0.01084069, 0.01301775, 0.004552327, 
    0.0233452, 0.01847719, 0.02141351, 0.02459274, 0.1015102, 0.04452211, 
    0.004846005, 0.008199224, 0.02404945, 0.003862437, 0.009112734, 
    0.009028444,
  6.425769e-05, 0.004808846, 0.03487131, 0.2550685, 0.00324305, 0.05204629, 
    0.1017658, 0.007137323, -0.0001109067, 0.004759578, 0.01998237, 
    0.01653295, 0.0353035, 0.0587816, 0.0335258, 0.06100309, 0.05773562, 
    0.06937899, 0.07456877, 0.2965915, 0.1005594, 0.03701246, 0.1603289, 
    0.1104774, 0.03999015, 0.06997719, 0.06326662, 0.03900452, 0.1090777,
  0.08497514, 0.2242061, 0.1573985, 0.3047073, 0.2031668, 0.2442962, 
    0.01758326, 0.08431857, 0.05089073, 0.06898735, 0.04651501, 0.4434099, 
    0.1469791, 0.1168938, 0.1543378, 0.1070605, 0.1416743, 0.06488506, 
    0.08770397, 0.3899585, 0.1342623, 0.1700064, 0.2437186, 0.394809, 
    0.1596441, 0.08935648, 0.1120412, 0.0587332, 0.0720479,
  0.03840378, 0.2492571, 0.2811657, 0.6034767, 0.6570811, 0.4376121, 
    0.4286589, 0.3468212, 0.4449546, 0.4641535, 0.4996593, 0.5315673, 
    0.2222484, 0.2808916, 0.1806771, 0.281837, 0.5152075, 0.2522117, 
    0.3700707, 0.355717, 0.6477455, 0.2648769, 0.2533733, 0.2132331, 
    0.3427956, 0.0376638, 0.10315, 0.0634482, 0.04831509,
  0.02435619, 0.02366344, 0.1797583, 0.0673025, 0.3709871, 0.5680469, 
    0.7714664, 0.5029964, 0.3332936, 0.4641258, 0.5630941, 0.4130129, 
    0.640073, 0.3684864, 0.4257164, 0.3112039, 0.529681, 0.5026876, 
    0.2748694, 0.388074, 0.2601278, 0.3299702, 0.4869734, 0.2627419, 
    0.2400357, 0.3800944, 0.2390294, 0.0994409, 0.08633754,
  0.6264374, 0.610549, 0.5715014, 0.5614708, 0.5551355, 0.5528134, 0.4445317, 
    0.5036764, 0.5346583, 0.5800551, 0.5320628, 0.5731481, 0.6190768, 
    0.582037, 0.5157991, 0.5178187, 0.5731633, 0.465911, 0.5143177, 
    0.5823689, 0.5402002, 0.2897814, 0.3063519, 0.3616715, 0.1219706, 
    0.1819395, 0.1044029, 0.2133965, 0.5497022,
  0.1407903, 0.1463517, 0.151913, 0.1574743, 0.1630357, 0.168597, 0.1741583, 
    0.1445951, 0.1459574, 0.1473198, 0.1486821, 0.1500445, 0.1514068, 
    0.1527692, 0.2118687, 0.2065376, 0.2012064, 0.1958753, 0.1905442, 
    0.1852131, 0.1798819, 0.2069919, 0.2053993, 0.2038068, 0.2022142, 
    0.2006217, 0.1990291, 0.1974366, 0.1363412,
  0.07865272, 0.1105382, 0.1045134, 0.1262088, 0.1064394, 0.04073989, 
    0.04581126, 0.06391767, 0.05346925, 0.0658246, 0.06953915, 0.03163157, 
    0.0539804, 0.02808747, 0.0942017, 0.04675585, 0.0233924, 0.0355989, 
    0.05206114, 0.02649273, 0.0774676, 0.1045564, 0.02755022, 0.03674175, 
    0.1271894, 0.1039199, 0.08251993, 0.01945607, 0.03187037,
  0.05715016, 0.06716732, 0.07151274, 0.0466411, 0.005176484, 0.1466419, 
    0.02377528, 0.007019782, 0.01203398, 0.03135784, 0.04256625, 0.08231669, 
    0.0272643, 0.09636347, 0.1343473, 0.1493759, 0.1689127, 0.1576135, 
    0.1795707, 0.2162943, 0.2705854, 0.3049395, 0.3629769, 0.188593, 
    0.2083792, 0.2090385, 0.1843259, 0.08641554, 0.04973803,
  0.2397487, 0.2148418, 0.1276196, 0.1393522, 0.1685195, 0.2608728, 
    0.2279813, 0.1124633, 0.2023752, 0.2380788, 0.2757352, 0.2667622, 
    0.2955645, 0.1483391, 0.1285159, 0.1803183, 0.2659851, 0.3389058, 
    0.2625813, 0.1772126, 0.1221771, 0.1209995, 0.09374326, 0.1197037, 
    0.190227, 0.2153449, 0.1771656, 0.1352488, 0.2154276,
  0.2029994, 0.1586732, 0.1857843, 0.2226937, 0.2462236, 0.1993667, 
    0.1754571, 0.09806146, 0.102759, 0.1244403, 0.08416209, 0.06900446, 
    0.06348691, 0.07571873, 0.01743087, 0.08216747, 0.1032892, 0.1304992, 
    0.1703835, 0.1980473, 0.1477563, 0.1052464, 0.09023988, 0.06033513, 
    0.01868982, 0.1701746, 0.2776481, 0.2563654, 0.244454,
  0.03281672, 0.01443106, 0.02292663, 0.05163448, 0.1285115, 0.0488452, 
    0.04216872, 0.01975266, 0.05572557, 0.01779068, 0.01664234, 0.007071437, 
    0.02555166, 0.03282174, 0.1114672, 0.02017239, 0.05952428, 0.05497618, 
    0.04892768, 0.1101353, 0.0617132, 0.01412394, 0.009622982, 0.139256, 
    0.016467, 0.04396561, 0.1623778, 0.1328566, 0.07192884,
  0.001532094, 0.001636304, 0.008716484, 0.00573097, 0.01141097, 
    0.0007159443, 0.001731951, 0.002951687, 0.006027563, 0.001494795, 
    -1.237594e-05, 4.171257e-08, 0.01093442, 0.002687867, 0.009255481, 
    0.002273611, 0.04041085, 0.05316277, 0.01015964, 0.001379748, 
    0.001977749, 0.00100211, 0.003666973, 0.02243667, 0.0200959, 0.01316953, 
    0.002779031, 0.001034388, 0.001769451,
  0.002192004, 0.03390918, 0.004429169, 0.0005468766, -0.002011524, 
    2.676279e-05, 0.0001349007, 0.000465401, 0.003944434, 0.003477302, 
    0.006532379, 0.000507, 0.000966863, 0.0003637948, 0.0004664687, 
    0.003177283, 0.0003618037, 0.0001197208, 4.101812e-06, 1.77478e-06, 
    1.024585e-06, 0.0001331603, 0.003352117, 0.0198994, 0.04628347, 
    0.05793632, 0.0001614963, 1.29944e-05, 0.0001012563,
  0.0141001, 0.006492692, 0.07034595, 0.0206856, 0.0003620597, 0.0001547266, 
    0.0005377085, 0.000129871, 0.0005099721, 0.0001771443, 0.0002813724, 
    6.032067e-05, -1.825782e-05, 0.0001959309, 6.995395e-05, 0.0003518014, 
    0.001055171, 0.0003100054, 0.0001526431, 0.0003251438, 0.0006654828, 
    0.002474446, 0.00533532, 0.005082901, 0.02883554, 0.003692894, 
    0.0001518997, 0.001007817, 0.003390679,
  9.362464e-05, 0.001801858, 0.0004021826, 0.008480122, 0.0003769445, 
    0.0005686199, 0.000996858, 0.0003045466, 0.05379174, 0.05117903, 
    0.001049432, 0.001288439, 0.0007019969, 4.788038e-05, 0.0005231468, 
    0.0002979904, 0.0001080157, 0.0004666476, 0.0003216545, 0.0005070149, 
    0.001471795, 0.004841974, 0.01115717, 0.0004959033, 0.00550218, 
    0.006719631, 8.739608e-05, 0.0004300484, 0.0004948937,
  5.541201e-09, 4.047189e-09, 7.774139e-10, 0.002449773, 0.003026922, 
    0.0005754973, -0.0005119827, 0.0008656382, 0.000437586, 0.0001080896, 
    0.00181861, 0.0008258999, 0.0007676792, 0.0003561378, 0.0002057243, 
    0.0004042946, 0.0008534081, 0.0003382374, 0.000929716, 0.000819444, 
    0.002342436, 0.001826557, 0.117554, 0.05372053, 8.933162e-05, 
    0.0007290777, 0.001892856, -2.555821e-07, -0.0001003067,
  -1.143615e-09, 1.448979e-09, 6.848079e-10, -7.74698e-05, 6.307407e-09, 
    0.0005215167, 0.0006970941, 0.0009414882, 0.04639468, 0.01878782, 
    0.001492949, 0.002796272, 0.002326609, 0.001699628, 0.001194045, 
    0.0010115, 0.0008731453, 0.0004913309, 0.004325126, 0.007328053, 
    0.006496488, 0.0675813, 0.001700736, -0.001087893, 0.0009987586, 
    0.0006213111, 0.0009736631, 4.710249e-05, 3.101362e-09,
  -4.711686e-05, 0.003941481, 0.0003465121, 0.00340808, 0.05310098, 
    -0.001203048, 0.00591831, 0.03514592, 0.01033552, 0.01977173, 0.01297365, 
    0.002324557, 0.002890616, 0.007468317, 0.004970161, 0.005510791, 
    0.002271352, 0.012691, 0.01006256, 0.01340323, 0.02171932, 0.08547341, 
    0.04009479, 0.002761526, 0.004991323, 0.01339782, 0.002227685, 
    0.00646349, 0.006188548,
  4.772764e-05, 0.003013671, 0.02657765, 0.2365774, 0.0024724, 0.04225422, 
    0.0943192, 0.004711003, -0.0001669143, 0.005680291, 0.02161562, 
    0.01413878, 0.02747018, 0.04717207, 0.02423405, 0.04335249, 0.03648613, 
    0.04982021, 0.05061983, 0.2709793, 0.09817239, 0.03263418, 0.1419283, 
    0.1004232, 0.02996829, 0.04762965, 0.04278732, 0.02418477, 0.07615769,
  0.05994558, 0.2148826, 0.1503127, 0.2909926, 0.1765468, 0.2141428, 
    0.01920741, 0.09748384, 0.09743437, 0.06442073, 0.03752028, 0.4234498, 
    0.1305536, 0.09700385, 0.1173549, 0.08932207, 0.1093874, 0.04764448, 
    0.06274512, 0.382889, 0.1144169, 0.1414377, 0.197294, 0.3558857, 
    0.1307781, 0.07456197, 0.08702622, 0.03847232, 0.04555556,
  0.0240949, 0.2724096, 0.2760013, 0.5414695, 0.5769092, 0.3723188, 
    0.3558303, 0.2900616, 0.3671798, 0.3936033, 0.4316052, 0.5952458, 
    0.2786058, 0.3073308, 0.1573059, 0.3031118, 0.5113417, 0.2490412, 
    0.3750383, 0.346292, 0.596404, 0.2875983, 0.2042607, 0.1980849, 
    0.3137629, 0.02948079, 0.07885054, 0.04810816, 0.03476682,
  0.02081605, 0.01929678, 0.2628232, 0.05686204, 0.3523632, 0.431311, 
    0.7062991, 0.4582355, 0.4130372, 0.4245386, 0.587779, 0.3720724, 
    0.4810619, 0.2640752, 0.3087854, 0.2710785, 0.471377, 0.4035644, 
    0.2157311, 0.2506976, 0.1890214, 0.2581855, 0.39922, 0.2387626, 0.237734, 
    0.2937425, 0.3414131, 0.09748051, 0.07407655,
  0.6689566, 0.6199248, 0.5175571, 0.4308732, 0.446236, 0.4046735, 0.2417237, 
    0.2324101, 0.3462856, 0.3689813, 0.3265024, 0.3837272, 0.3976541, 
    0.3626725, 0.3685067, 0.3730989, 0.4762661, 0.4723472, 0.3300754, 
    0.3871473, 0.3499554, 0.2838666, 0.3117991, 0.4605854, 0.162753, 
    0.1519902, 0.09633106, 0.2089419, 0.4387113,
  0.09309179, 0.09744438, 0.101797, 0.1061495, 0.1105021, 0.1148547, 
    0.1192073, 0.09646735, 0.09859093, 0.1007145, 0.1028381, 0.1049617, 
    0.1070853, 0.1092089, 0.1569795, 0.1518123, 0.1466451, 0.1414779, 
    0.1363107, 0.1311435, 0.1259762, 0.1355557, 0.1342467, 0.1329377, 
    0.1316288, 0.1303198, 0.1290109, 0.1277019, 0.08960973,
  0.0689756, 0.1030117, 0.09412244, 0.1238292, 0.1556198, 0.03436021, 
    0.04023277, 0.09017467, 0.07772242, 0.066554, 0.05703929, 0.02587799, 
    0.04338637, 0.02405511, 0.09619343, 0.03553382, 0.01788937, 0.02979054, 
    0.04730627, 0.02659159, 0.06845894, 0.0917758, 0.02311781, 0.03750287, 
    0.1220693, 0.09651643, 0.07597479, 0.01802537, 0.03108344,
  0.05242927, 0.05701511, 0.05978625, 0.05012678, 0.003885041, 0.134996, 
    0.03119675, 0.006820034, 0.01521377, 0.03070742, 0.03598955, 0.07673238, 
    0.02430202, 0.081146, 0.1102222, 0.125322, 0.1384143, 0.1338057, 
    0.1545601, 0.1845286, 0.2310846, 0.2534638, 0.317275, 0.1664262, 
    0.1833717, 0.1778354, 0.1517879, 0.06701052, 0.04088881,
  0.2024251, 0.182828, 0.1030833, 0.1157735, 0.1417542, 0.2183203, 0.1902089, 
    0.08866904, 0.1688438, 0.2002505, 0.2212763, 0.2123963, 0.253125, 
    0.1169321, 0.09646872, 0.144566, 0.2107679, 0.2771822, 0.2140486, 
    0.1437287, 0.09708302, 0.0924142, 0.07587973, 0.08907857, 0.1427906, 
    0.1782154, 0.1558028, 0.1100988, 0.1858404,
  0.1733419, 0.1343289, 0.1585904, 0.1792494, 0.194917, 0.1626009, 0.1429978, 
    0.0825865, 0.08354663, 0.1014388, 0.06469923, 0.05163884, 0.04760919, 
    0.05529116, 0.01197476, 0.06696392, 0.07571307, 0.09864561, 0.1329495, 
    0.1581313, 0.1179232, 0.08212306, 0.06968469, 0.06366789, 0.01486706, 
    0.1410661, 0.2254176, 0.222748, 0.2095442,
  0.0245966, 0.01074533, 0.01513319, 0.03859692, 0.09574513, 0.0335275, 
    0.02954731, 0.01454513, 0.03854714, 0.0133572, 0.01132789, 0.005727855, 
    0.02104112, 0.02482383, 0.1120228, 0.01227868, 0.03731824, 0.03422604, 
    0.03151144, 0.07382964, 0.04428212, 0.009260722, 0.007763017, 0.1395702, 
    0.01318855, 0.02893815, 0.122273, 0.0968466, 0.05318245,
  0.001270608, 0.001366228, 0.01034082, 0.003930437, 0.007941216, 
    0.0005696613, 0.001469299, 0.002513427, 0.005160666, 0.001196918, 
    -9.629705e-06, 4.099732e-08, 0.01265641, 0.002084411, 0.006220329, 
    0.001918947, 0.02758453, 0.03721194, 0.007523206, 0.001064478, 
    0.001641074, 0.0008368678, 0.003140233, 0.01906655, 0.02070818, 
    0.006894146, 0.001744508, 0.0008549078, 0.001479034,
  0.001768884, 0.0272278, 0.00414277, 0.0004430155, -0.001735531, 
    2.197902e-05, 0.0001069457, 0.0003904702, 0.003280228, 0.002647907, 
    0.004473354, 0.001282553, 0.000550916, 0.0002862912, 0.0003787272, 
    0.001996774, 0.0002920913, 9.513598e-05, 3.348634e-06, 1.672096e-06, 
    8.582938e-07, 0.0001064733, 0.002710776, 0.01645747, 0.04546513, 
    0.1232118, 0.0001246204, 1.039752e-05, 8.238434e-05,
  0.01166424, 0.00522978, 0.1057478, 0.07208697, 0.000263938, 0.0001265441, 
    0.0004488403, 9.856051e-05, 0.0004226025, 0.0001301735, 0.0002040158, 
    4.372877e-05, -6.042555e-06, 0.0001529395, 5.397847e-05, 0.000271077, 
    0.0006811998, 0.0002321947, 0.0001245955, 0.0002725377, 0.0005626637, 
    0.002069143, 0.004433976, 0.1131935, 0.07599396, 0.04320728, 
    0.0001421631, 0.0008483317, 0.002795282,
  6.879762e-05, 0.01140657, 0.006184611, 0.00914978, 0.0002806795, 
    0.0004153477, 0.0007715863, 0.0002448067, 0.08486208, 0.1149356, 
    0.0008346504, 0.001029335, 0.0004958443, 4.033074e-05, 0.0004030844, 
    0.0002404612, 8.649097e-05, 0.0003863301, 0.0002507622, 0.0003906697, 
    0.001168725, 0.003733353, 0.008830281, 0.0278251, 0.0312149, 0.004040818, 
    7.530957e-05, 0.0003420966, 0.0004239881,
  5.759461e-09, 4.145226e-09, 7.923849e-10, 0.003272098, 0.002367491, 
    0.0004832021, -0.0004024403, 0.0007179228, 4.232918e-05, 8.18362e-05, 
    0.001224687, 0.0005680584, 0.0005243444, 0.0002645844, 0.0001721072, 
    0.0003382581, 0.0006887718, 0.0002426794, 0.0006381755, 0.0004836691, 
    0.001280354, 0.001186571, 0.1221943, 0.04607373, 7.904445e-05, 
    0.0006091343, 0.001599684, -2.021888e-07, -0.0001368478,
  -1.355854e-10, 1.401473e-09, 6.570423e-10, -6.535026e-05, 6.225227e-09, 
    0.0004556228, 0.0006382465, 0.0007558014, 0.04866432, 0.01524997, 
    0.001286859, 0.001903299, 0.001674647, 0.001421307, 0.0009922346, 
    0.0008780517, 0.0007279413, 0.0004121136, 0.00350351, 0.006328489, 
    0.004396712, 0.06223409, 0.001453919, -0.001195706, 0.0008556247, 
    0.0005224463, 0.0008203438, 4.175008e-05, 3.131189e-09,
  -3.534667e-05, 0.003111568, 0.0002902628, 0.002537589, 0.04977689, 
    -0.001054371, 0.005004631, 0.1016953, 0.01095096, 0.01702197, 0.01191751, 
    0.001938962, 0.002119085, 0.004111916, 0.002903971, 0.003151275, 
    0.00154119, 0.007984052, 0.007076402, 0.01014538, 0.01886568, 0.07754739, 
    0.04756404, 0.002212321, 0.003276826, 0.008906422, 0.001682702, 
    0.005319866, 0.004724144,
  -8.417931e-06, 0.002177098, 0.02258915, 0.2429622, 0.002080277, 0.03566441, 
    0.09012529, 0.003693006, -0.0003173901, 0.01153277, 0.03280086, 
    0.01323135, 0.02374426, 0.03919687, 0.02067356, 0.03481719, 0.02768927, 
    0.04147471, 0.03897242, 0.268165, 0.1066845, 0.03655981, 0.1431271, 
    0.09567156, 0.02543081, 0.03392585, 0.03269562, 0.01649659, 0.06363418,
  0.04421965, 0.2360741, 0.1684291, 0.2714603, 0.1637595, 0.194269, 
    0.02358634, 0.2249249, 0.2088969, 0.08570254, 0.06969053, 0.4457878, 
    0.1231261, 0.08255305, 0.09591463, 0.07689153, 0.09093051, 0.03901308, 
    0.04931368, 0.3997569, 0.1094159, 0.1379866, 0.2046601, 0.3547317, 
    0.1245035, 0.0658425, 0.07385153, 0.028106, 0.02863734,
  0.01835277, 0.3854816, 0.2866822, 0.5010606, 0.5494003, 0.3913451, 
    0.3362578, 0.3197618, 0.471766, 0.433368, 0.4330679, 0.5706968, 
    0.3685231, 0.3338969, 0.1498489, 0.311883, 0.5166655, 0.2703153, 
    0.4211561, 0.4050296, 0.5786675, 0.3190029, 0.1889683, 0.2409953, 
    0.3005614, 0.0277196, 0.06496029, 0.03891117, 0.02747087,
  0.01910986, 0.01716542, 0.360254, 0.05004767, 0.3392227, 0.3460312, 
    0.6290941, 0.4148914, 0.4766485, 0.4078301, 0.5536979, 0.3635474, 
    0.3823926, 0.2439873, 0.2463037, 0.2339019, 0.4553696, 0.3756558, 
    0.1943936, 0.1937041, 0.1536088, 0.2555997, 0.3551404, 0.2544389, 
    0.2174062, 0.2607943, 0.5085396, 0.09806845, 0.06893129,
  0.6665547, 0.6372163, 0.4773426, 0.3542478, 0.3376139, 0.3572395, 
    0.1948959, 0.1721421, 0.2740762, 0.2555507, 0.2418059, 0.3051251, 
    0.3060376, 0.2770521, 0.2904593, 0.2947485, 0.3771445, 0.3022695, 
    0.1947332, 0.2604352, 0.296063, 0.1984071, 0.3689261, 0.4528977, 
    0.1550683, 0.1195659, 0.1109531, 0.2337539, 0.3833161,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, -3.272096e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -2.258097e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, -5.411911e-05, 0, 0.0001237273, 0, -2.996374e-05, 0, 
    -2.129675e-05, 0, 0, 0.001069514, 0, 0.0007197918, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -3.361465e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 2.394752e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, -0.000139622, -2.08553e-05, 0.0002403983, 0, 0.003341083, 0, 
    0.0003061036, 0, 0, 0.00116565, -2.200659e-05, 0.002266245, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 9.5057e-05, -1.858197e-07, 0.0002323879, 0, -5.927597e-06, 
    -2.685445e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.844265e-07, 
    0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -3.291725e-05, 0, 0, -4.962773e-05, 
    3.581404e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, -4.530026e-05, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -9.707285e-06, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, -1.999187e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0.002377653, 0, 0, 0, 0, 0, 0, 0, 0, -1.319825e-05, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, -7.572062e-05, 0, 0, 0,
  0, 0, 3.76484e-05, -0.0001651792, -0.0001322046, 0.0009821514, 0, 
    0.007637457, 0, 0.004323487, -2.25391e-05, 0, 0.00198667, -3.436801e-05, 
    0.003051532, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0003538794, 1.162006e-05, 0, 0, 0,
  0, 0, 0, 0.0008207273, -1.19175e-05, 0.0003888232, -2.211805e-05, 
    0.001100544, -0.0001180158, -1.76594e-05, -9.701998e-06, 0, 0.0001154995, 
    0, 0, 0, -2.010702e-05, -1.513759e-06, 0, 0, 0, 0, 0, -3.7891e-06, 
    -0.0001043366, 0, 0, 0, 0,
  0, 0, 0, 0, 0, -3.359565e-07, 0, 0, 0, 0.0001027106, 0, 0, 3.583495e-05, 
    0.0002923862, 0, 0, 0, -3.609238e-06, 0, 0, 0, 0, 0, -5.366025e-05, 
    0.000226327, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -4.889254e-05, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0.0005302365, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, -5.231447e-08, 0, 0, 0,
  0, 0, 0, 0, 0.006452222, 0, 0, 0, 0, -4.500825e-05, 0, 0, 0, -2.263788e-05, 
    0, 0, 0.0001134566, 0.0004998008, 0.003294205, 2.220525e-05, 0, 0, 0, 0, 
    0, -0.0002423417, 0, 0, 0,
  0, 0, 0.0004822205, 0.001419441, -0.0001749947, 0.003628934, 9.487441e-05, 
    0.01386049, 0, 0.007945134, 1.931894e-05, 0, 0.004480835, 0.0004302075, 
    0.002977256, 0.000201076, 0, -9.562138e-06, 0, 0, 0, 0, 0, 0, 
    0.004211077, 0.001372374, 0, 0, 0,
  0, 0.0006122625, 0.0002166939, 0.002903021, -6.713301e-05, 0.001145215, 
    -3.870659e-05, 0.00367996, 0.0004655358, 0.0002400023, -3.504215e-05, 
    -9.56289e-07, 0.0005892098, -1.275336e-05, 6.729718e-05, 0, 
    -0.0001503981, -3.688515e-05, 0, 0, 0, 0, 0, 2.540032e-05, 0.0001480966, 
    0, 0, 0, 0,
  0, 0, 0, 0, 5.477661e-05, -5.329474e-05, 0, 0, 0.0001911442, 0.001375373, 
    0, 0, 8.869238e-07, 0.003978942, 1.149479e-05, -5.000653e-06, 0, 
    -2.397817e-05, 0, 0, 0, 0, -3.035417e-07, -6.143945e-05, 0.0003993004, 
    -2.406904e-05, 0, 0, 0,
  0, 0, 0, 0, -1.818018e-05, 0, 0, 0, 0, 0, 0.001565164, -0.0001685273, 
    -0.0001037156, 0, 0, 0, -5.576705e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, -1.882614e-07, -2.763422e-07, 0.001832299, 0, 0, 0, 0, 
    -1.833589e-05, 0, 0, -1.610615e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -4.09401e-05, -2.71926e-05, 0, 0,
  0, 0, 0, 0, 0.0211058, 0, 0, 0, 0, 0.0003083376, 0, 0, 0, 0.0004545755, 0, 
    0, 0.002980957, 0.00151052, 0.01349775, 0.0001137508, 0, 0, 0, 0, 0, 
    0.003106933, 0, 0, 0,
  0, 0, 0.0007984476, 0.003559012, 0.0004534899, 0.005098184, 0.0003708061, 
    0.02887917, 0, 0.009787043, 2.733017e-05, 3.557123e-05, 0.01259559, 
    0.001284974, 0.00367805, 0.0009411941, 0, 0.001012743, 0, -4.318381e-05, 
    0, 0, 0, 0, 0.007425166, 0.002346999, 0, 0, 0,
  0, 0.00240534, 0.0007612891, 0.00580663, -0.0003179884, 0.002096667, 
    -1.232743e-06, 0.005187138, 0.003754945, 0.0007932619, 0.002770704, 
    4.127642e-06, 0.001012168, 0.0001939578, 0.003054924, 0, -0.00035309, 
    -5.999386e-05, 0, 0, 0, 0, 0, 0.0001848337, 0.001742691, 0, 0, 0, 0,
  0, 0, 0, 0, 0.0005871342, -5.753078e-05, 4.333173e-07, 0, 0.0002357764, 
    0.009052248, 0, 4.488119e-05, 3.338741e-05, 0.005314807, 3.727938e-06, 
    -7.90307e-06, 0, 6.294787e-05, -3.481988e-05, 0, 0, 0, 2.011487e-05, 
    2.050709e-05, 0.0004560586, -6.400225e-05, 0, 0, 0,
  0, 0, 0, 0, -4.363244e-05, 0, 0, -4.430554e-05, 0, 0, 0.00381616, 
    -0.0002776643, 0.001585661, -2.043815e-06, 0, 0.000739571, 0.0003690057, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -4.395626e-06, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -2.392572e-07, -1.975889e-05, 2.734217e-05, 0.006202423, 0, 0, 0, 0, 
    0.0006315787, 0, 0, 0.001008597, -4.158838e-05, -3.224807e-05, 
    9.495582e-06, -2.590988e-06, 0.001240671, -2.276846e-06, 0, 0, 0, 0, 
    0.0004209879, 0.0007656695, 1.108584e-05, 0, 0,
  0, 0, 0, 0, 0.0480656, -3.647678e-05, 0, 0, 0, 0.0006468108, 0, 0, 0, 
    0.003775577, -1.430597e-05, 0, 0.007350116, 0.002974657, 0.01944494, 
    0.0008376256, 0, 0, 0, 0, 0, 0.008385321, -2.703342e-05, 0, 3.173522e-05,
  0, -6.802623e-05, 0.002199585, 0.01137339, 0.007534923, 0.01454155, 
    0.0007061174, 0.04602658, 0, 0.01168265, -8.569855e-05, 0.0002622688, 
    0.03567641, 0.002751786, 0.005828618, 0.004262169, -2.595025e-05, 
    0.003242763, 0, 0.001108344, 0, 0, 0, -6.811074e-06, 0.0117196, 
    0.004343232, 0, 0, 0,
  0, 0.004933857, 0.001547842, 0.01135398, 0.000261555, 0.007177924, 
    0.0001652168, 0.007542909, 0.008682426, 0.003297984, 0.008117574, 
    -0.0001309802, 0.003759218, 0.0005752886, 0.007367961, -1.643983e-05, 
    -0.0002661871, -9.464402e-05, 0, 0, 0, 0, 0, 0.002319553, 0.004572203, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0.0006610423, 0.004138767, 0.004402874, 1.216247e-05, 
    0.001926066, 0.01552612, -8.687213e-06, 8.426757e-05, 0.0006678827, 
    0.007500239, 0.003238604, -1.502425e-05, 0, 0.0002115382, -9.883933e-05, 
    -1.00127e-05, 0, 0, 6.316555e-05, 0.0002054969, 0.001250239, 
    -0.0001426662, -7.333886e-06, 0, 0,
  0, 0, 0, 0, -7.001153e-05, 0, 0, -0.0001822639, 0, 0, 0.005602339, 
    0.000636235, 0.001393811, 0.000663791, -2.908347e-05, 0.001200073, 
    0.006282111, -2.176523e-05, -2.044404e-05, -8.892867e-05, 0, 
    -9.132321e-05, 0, 0, -3.274322e-07, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.703859e-05, 0, 0, 0, 
    0, 0, 0, 0, -1.197738e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -8.551317e-06, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 1.335843e-05, 1.805111e-05, 0, 0, 0, 0, 0, 0, 4.177674e-05, 0, 
    -3.08146e-05, 0.0003636776, 0.0005647074, 0, 0, 0, 0, 0, 0.001232049, 0, 
    0, 0, 0, 0, -6.795551e-07,
  -3.063633e-05, 0, -5.749137e-06, -2.529054e-05, 0.00581195, 0.01012165, 
    0.0006858496, 0, 0, 0, 0.00362299, 0, 0, 0.006043101, 0.0003531686, 
    8.791346e-05, 0.003436345, -0.0001099371, 0.004426538, 0.0002548445, 0, 
    0, 0, 0, 0.002585299, 0.002846847, -0.0003739538, 0.001378342, 0,
  0, 0, 7.248998e-06, 0, 0.08844204, 0.004818965, 0.001440534, 0, 0, 
    0.001364154, -3.648788e-05, 0, 0, 0.01646808, -6.626015e-05, 0, 
    0.01355486, 0.005866987, 0.02825727, 0.002775763, 0, 0, 0, 0, 
    -0.0001311795, 0.03386584, 0.0008393999, 0, 0.0008250407,
  0, -0.0003245168, 0.00272873, 0.02206809, 0.0201939, 0.03433369, 
    0.001170992, 0.06802332, 0, 0.0168117, -0.0001421591, 0.0006333815, 
    0.05984474, 0.008619494, 0.009226091, 0.01957088, -0.0002253999, 
    0.006036628, 0.003702888, 0.001817483, 0, 0, 0, 0.0006423261, 0.03296691, 
    0.007549216, 0, 0, 0,
  0, 0.006559136, 0.005135134, 0.01828152, 0.005165784, 0.02647823, 
    0.004465272, 0.012325, 0.02293439, 0.007721144, 0.01436605, 0.0005639067, 
    0.008165022, 0.008876716, 0.01920108, 0.0008899248, 0.002843227, 
    0.0002794992, 0, 0, 0, 0, 0, 0.009731987, 0.01186101, 0.0003323308, 0, 0, 0,
  0, 0, 0, 0, 0.003476161, 0.01449849, 0.008767401, 0.0006260711, 
    0.004111971, 0.02214367, 7.523674e-05, 3.127898e-05, 0.008129742, 
    0.01024073, 0.008114811, 3.219305e-05, -5.933337e-05, 0.005346263, 
    -0.0001051618, -8.507293e-05, 0, 0, 0.001317041, 0.004385085, 
    0.004917336, 0.0003764072, -2.243262e-05, 0, 0,
  0, 0, 0, 0, -8.208704e-05, 0, -2.5785e-05, 3.852499e-05, 0, 0, 0.01283632, 
    0.007419048, 0.002199926, 0.006507052, -0.0003452583, 0.002228835, 
    0.01386642, -0.000172641, -0.0001170462, -0.0002404698, -2.84248e-05, 
    -0.0004964496, -3.166035e-07, 0, 5.530625e-06, 0.00186328, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3.013349e-06, 0, 
    -1.562459e-05, -7.214621e-11, 0, 0, -7.375993e-07, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -5.225545e-06, 0.0001701444, 0, 0, 0, 
    5.380872e-05, 0.008772696, -2.827245e-06, 0, 0, 0, 0, 8.46303e-05, 0, 
    0.005918622, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.02174e-05, 0, 0, 
    0, 0, 0.00335158, 0.0002376898, 0.002009035, -1.626434e-05, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -4.16447e-05, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.00516853, -0.0002306234, 
    0.003628255, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  -5.90577e-06, -1.604224e-05, 0, 0.002486607, 0.004481117, 0.002542829, 0, 
    0, 0, 0, 0, 0, 0.001781765, 0.001398816, -0.0001137131, 0.007453722, 
    0.005559548, 0, 0, 0, 0, -4.006502e-05, 0.003224884, 0, 0, 0, 
    0.0001602701, 0.0005831393, -2.323935e-05,
  3.585527e-05, -3.680615e-05, -2.171274e-05, 0.0006608547, 0.02338172, 
    0.01520322, 0.004895156, -2.287695e-05, 0, -1.505243e-06, 0.01046195, 
    -3.422e-05, 0.0006658557, 0.02671613, 0.007086668, 0.009811268, 
    0.008552222, 0.00347367, 0.00772919, 0.00412708, 5.67224e-06, 0, 0, 0, 
    0.005061489, 0.006259201, 0.005362523, 0.002799379, 0.0006891392,
  -3.926164e-05, 0, 0.0004779676, -3.700833e-05, 0.1245132, 0.01092826, 
    0.007169113, -4.301903e-06, 0.01027927, 0.00222026, 0.001022645, 
    -5.227574e-06, -0.0001140512, 0.04833345, 0.001326687, 5.115823e-05, 
    0.02232243, 0.01482236, 0.05043749, 0.004059635, 0, 0, 0, 0, 0.002112177, 
    0.07083741, 0.004890607, 0, 0.006891154,
  3.886502e-06, 0.00291753, 0.005196075, 0.03513964, 0.03161112, 0.06272025, 
    0.0053191, 0.08519811, 1.101209e-05, 0.02759208, 0.01493773, 0.01177724, 
    0.09466433, 0.014109, 0.0169064, 0.04356845, 5.080931e-05, 0.01440127, 
    0.005855237, 0.008420823, 0, 0, 0, 0.003577769, 0.06016842, 0.01124072, 
    0, 0, 0,
  0, 0.01074692, 0.01278077, 0.04268932, 0.02718754, 0.04410405, 0.01516088, 
    0.02110086, 0.05591595, 0.01908281, 0.03121649, 0.01684493, 0.02783467, 
    0.04657789, 0.03921994, 0.004992542, 0.01720743, 0.001095551, 
    -2.130098e-05, 0, 0, 0, 0, 0.08054665, 0.03233108, 0.00200672, 
    0.0001843346, 0, 0,
  0, -1.299359e-05, 0, 0, 0.007321258, 0.02522864, 0.02797648, 0.001854538, 
    0.009612472, 0.03395759, 0.004324893, 0.003257414, 0.03006127, 0.0272182, 
    0.02340527, 0.000198347, -8.360198e-05, 0.01252367, 0.002181988, 
    -0.0001941853, -4.637869e-05, 0, 0.00542245, 0.02784685, 0.02555512, 
    0.00406758, 0.0007163126, 0, 0,
  0, 0, 0, 0, 0.001699383, -1.651948e-06, 0.0001859998, 0.0002692874, 0, 0, 
    0.02687973, 0.01750419, 0.005073487, 0.02414191, 0.001549231, 
    0.003247401, 0.03700129, 0.0001559331, -3.750501e-06, 0.001152621, 
    -0.0003288006, 0.00154817, 0.003658192, 0, 0.0003286453, 0.006455902, 
    -8.003129e-05, -1.584925e-06, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0005827395, 0.0003436318, 
    0.001650015, 0.003404944, 0.001698344, 0.004719097, 0, 0, -0.0001489254, 
    -1.149213e-07, 0, 3.795985e-06, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 2.176365e-05, -1.872809e-05, 0.0006151638, 
    0.0007483537, 0.000234379, 0, 0, 0.001923533, 0.0318419, -2.728329e-05, 
    0, -8.44759e-06, 0.0006806088, 0.003319862, 0.01290503, 0.0001258118, 
    0.01789816, -2.64492e-08, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002717544, 0, 0, 0, -5.822219e-05, 
    6.872793e-06, -1.986431e-05, -6.23227e-05, 0, -2.067594e-05, 
    0.0002330332, 0.009911494, 0.005098997, 0.008112391, 0.001249795, 0, 0,
  -7.510935e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, -9.898938e-05, -1.853812e-05, 0.0008783236, 0, 0.001740339, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, -1.499234e-06, 0, 0, 0, 0, 0, 0, 0, -5.994863e-06, 
    -4.645693e-05, -3.984291e-07, 0.01073912, 0.007241705, 0.0103501, 0, 0, 
    0, 0, 0, 0, 0, -2.231543e-06, -2.138929e-06, 0,
  0.0009008495, 0.0009980954, -2.241884e-05, 0.008652275, 0.01131304, 
    0.007983485, 0.0009908091, 0.003077064, 0.002205631, 0.002580411, 
    0.000459344, 0, 0.01041496, 0.01321495, 0.005659441, 0.01479613, 
    0.008829874, -1.98548e-05, -5.014612e-05, -9.829218e-05, 0, 0.003433067, 
    0.008894831, 0.001032655, -4.484191e-05, -2.972953e-05, 0.002273215, 
    0.003881231, 0.0001561025,
  0.008074108, 0.001479095, -0.0001214462, 0.007465811, 0.03946779, 
    0.02847148, 0.01026948, 0.004154307, 0, 0.0004631863, 0.03264607, 
    0.008022515, 0.005505378, 0.05610051, 0.02063372, 0.03238807, 0.01627953, 
    0.008824287, 0.01106114, 0.01885667, 0.00875949, 0.000768633, 0.00025313, 
    1.410151e-07, 0.01212019, 0.01114735, 0.02590575, 0.01852337, 0.009848475,
  -0.0002039394, -9.919993e-07, 0.01480405, 0.002740702, 0.1837984, 
    0.06720061, 0.02540467, 0.001074484, 0.03005466, 0.00391066, 0.009860504, 
    0.02249618, 0.006384146, 0.117447, 0.01084049, 0.003375661, 0.04521755, 
    0.02961727, 0.07848626, 0.006322858, -6.594276e-06, 7.791258e-05, 
    2.749317e-10, 0, 0.01270641, 0.1275496, 0.01047985, 2.884487e-05, 
    0.02001093,
  0.0005638681, 0.02596518, 0.01316492, 0.1305849, 0.1258456, 0.14493, 
    0.01945161, 0.10849, 0.001898969, 0.07528349, 0.1657932, 0.06096563, 
    0.2366, 0.04240479, 0.05115368, 0.1076373, 0.07618091, 0.06065888, 
    0.01201149, 0.01806879, 4.399919e-09, 2.577823e-06, -2.60416e-05, 
    0.01320351, 0.2394589, 0.01754651, 0.0001352022, -3.889007e-12, 
    -2.689558e-07,
  0, 0.02836096, 0.0605733, 0.1273311, 0.08377281, 0.1291748, 0.06631081, 
    0.1072539, 0.1548773, 0.2338345, 0.1707943, 0.1731222, 0.2445378, 
    0.2691281, 0.1354055, 0.07166168, 0.08714055, 0.03638955, 0.0003537139, 
    0.0003010874, 0, -9.360527e-09, 0.03106296, 0.2256086, 0.1710883, 
    0.00711967, 0.003283761, 0, 0,
  -2.540613e-11, 0.001263013, 0.0001163525, -6.654998e-05, 0.01081133, 
    0.04784959, 0.1211167, 0.03966962, 0.06957307, 0.06665033, 0.0855689, 
    0.07646972, 0.1948351, 0.2071213, 0.06792609, 0.008008951, 0.0002497558, 
    0.03249401, 0.01278339, 0.006753401, -4.600091e-05, 3.935634e-09, 
    0.008366109, 0.1341573, 0.119181, 0.01268187, 0.002770886, 0, 0,
  0, 0, -2.686414e-08, 0, 0.01188566, 0.0006317347, 0.0007672865, 0.01638065, 
    -6.743184e-05, -2.551459e-05, 0.07880585, 0.08082356, 0.06935158, 
    0.05765602, 0.03840086, 0.007023019, 0.07915439, 0.007347216, 
    0.008767538, 0.01300904, 0.0005867226, 0.007861841, 0.009124758, 
    3.813918e-05, 0.0006646822, 0.01388011, -0.0001772213, -4.276794e-05, 
    1.844165e-05,
  -3.173205e-06, 0, 0, 2.898355e-08, 1.663148e-07, 0, 0, 0, 0, 3.519314e-09, 
    1.658865e-08, 1.637225e-07, 4.480599e-08, 1.095432e-06, -1.9363e-09, 
    5.063755e-06, 0.004126613, 0.01179234, 0.01615602, 0.01187644, 
    0.01241414, 0.02017475, -3.659092e-05, -1.598143e-07, -0.0009010612, 
    -7.129517e-06, -2.753523e-09, 0.002592745, 4.628735e-05,
  0, 0, 0, 0, 0, -3.476985e-12, -5.695005e-11, 0, 0, 0.001768461, 
    -0.0001041913, 0.006168092, 0.004380808, 0.005275139, 7.971797e-10, 
    -2.879229e-05, 0.005146589, 0.065708, 0.002740575, -2.750817e-05, 
    -0.0001013401, 0.005409173, 0.008807568, 0.01929629, 0.008543381, 
    0.03052003, 2.531731e-06, -4.916615e-06, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0001164306, 0.01003697, 0, 
    -1.960445e-05, 0.001790328, -0.0002365818, 0.01333513, 0.001597631, 
    0.003861232, 0, -0.0001022466, 0.00628943, 0.01524774, 0.01066898, 
    0.01584942, 0.009257383, 0, 0,
  -4.070537e-05, 0.0009799806, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.820526e-05, 
    0, 0, 0, 0, 0, 0.0008524499, -9.12683e-06, 0, -3.391613e-05, 
    -3.058227e-05, 0.000625517, -9.494871e-05, 0.007285747, 0, 0.007940819, 
    0.00141765,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -8.383953e-06, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  -0.0001104346, 0, -1.129079e-08, 0, 0, -5.752087e-06, 0, 0, -1.621491e-05, 
    -6.413152e-07, 0, 0, 0, 0.0001116215, 0.003162745, 0.005155423, 
    0.02026803, 0.01212072, 0.01825139, -4.472164e-05, 0, 0, -1.256641e-05, 
    0.0002615602, -1.001696e-05, -0.0001334844, 0.0006485218, 0.0006391614, 
    -0.0001620095,
  0.008324857, 0.004674423, 0.0009862063, 0.01419459, 0.01951364, 0.02720945, 
    0.009789402, 0.008841522, 0.004361827, 0.00652744, 0.004467772, 0, 
    0.02523373, 0.02864453, 0.02394071, 0.02513066, 0.02317058, 0.002784106, 
    0.004645813, 0.001997617, -3.943061e-05, 0.0139441, 0.02051608, 
    0.009929686, 0.000238099, 0.00230029, 0.01068136, 0.01720808, 0.00826276,
  0.03734948, 0.01379813, 0.001834172, 0.01929916, 0.09108433, 0.07947812, 
    0.04862032, 0.01733633, -1.642488e-08, 0.006606814, 0.05155347, 
    0.03872884, 0.0130341, 0.09193996, 0.07011394, 0.07693569, 0.04367013, 
    0.02488873, 0.02961779, 0.03502368, 0.04034087, 0.008708108, 0.001797486, 
    0.003039274, 0.0263504, 0.0439085, 0.0957309, 0.06335934, 0.05640273,
  -0.0003498599, 9.665061e-07, 0.1181191, 0.008218151, 0.1704277, 0.08785195, 
    0.1061314, 0.05326154, 0.1224794, 0.02785929, 0.03469955, 0.04528634, 
    0.03626584, 0.2903683, 0.09929576, 0.06841008, 0.1408042, 0.1673349, 
    0.2273838, 0.08134984, 0.001865924, 0.009136318, 0.007111723, 
    -9.153964e-07, 0.1053974, 0.298134, 0.18009, 0.05053977, 0.05000747,
  0.00864227, 0.1274096, 0.07327466, 0.1018122, 0.1159948, 0.1623378, 
    0.0290666, 0.1087475, 0.001826929, 0.05808009, 0.1412531, 0.06196891, 
    0.2069978, 0.03496675, 0.04438787, 0.1043505, 0.1672547, 0.2221749, 
    0.1277646, 0.1494958, 0.0007036671, 0.02710372, 0.0211747, 0.01491775, 
    0.2435531, 0.104607, 0.02633729, 1.498057e-05, -0.0001599321,
  2.148102e-05, 0.09797137, 0.4509045, 0.4208148, 0.1404834, 0.2268252, 
    0.112823, 0.1306355, 0.1641929, 0.2027577, 0.1854454, 0.126179, 
    0.2015142, 0.1982049, 0.1207079, 0.06822289, 0.09780176, 0.04552338, 
    0.02912178, 0.006075441, 0.0001420088, 9.646642e-07, 0.09074508, 
    0.4405788, 0.3283208, 0.15171, 0.1435926, 2.837289e-06, 1.595329e-06,
  5.252999e-06, 0.05589659, 0.1455639, 0.0907541, 0.04003193, 0.1470684, 
    0.2178572, 0.2120367, 0.2824103, 0.2334089, 0.0941575, 0.1279544, 
    0.1959757, 0.1663601, 0.04247936, 0.001009427, 0.000739463, 0.04779259, 
    0.01878845, 0.01962317, 0.01201091, 1.567652e-06, 0.01828187, 0.4393822, 
    0.4349325, 0.1592545, 0.08342532, 5.60369e-06, 5.465924e-06,
  8.432376e-06, 6.678295e-06, 0.0001778191, 9.879303e-05, 0.06159, 
    0.02346136, 0.03652851, 0.03369175, 0.0003805711, 9.509965e-05, 
    0.1038704, 0.08218335, 0.0438039, 0.03900178, 0.03008444, 0.006978344, 
    0.08090642, 0.005701835, 0.04842861, 0.1070644, 0.1276285, 0.04273811, 
    0.01514106, 5.679508e-06, 0.01188644, 0.1201985, 0.1126919, 0.1031646, 
    0.000116827,
  0.000435339, 1.879733e-06, -1.148441e-08, 1.402292e-05, 6.280357e-05, 
    6.608082e-06, -3.915712e-07, 4.07432e-05, 3.561507e-07, -2.076515e-08, 
    2.413336e-06, 7.149153e-08, 6.014609e-07, 1.449882e-06, 1.665089e-07, 
    1.433119e-06, 0.02176002, 0.03944245, 0.02890568, 0.0471262, 0.09025907, 
    0.07010396, 0.01195529, 0.00253842, 0.002259234, -0.0001231927, 
    0.0008683827, 0.05991014, 0.005788839,
  -5.595385e-06, -8.634103e-06, 0.0004294776, 0, -1.522805e-06, 1.707213e-08, 
    0.0002069139, 0, 0, 0.007218728, 0.004515316, 0.01986754, 0.01287783, 
    0.01184666, -6.917636e-05, 0.004271877, 0.01032324, 0.1152258, 
    0.03130846, 0.0003949818, 0.002084436, 0.01496877, 0.01443781, 
    0.02493032, 0.01815823, 0.04120598, 0.002713967, -7.204501e-06, 0,
  0.004043195, 0, 2.799548e-07, 0, 0.0006110424, 0, 0, 0, 0, 0, 0, 
    0.0005622898, 0.01483515, 0.00134837, 0.00340481, 0.005882658, 
    0.006341767, 0.04394829, 0.01440836, 0.02173971, -1.385375e-05, 
    -0.0004307514, 0.01195252, 0.02996548, 0.02300727, 0.0325837, 0.01969177, 
    2.545818e-05, 0,
  0.003121848, 0.003661923, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002418939, 0, 0, 
    0, 0, 0, 0.001272363, -2.637859e-05, 0, -5.836306e-05, -0.0001869469, 
    0.003452125, 0.002501502, 0.01459231, 0.004279483, 0.01711028, 0.00511451,
  6.348469e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, -1.662859e-05, 9.420478e-05, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.064227e-08, 0, -7.708013e-05, 0, 
    -2.449247e-05, -9.609469e-05, -7.35263e-07, -4.294553e-08, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0.001159247, 5.38388e-05, 0.001479909, 0, 0.0001938002, 0.001258941, 
    -7.1727e-05, 0.0001593904, 0.002182918, -0.000108232, 0.002579164, 
    0.006828663, -0.0001352752, 0.0002330353, 0.03409965, 0.04493832, 
    0.04271046, 0.03364615, 0.02457773, -6.547618e-05, -9.763971e-10, 
    -1.441502e-05, -1.663839e-05, 0.005619551, 0.004357354, 0.001134619, 
    0.006249185, 0.006467175, 0.003682728,
  0.04111271, 0.0511591, 0.03478522, 0.05666604, 0.05297447, 0.06361711, 
    0.05597663, 0.03125988, 0.03648434, 0.02688401, 0.04849361, 0.062769, 
    0.04420208, 0.05904024, 0.08788161, 0.1353116, 0.1781022, 0.08875746, 
    0.05320168, 0.02117977, -0.0003269275, 0.0395625, 0.0552818, 0.02296321, 
    0.009800616, 0.02008883, 0.01757671, 0.06685989, 0.06450663,
  0.1486223, 0.08816967, 0.03789948, 0.05017511, 0.1129862, 0.1329419, 
    0.09573328, 0.06541423, 0.05983735, 0.122178, 0.1172433, 0.08751134, 
    0.01810528, 0.1102704, 0.08847878, 0.1184011, 0.1701021, 0.1005233, 
    0.08130215, 0.09388146, 0.1155504, 0.08263843, 0.01550995, 0.004991822, 
    0.04629287, 0.06893416, 0.1250135, 0.08498098, 0.1035956,
  -0.0004775412, 2.480018e-07, 0.1175146, 0.002717054, 0.1650336, 0.08639379, 
    0.1252517, 0.0556235, 0.1124688, 0.02162287, 0.03070797, 0.03193891, 
    0.03338557, 0.2645597, 0.08030929, 0.07588469, 0.1895677, 0.1786557, 
    0.2770336, 0.1977506, 0.08704134, 0.01501924, 0.001625312, 2.406931e-06, 
    0.11079, 0.2822563, 0.1426264, 0.04598917, 0.1207193,
  0.0009717867, 0.08773662, 0.0474956, 0.08227776, 0.09232098, 0.1556288, 
    0.01432758, 0.1232739, 0.002404652, 0.03786289, 0.1275046, 0.0523057, 
    0.1920011, 0.03184209, 0.03945597, 0.1003833, 0.1215241, 0.1736542, 
    0.0996578, 0.1335581, 0.005126518, 0.02091218, 0.008238124, 0.01870791, 
    0.1938431, 0.09269562, 0.005418754, 1.65404e-06, -7.844033e-06,
  3.507315e-05, 0.07229835, 0.426241, 0.3822088, 0.0912622, 0.1649478, 
    0.09032051, 0.09750082, 0.1573198, 0.17403, 0.153074, 0.09803694, 
    0.1419281, 0.1524795, 0.09939783, 0.04731299, 0.06887089, 0.0256847, 
    0.01587547, -0.0001397852, 1.042391e-05, 1.61784e-07, 0.03843822, 
    0.4083462, 0.2953956, 0.1141975, 0.1087031, 1.426024e-06, 2.879889e-07,
  6.98851e-06, 0.02542463, 0.04301178, 0.08257659, 0.0213449, 0.1145392, 
    0.1650631, 0.1508597, 0.2048933, 0.187093, 0.05513107, 0.08743931, 
    0.152683, 0.1333655, 0.03173245, 0.0002968585, 8.213979e-05, 0.02944576, 
    0.006209388, 0.008982552, 0.004904469, 4.500588e-07, 0.006772656, 
    0.243605, 0.3999714, 0.09810504, 0.04938143, 5.680929e-07, 3.804222e-06,
  3.865037e-05, 3.815561e-06, 0.0003455205, 0.001932913, 0.02688344, 
    0.01835621, 0.01627564, 0.02041215, 5.946117e-05, 0.001737875, 0.1071478, 
    0.07764827, 0.02737826, 0.04032518, 0.01314645, 0.006384152, 0.06190987, 
    0.006037584, 0.04517117, 0.06184813, 0.08436423, 0.03381485, 0.01654349, 
    -2.433789e-05, 0.003291376, 0.07214757, 0.09285118, 0.07455061, 
    0.0001142272,
  0.09251171, 0.005847381, -3.074729e-06, 2.488365e-06, 9.446599e-06, 
    5.106575e-06, -2.319236e-07, 3.239654e-05, 2.513862e-07, -1.663877e-08, 
    1.297282e-06, 3.559588e-06, 0.0002040377, 2.127341e-06, 1.478188e-07, 
    -7.484367e-06, 0.01944886, 0.02250157, 0.04359502, 0.05006518, 
    0.06370403, 0.07572227, 0.03568256, 0.03326897, 0.0157334, 1.854023e-05, 
    0.005473372, 0.08329198, 0.1820554,
  0.009912196, 0.001708446, 0.005649833, -1.226003e-10, -6.878132e-05, 
    0.0003207415, 0.003848823, 0, -1.02547e-13, 0.02494233, 0.02521879, 
    0.04902043, 0.04623504, 0.03152, 0.007975429, 0.0314335, 0.03187961, 
    0.1511289, 0.1386244, 0.0352242, 0.012163, 0.05407246, 0.05650939, 
    0.03725016, 0.0572072, 0.06050192, 0.02499298, 0.0001877858, -0.0001791703,
  0.01421863, 0.0003861815, 6.45067e-05, 0, 0.001323291, 0, 0, 0, 0, 0, 0, 
    0.002302856, 0.01894707, 0.01429129, 0.01387281, 0.01613053, 0.03157498, 
    0.07990986, 0.03305155, 0.05446532, 0.00138938, 0.002651501, 0.01964439, 
    0.05618351, 0.03227604, 0.05774442, 0.06143241, 0.01624511, 3.526123e-05,
  0.01408289, 0.005487412, 0, 0, 7.640374e-06, 0, 0, 0, 0, 0, 0, 0, 
    0.007944349, -8.415221e-06, 0.000429515, 0, 0, -1.837907e-05, 
    0.002827574, 0.0006116432, -1.395245e-09, 0.0005761131, 0.0003619326, 
    0.009152109, 0.008763631, 0.02899525, 0.01517062, 0.04905058, 0.01529101,
  0.002215102, -2.933366e-05, -2.423418e-05, 0.0001632842, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -8.702737e-05, 0.0001396386, 
    0.003252119, 0.001191006,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -1.052863e-05, -7.752717e-05, -0.0001126024, 
    -1.738871e-05, 0, 0, -1.34157e-07, 8.491014e-07, 0.0005586476, 
    0.002949284, 0.007390793, 0.003368996, -5.190637e-05, -1.822252e-05, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0.01587776, 0.01202655, 0.01124599, -6.121978e-05, 0.0203152, 0.01531815, 
    0.01031044, 0.008312035, 0.04895558, 0.04213975, 0.04470633, 0.03565496, 
    0.02629138, 0.03190925, 0.09468035, 0.08254689, 0.09692697, 0.07251935, 
    0.05245033, 0.002972257, 0.0004634105, -3.265598e-06, 0.0006607732, 
    0.03693889, 0.03709373, 0.0214366, 0.05333912, 0.05239932, 0.0346312,
  0.09289988, 0.09512857, 0.1131185, 0.1311194, 0.1399589, 0.1581812, 
    0.1069985, 0.1556694, 0.1053223, 0.09260914, 0.1416716, 0.1572557, 
    0.1090295, 0.1142566, 0.1117602, 0.2231621, 0.2051424, 0.132657, 
    0.1276026, 0.1259424, 0.120154, 0.1450762, 0.1156846, 0.05121835, 
    0.1143764, 0.110929, 0.07255638, 0.1014498, 0.1127897,
  0.1201755, 0.1015186, 0.03691269, 0.0448484, 0.07940747, 0.1147828, 
    0.08730992, 0.06957465, 0.05344374, 0.1098924, 0.1090285, 0.1042999, 
    0.02974068, 0.1117758, 0.08906678, 0.1202943, 0.1631528, 0.06857293, 
    0.0725591, 0.09181091, 0.1295685, 0.07760482, 0.02105629, 0.005011449, 
    0.04653744, 0.04927713, 0.1083611, 0.08175838, 0.1028495,
  -0.0004810645, 7.290376e-07, 0.1007907, 0.004047168, 0.1477496, 0.07560984, 
    0.1162269, 0.06294389, 0.09957991, 0.03153817, 0.03735731, 0.02969401, 
    0.03032287, 0.2420373, 0.06932238, 0.06307267, 0.1730089, 0.1488915, 
    0.240963, 0.180679, 0.06167668, 0.005154373, 0.0003317395, -3.663162e-06, 
    0.08272582, 0.2628134, 0.1359765, 0.03035597, 0.1082331,
  0.0004046985, 0.06923097, 0.03718581, 0.07803854, 0.08028354, 0.1402427, 
    0.01518496, 0.1118929, 8.182928e-05, 0.03233862, 0.124366, 0.04977521, 
    0.1717516, 0.02849146, 0.0402789, 0.09548341, 0.1169618, 0.1546564, 
    0.0965345, 0.1120114, 0.01700789, 0.01430953, 0.0001543812, 0.01644027, 
    0.1627461, 0.08407193, 0.002880138, 2.852232e-06, 1.072166e-06,
  5.179232e-05, 0.05088633, 0.3976586, 0.3470675, 0.07893822, 0.1304137, 
    0.08032829, 0.08039802, 0.1550439, 0.1561767, 0.1307052, 0.08430748, 
    0.09232448, 0.1171764, 0.1017706, 0.04724375, 0.06373088, 0.01719701, 
    0.004880185, -5.600378e-06, 6.748819e-07, -1.9065e-08, 0.01753688, 
    0.3934285, 0.2986278, 0.08647166, 0.06654194, 1.129082e-07, 8.465599e-08,
  4.67582e-06, 0.01510493, 0.005527591, 0.02381155, 0.02003435, 0.09210509, 
    0.1419592, 0.1238985, 0.1640968, 0.173371, 0.03770155, 0.06635956, 
    0.1453993, 0.1154085, 0.03005114, 0.000178936, 0.0004536597, 0.01918849, 
    0.004143683, 0.003275255, 0.002260258, 6.556657e-08, 0.004329766, 
    0.1497141, 0.3380229, 0.07328083, 0.02761295, 3.54466e-05, 8.84559e-07,
  7.156361e-06, 2.431823e-06, 7.959936e-05, 0.0007211493, 0.01737997, 
    0.01527287, 0.01094698, 0.01428742, 0.0005561746, 0.004020968, 0.1170854, 
    0.0802846, 0.02459529, 0.03920581, 0.0096949, 0.0109198, 0.05424854, 
    0.01339828, 0.04604274, 0.04630961, 0.05392031, 0.02233714, 0.01353751, 
    1.111669e-05, 0.003688199, 0.04671171, 0.08946379, 0.04668882, 
    3.785257e-05,
  0.09270131, 0.00410516, 9.022731e-07, 3.510054e-07, 2.581591e-06, 
    8.158522e-06, -3.971423e-07, 1.602721e-05, 3.34745e-07, 8.621999e-08, 
    2.040972e-06, 6.524881e-05, 0.008850649, 2.624463e-05, 1.986876e-09, 
    1.271544e-06, 0.01583105, 0.02315039, 0.03416381, 0.02850829, 0.03031629, 
    0.06558285, 0.0261952, 0.03237686, 0.01754059, 0.001286173, 0.02368115, 
    0.1045812, 0.1824106,
  0.03876793, 0.03332373, 0.006254409, 2.966461e-05, 0.004221553, 
    0.003273267, 0.008628499, 0, -2.011852e-12, 0.04959287, 0.07570405, 
    0.07677727, 0.07830505, 0.04202962, 0.0427825, 0.08324278, 0.1062044, 
    0.2556611, 0.2251137, 0.1400378, 0.04992738, 0.1234193, 0.1148249, 
    0.09060817, 0.1221907, 0.06399662, 0.04744172, 0.01427142, 0.01323742,
  0.02446734, 0.00247943, 0.00162301, 0.002622036, 0.00814652, 0.005368438, 
    -5.69439e-05, 0, 0, 0, 0, 0.009275798, 0.03192655, 0.04676123, 
    0.02662031, 0.04332718, 0.06263996, 0.1051097, 0.08289476, 0.09466103, 
    0.004457382, 0.03435196, 0.06797981, 0.1367683, 0.1527365, 0.1381886, 
    0.1239503, 0.04637093, 0.004261091,
  0.06739099, 0.01111369, 0.0010968, 6.508097e-05, 0.00174711, 0, 0, 0, 0, 0, 
    0, 0, 0.01677228, 0.00252511, 0.001426086, 0, -4.00912e-11, 0.000112867, 
    0.01100993, 0.01100425, 7.881057e-05, 0.005806797, 0.009694689, 
    0.01760655, 0.01886288, 0.04442019, 0.04405819, 0.07576872, 0.06366943,
  0.01335698, 0.0008889289, 0.003599317, 0.002907537, 0.0007921132, 0, 0, 0, 
    0, 0, 0, 0, -1.558891e-05, -2.41e-06, 0, 0, 0, 0, 0, 0, 1.273597e-10, 0, 
    0, 0, -1.240673e-05, 0.000326067, 0.006208509, 0.008249831, 0.00368519,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  -6.563026e-06, -3.679191e-05, 0, -4.705772e-07, -7.98687e-05, 0, 
    0.0003335318, 0.00235116, -2.529244e-05, -0.00181598, -4.510734e-05, 
    -2.223118e-07, -0.0003526684, -0.0008569325, 0.04029131, 0.03862963, 
    0.02390742, 0.02373825, 0.01639991, 0.005061181, 0, -1.277549e-05, 0, 
    -1.081034e-05, 8.988622e-06, 0.00172677, -1.612686e-07, 0, -1.556543e-05,
  0.06576779, 0.0465058, 0.02536052, 0.04522037, 0.03645819, 0.04848013, 
    0.03055512, 0.03975983, 0.1183102, 0.1379955, 0.1202774, 0.1485344, 
    0.150357, 0.1347435, 0.1497031, 0.1122078, 0.1262641, 0.09462484, 
    0.08362702, 0.05468964, 0.04018242, 0.03921551, 0.02908964, 0.07451517, 
    0.07596759, 0.09596148, 0.121863, 0.1387547, 0.07867461,
  0.1340225, 0.1280567, 0.1642371, 0.1862919, 0.1997954, 0.1878725, 
    0.1550836, 0.1653398, 0.1292325, 0.1530821, 0.1617389, 0.1588539, 
    0.1597891, 0.1452382, 0.1081774, 0.2052433, 0.1802914, 0.126142, 
    0.1331419, 0.1335519, 0.1702291, 0.1790782, 0.1544412, 0.09723771, 
    0.127108, 0.1478099, 0.09013153, 0.1122114, 0.1467987,
  0.09639008, 0.08851001, 0.03079683, 0.03522561, 0.07007569, 0.1203435, 
    0.06974157, 0.06419558, 0.03070108, 0.08337946, 0.07809108, 0.09882882, 
    0.03556591, 0.09503783, 0.09040376, 0.1103568, 0.1559446, 0.04339304, 
    0.07531261, 0.09819436, 0.1131464, 0.05435019, 0.02778942, 0.00348511, 
    0.04591187, 0.03566919, 0.0898113, 0.08388876, 0.07932371,
  -0.0002047384, 5.852665e-08, 0.09799288, 0.01998956, 0.1393365, 0.05786959, 
    0.1063546, 0.04754244, 0.09916948, 0.02714971, 0.03648791, 0.02475826, 
    0.02477132, 0.2287961, 0.06647161, 0.0503512, 0.152044, 0.1135351, 
    0.1929532, 0.188198, 0.03629482, 0.003945613, 3.565628e-05, 
    -4.905385e-07, 0.06328368, 0.2415418, 0.1542609, 0.03055174, 0.09145534,
  2.933219e-05, 0.05158447, 0.0310126, 0.06506511, 0.08780868, 0.11786, 
    0.01275168, 0.1160779, 3.306096e-05, 0.03211314, 0.1317618, 0.04676847, 
    0.1580265, 0.02382213, 0.04255847, 0.08366286, 0.09966595, 0.1392646, 
    0.08724342, 0.1032475, 0.002456968, 0.01186936, 6.924375e-05, 0.012025, 
    0.1280656, 0.07942016, 0.002211369, 3.278255e-06, -2.21539e-08,
  3.251416e-05, 0.04527751, 0.3785273, 0.3013668, 0.07344866, 0.1011025, 
    0.08030184, 0.07001932, 0.1454978, 0.1351626, 0.1168471, 0.07801716, 
    0.06099927, 0.08915821, 0.1062955, 0.03991392, 0.05777223, 0.01149858, 
    0.003263826, 5.601757e-05, 2.380712e-07, -1.474479e-08, 0.01039872, 
    0.3457841, 0.2975983, 0.04667817, 0.02406931, -7.601963e-08, 2.845454e-09,
  1.965185e-06, 0.01179098, 0.004132214, 0.005509551, 0.02282284, 0.06608324, 
    0.107205, 0.0961953, 0.1160959, 0.1553001, 0.02018913, 0.046619, 
    0.1208724, 0.09141962, 0.02943046, 0.0002857428, 2.306696e-05, 
    0.01301392, 0.01852066, 0.001570437, 0.001220605, 6.682246e-08, 
    0.004322428, 0.07653262, 0.2506104, 0.07890029, 0.01995216, 0.0002965997, 
    8.02392e-07,
  2.427928e-06, 9.224268e-07, 6.293084e-06, 0.0004269296, 0.0131894, 
    0.009300324, 0.004604129, 0.01103857, 0.00117681, 0.0004594948, 
    0.1147772, 0.07328223, 0.01606741, 0.03710585, 0.006992077, 0.01659972, 
    0.05668736, 0.02483736, 0.02811787, 0.04261469, 0.03831118, 0.00296192, 
    0.02245781, -2.500656e-05, 0.005297956, 0.0437538, 0.08065422, 
    0.01979172, 4.380695e-05,
  0.09922805, 0.002274069, -1.454441e-06, 9.821814e-08, 7.554221e-07, 
    1.739011e-05, -4.225948e-07, 4.0482e-06, 3.694933e-07, 1.328771e-07, 
    4.788392e-06, 0.0003117161, 0.00191252, 6.370507e-05, -1.016163e-06, 
    8.999576e-06, 0.02378794, 0.02008492, 0.01625758, 0.03328979, 0.01911413, 
    0.05070261, 0.01786575, 0.03378244, 0.01540903, 0.003765648, 0.05888227, 
    0.074196, 0.1675424,
  0.06621592, 0.07801828, 0.03142456, 0.009567959, 0.008440387, 0.03566212, 
    0.02230731, -1.839235e-09, -4.471835e-07, 0.1225206, 0.1286068, 
    0.08037799, 0.07327583, 0.0508622, 0.07470124, 0.1131981, 0.1568574, 
    0.2405815, 0.1748061, 0.09204043, 0.09086058, 0.1071571, 0.1151206, 
    0.06965666, 0.08828245, 0.06496408, 0.03267191, 0.02272821, 0.01533672,
  0.02856591, 0.02306588, 0.003744179, 0.01702759, 0.01093108, 0.009940441, 
    -0.0001218913, 0, 0, -5.642944e-13, -2.549104e-05, 0.0362652, 0.07841018, 
    0.09226692, 0.06419972, 0.08129597, 0.1335164, 0.1698526, 0.1621892, 
    0.1313187, 0.01423014, 0.1424102, 0.162056, 0.2233273, 0.1885908, 
    0.1929071, 0.1668646, 0.1011915, 0.05343832,
  0.1027685, 0.02963194, 0.001151703, 0.007234456, 0.005884439, 0, 0, 0, 0, 
    0, 0, 0, 0.01809102, 0.01871566, 0.02851608, 0.005461233, -8.671924e-08, 
    0.003326823, 0.04062655, 0.02580463, 0.005438676, 0.04312821, 0.0647551, 
    0.04291825, 0.08781707, 0.1171219, 0.1098337, 0.141566, 0.1060358,
  0.04937569, 0.02526095, 0.0120631, 0.01301744, 0.001798001, -5.205464e-06, 
    0, 0, 0, 0, 0, -3.178459e-06, -0.0001794769, 0.007762837, 0.007225167, 
    8.106412e-08, -5.649851e-06, 0.0003500416, -4.489512e-06, -3.961856e-05, 
    0.00173532, 0, 3.188418e-07, -1.720246e-08, 0.002235915, 0.006167639, 
    0.01596685, 0.02079183, 0.03365774,
  0.0008265651, -9.480867e-05, 0, -1.610135e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.49135e-05, 0.001879085,
  -1.817017e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.0005189393,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0006144099, -0.0003167927, 
    0, 0, 0, 0, 0, 0, -3.895277e-05, 0, -4.111895e-07, 0, 0, 0,
  0.03459467, 0.02125119, 9.389594e-05, -7.895546e-06, -0.0004505037, 
    -0.000474179, 0.01935699, 0.003360037, 0.009876738, 0.01189599, 
    0.00621233, -0.0001951875, 0.001220295, 0.01434648, 0.0737502, 0.1087505, 
    0.1850141, 0.1455784, 0.1532465, 0.06999953, 0.05300339, 0.02330501, 
    0.008993748, 0.01191343, 0.1076299, 0.09177702, 0.014086, 0.006442958, 
    0.007496447,
  0.128238, 0.07964644, 0.04757223, 0.08696281, 0.1008617, 0.09260178, 
    0.09688887, 0.113355, 0.163528, 0.1845594, 0.2157221, 0.1893965, 
    0.1809142, 0.1647079, 0.1886483, 0.1227429, 0.1164676, 0.09763226, 
    0.1263813, 0.1001446, 0.07738008, 0.0614754, 0.07740041, 0.1635237, 
    0.143259, 0.1132991, 0.1597937, 0.1710874, 0.1392372,
  0.1633353, 0.1869826, 0.2129694, 0.1803404, 0.1873605, 0.1691696, 
    0.1485902, 0.1657921, 0.1512759, 0.1821077, 0.1407793, 0.1490885, 
    0.1943112, 0.1752661, 0.09755322, 0.1917533, 0.1551421, 0.125085, 
    0.1336938, 0.141627, 0.1568224, 0.1654869, 0.1492806, 0.09883599, 
    0.1175095, 0.1550542, 0.09264076, 0.1130825, 0.1698591,
  0.08048245, 0.08256321, 0.03022206, 0.03950936, 0.06381069, 0.1132384, 
    0.06149534, 0.05494503, 0.02001185, 0.06798165, 0.05829581, 0.08216311, 
    0.03732301, 0.08905571, 0.08939298, 0.09762971, 0.1315477, 0.0266253, 
    0.08165909, 0.1082328, 0.1043592, 0.06265043, 0.02592651, 0.003164902, 
    0.04766512, 0.02859673, 0.06853034, 0.0831747, 0.05590659,
  0.00175335, -8.556468e-07, 0.08783845, 0.005079478, 0.1383863, 0.05850988, 
    0.09760801, 0.04481454, 0.05679426, 0.03926296, 0.03953752, 0.0137648, 
    0.01946113, 0.2117058, 0.07892939, 0.03094626, 0.1499665, 0.09293534, 
    0.1757939, 0.1970556, 0.01869132, 0.004337875, 1.068798e-06, 
    -2.763474e-06, 0.05581819, 0.2207308, 0.1316096, 0.0181517, 0.08248125,
  1.263201e-05, 0.04604963, 0.02507539, 0.05561918, 0.09437575, 0.1066852, 
    0.007165831, 0.116461, 7.701742e-05, 0.02921865, 0.09731879, 0.03700819, 
    0.1462921, 0.01795842, 0.04312927, 0.07709786, 0.0840052, 0.1141508, 
    0.06944415, 0.08304746, 0.0001024737, 0.00682571, 4.743041e-05, 
    0.0105196, 0.113851, 0.0567187, 0.001890923, 1.927297e-06, 3.908782e-08,
  1.209947e-05, 0.03426908, 0.3290854, 0.2479399, 0.05587196, 0.07589347, 
    0.06498481, 0.06106403, 0.1286652, 0.1203606, 0.09619172, 0.0741355, 
    0.04632069, 0.0574539, 0.1103071, 0.02470548, 0.04126654, 0.009646465, 
    0.003111193, 5.530024e-05, 8.848299e-10, -2.289552e-08, 0.003541253, 
    0.2851835, 0.2775128, 0.02974604, 0.01518401, -3.659473e-07, -4.410834e-09,
  -4.138655e-06, 0.01142329, 0.004152327, 0.0009491846, 0.02222469, 
    0.03797492, 0.07436397, 0.06270672, 0.07172848, 0.1463019, 0.01189991, 
    0.03280012, 0.09776457, 0.06109616, 0.02327422, 0.0007731015, 
    0.0004339143, 0.013845, 0.01718077, 0.0009584669, 0.0005502804, 
    -6.157323e-09, 0.02737316, 0.04454075, 0.1607011, 0.06914006, 0.01321067, 
    0.0003589458, 1.004182e-06,
  7.389472e-07, 3.635256e-07, 2.736778e-06, 0.0005482589, 0.007312596, 
    0.004741491, 0.005122755, 0.005117676, 0.0009009153, 0.0008443053, 
    0.09513982, 0.06737929, 0.01347999, 0.03806718, 0.006569139, 0.01834323, 
    0.05494983, 0.0365609, 0.02175673, 0.0300282, 0.02494808, 0.002629773, 
    0.007779478, 0.0001999014, 0.006072612, 0.04017913, 0.07006778, 
    0.01995945, 1.557447e-05,
  0.104755, 0.001570084, 0.0003776563, -1.28158e-06, 8.573867e-07, 
    1.963826e-05, -5.571881e-07, 1.514914e-06, 4.603643e-07, 4.184719e-08, 
    4.545489e-05, 0.001229386, 0.0001433319, 0.005888492, 0.0009736831, 
    0.005028641, 0.03113517, 0.01909636, 0.008131569, 0.041411, 0.01465223, 
    0.04728474, 0.007136223, 0.03554828, 0.01397578, 0.006992743, 0.03799325, 
    0.05296183, 0.1621747,
  0.03629752, 0.06890281, 0.03402162, 0.02447532, 0.011224, 0.04264117, 
    0.02854699, -2.596605e-08, 0.0001833038, 0.1581109, 0.1639892, 0.0886275, 
    0.06594313, 0.05826949, 0.08203864, 0.1195935, 0.1398848, 0.1668225, 
    0.1425823, 0.07535032, 0.09698217, 0.08780514, 0.1102433, 0.05423359, 
    0.074312, 0.05803533, 0.02204934, 0.02386277, 0.009743251,
  0.05985591, 0.08796176, 0.05912701, 0.05698038, 0.008864018, 0.01203283, 
    0.0003212407, 0.001215109, -5.199379e-07, -6.267042e-09, 0.004297975, 
    0.09063438, 0.1133279, 0.1291053, 0.132985, 0.1204073, 0.1859971, 
    0.2018835, 0.176421, 0.2206331, 0.05996671, 0.1603387, 0.1812555, 
    0.2101689, 0.1830041, 0.176076, 0.1620932, 0.1131029, 0.1093447,
  0.1732879, 0.110167, 0.08265769, 0.05483398, 0.03863671, 0.00577673, 0, 
    -1.0136e-05, 0, 0, 0, 0, 0.09399832, 0.06060178, 0.08886948, 0.04815042, 
    0.004334344, 0.01039274, 0.1075744, 0.04648835, 0.03768608, 0.09449413, 
    0.1584347, 0.1267491, 0.1976124, 0.1616301, 0.1284032, 0.1666798, 
    0.1759849,
  0.09628871, 0.09690259, 0.0573087, 0.03780044, 0.004175424, 0.0003343763, 
    1.942814e-05, -5.43819e-09, 0, 0, 0, -1.271384e-05, 0.002493357, 
    0.01894291, 0.01561236, 0.02946636, -0.0001180529, 0.001666655, 
    0.000450979, 0.004512607, 0.02628012, 0.02552105, 0.02511886, 0.00138609, 
    0.01606998, 0.02154415, 0.02834799, 0.03974297, 0.08543134,
  0.006146032, 0.009030391, -0.0003220982, 0.0006859038, 0, -5.18946e-05, 
    -3.532122e-05, 0.00276775, 0, 0, 0, 0, -3.269555e-05, 0.02285318, 
    0.05863459, 0.03139314, 0.03107483, -1.028494e-05, 1.483986e-07, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.0002124823, 0.009763707,
  -3.089996e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, -6.280977e-05, 0.0008760073,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.671277e-07, 0.00143072, 
    0.01081199, 0.09872597, 0.06934932, 0.004021883, 0, -4.370186e-06, 0, 
    0.004400969, 0.03411278, 0.00390594, 0.00895083, 0.006083048, 
    -1.650017e-05, 0,
  0.1953449, 0.07802235, 0.06331675, 0.02662629, -0.000496955, 0.003743013, 
    0.09095066, 0.005025927, 0.04455578, 0.07023378, 0.03321811, 
    -0.0005018571, 0.0117667, 0.07957537, 0.1238611, 0.1635115, 0.1998932, 
    0.1885769, 0.1896924, 0.09925342, 0.08240724, 0.07208484, 0.06166219, 
    0.1627249, 0.3181249, 0.2245979, 0.06855676, 0.04989437, 0.1706473,
  0.1765465, 0.1210613, 0.1200288, 0.1708492, 0.1850464, 0.1256945, 
    0.1779299, 0.2096881, 0.2303224, 0.2655971, 0.2435735, 0.1811553, 
    0.1744763, 0.1733405, 0.1634239, 0.1192598, 0.1133788, 0.1109223, 
    0.1539535, 0.1858898, 0.1504303, 0.1144149, 0.151699, 0.2392764, 
    0.2355448, 0.1703209, 0.199864, 0.1935605, 0.2068974,
  0.1870947, 0.2086738, 0.2225161, 0.1739268, 0.1763288, 0.153316, 0.1329262, 
    0.1624149, 0.1552642, 0.1675805, 0.154162, 0.1316644, 0.1833621, 
    0.1741237, 0.09697621, 0.1786592, 0.1459489, 0.1310107, 0.1335105, 
    0.1524365, 0.1499466, 0.1585101, 0.1396239, 0.09342858, 0.09734552, 
    0.1474919, 0.1071433, 0.1292048, 0.1815072,
  0.07449353, 0.07065284, 0.02509777, 0.03858677, 0.0569164, 0.1061375, 
    0.07216921, 0.05957055, 0.01187736, 0.04632375, 0.0366033, 0.07710803, 
    0.03977054, 0.08762643, 0.08360616, 0.1144419, 0.09994626, 0.02461576, 
    0.0756292, 0.07620493, 0.07928319, 0.07134674, 0.02564893, 0.00211122, 
    0.04734675, 0.02790223, 0.04965219, 0.07402315, 0.04687364,
  0.004141381, -7.673587e-07, 0.08054509, 0.002502914, 0.1371855, 0.04611719, 
    0.09288184, 0.03180651, 0.04040518, 0.04222661, 0.04330684, 0.0154172, 
    0.0179904, 0.1962256, 0.08140107, 0.02639109, 0.1550402, 0.08370283, 
    0.1506421, 0.1402352, 0.01114818, 0.002913765, 2.327852e-07, 
    -7.44892e-06, 0.05384937, 0.2245324, 0.09064846, 0.01050451, 0.07270946,
  3.36725e-05, 0.03969544, 0.02337503, 0.06762379, 0.1178021, 0.09893447, 
    0.007205699, 0.1193971, 0.000181483, 0.02457653, 0.06888177, 0.0268848, 
    0.1322623, 0.01634923, 0.05446432, 0.07205801, 0.06455392, 0.09396136, 
    0.04985595, 0.06893735, 1.893443e-05, 0.002711044, 6.045397e-06, 
    0.01013605, 0.09973177, 0.04261049, 0.001404236, 2.498469e-07, 
    1.617834e-07,
  4.515652e-06, 0.02477595, 0.2726038, 0.1707915, 0.04443996, 0.05307323, 
    0.0661896, 0.05843472, 0.09947816, 0.1022891, 0.0818511, 0.06976558, 
    0.04152808, 0.03758474, 0.1111697, 0.01726148, 0.03591143, 0.008867031, 
    0.002893823, 8.883686e-05, 0, 1.903568e-08, 0.0005011407, 0.2202734, 
    0.2613218, 0.02664553, 0.01001952, -2.322476e-06, 8.613269e-08,
  2.003845e-05, 0.008261035, 0.004336298, 0.000529229, 0.02364078, 
    0.03910206, 0.06482847, 0.04814348, 0.04675405, 0.1408549, 0.009232153, 
    0.02135993, 0.07602526, 0.04417401, 0.01537, 0.005106878, 0.0005393783, 
    0.01268058, 0.01670766, 0.0001622976, 0.0007730412, 1.240641e-07, 
    0.04313658, 0.036305, 0.09710519, 0.04915965, 0.01275177, 0.000358476, 
    4.095707e-06,
  1.760384e-07, 7.542698e-08, 7.86637e-07, 0.001416223, 0.001922678, 
    0.002045488, 0.002172835, 0.00295508, 0.0009562274, 0.0008104014, 
    0.08752988, 0.06032872, 0.01234896, 0.0359485, 0.02624881, 0.01628638, 
    0.05883914, 0.04420496, 0.02254459, 0.01193075, 0.02175939, 0.002185812, 
    0.001494353, 0.0003580921, 0.008609345, 0.03944426, 0.0345605, 
    0.02269457, -6.669966e-05,
  0.0790977, 9.644464e-05, 2.675584e-05, -3.567777e-06, 5.138106e-07, 
    2.085997e-05, -8.096393e-07, 4.321122e-07, 1.37014e-07, 8.773588e-08, 
    0.0004348326, 0.005156998, 1.860224e-05, 0.004356022, 0.005608141, 
    0.02737649, 0.02278053, 0.01298956, 0.003676907, 0.04366443, 0.01784534, 
    0.04122989, 0.003289162, 0.01962992, 0.01229885, 0.007847997, 0.01092268, 
    0.03618165, 0.1155866,
  0.02509058, 0.05530812, 0.03746093, 0.03400824, 0.01416911, 0.04533198, 
    0.03203595, 6.510091e-06, 0.003662994, 0.178648, 0.1959582, 0.08259467, 
    0.06921794, 0.08309145, 0.09210625, 0.1251226, 0.1337691, 0.1442744, 
    0.1294161, 0.0666451, 0.08736241, 0.07691738, 0.08283915, 0.03740831, 
    0.0609137, 0.05334228, 0.01806797, 0.01536298, 0.01236997,
  0.06659113, 0.09403037, 0.05771724, 0.06013863, 0.08060235, 0.04691376, 
    0.008366188, 0.05442159, 0.005345318, -0.0003134079, 0.03891735, 
    0.1269576, 0.1606981, 0.1312222, 0.1298761, 0.1316264, 0.2413525, 
    0.2128279, 0.187831, 0.2456632, 0.1677203, 0.1622011, 0.1799991, 
    0.2034592, 0.1491921, 0.1569349, 0.1678696, 0.09918685, 0.08948299,
  0.1858682, 0.1727403, 0.1584661, 0.166154, 0.1575465, 0.1603722, 
    0.04158422, -4.397566e-05, 0.0002346785, 0, 4.244074e-07, -0.0007591399, 
    0.1653284, 0.1296173, 0.1518463, 0.1035114, 0.077721, 0.01764932, 
    0.1405371, 0.09089869, 0.05966368, 0.1136104, 0.2073645, 0.1928296, 
    0.2077682, 0.15692, 0.1364251, 0.1842754, 0.1876148,
  0.1473716, 0.135763, 0.1248378, 0.1370757, 0.1289417, 0.04540066, 
    0.03243283, 0.01181833, 0.01087083, 0.00234237, 0, 8.942423e-05, 
    0.01527306, 0.1050356, 0.05091997, 0.0151748, -3.911937e-05, 0.007123931, 
    0.003757621, 0.02752782, 0.05320338, 0.08454469, 0.05750172, 0.05258003, 
    0.05460559, 0.04141209, 0.05704262, 0.1028686, 0.1269686,
  0.05378, 0.02148069, 0.0006606919, 0.02210126, 0.01612856, 0.02307249, 
    0.01647369, 0.006456678, 0, 0, -2.865961e-07, -6.641282e-05, 0.03023269, 
    0.11672, 0.08839456, 0.06767986, 0.06972051, 0.07003356, -9.995805e-05, 
    0, 0, -2.177763e-10, 0, 0, 0.002218597, 0, -1.21052e-05, 0.009710737, 
    0.04649156,
  0.000965354, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, -6.821496e-06, 3.325992e-05, -2.454268e-05, -0.000623417, 
    0.007054899,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001714159, 0.006405239, 0.1073702, 
    0.1886564, 0.2628158, 0.1593984, 0.009979841, 0.0005855021, 
    -0.0003289302, 0.02748275, 0.08685387, 0.0462179, 0.02404216, 0.05787311, 
    -0.002544805, 0,
  0.2194079, 0.192568, 0.1437881, 0.1435035, 0.003630867, 0.01621077, 
    0.1623148, 0.01407163, 0.09139539, 0.10059, 0.0786046, 0.01865013, 
    0.06830983, 0.1159926, 0.1567929, 0.1809673, 0.2021642, 0.2156147, 
    0.2226384, 0.1306447, 0.09155595, 0.1433545, 0.2267918, 0.2257865, 
    0.4023888, 0.2265963, 0.1142833, 0.1545323, 0.2248119,
  0.2114569, 0.1542712, 0.1722978, 0.2406655, 0.2109549, 0.1277052, 
    0.1837872, 0.2211422, 0.2628506, 0.2734823, 0.2394244, 0.1918194, 
    0.1559485, 0.173477, 0.1692322, 0.121194, 0.1139357, 0.1230281, 
    0.1654652, 0.203073, 0.183151, 0.1869314, 0.1720638, 0.2328168, 
    0.2542095, 0.1782759, 0.2047081, 0.2207999, 0.2479151,
  0.1922873, 0.2130446, 0.2280847, 0.1767762, 0.1759439, 0.1714887, 
    0.1257831, 0.167166, 0.1504177, 0.1548098, 0.1546986, 0.1109716, 
    0.1747207, 0.160732, 0.1003524, 0.1867395, 0.1466828, 0.133211, 
    0.1216701, 0.1414014, 0.1290968, 0.1489033, 0.1429073, 0.09147725, 
    0.09609959, 0.143264, 0.09529038, 0.134426, 0.1939831,
  0.07286762, 0.06991953, 0.01966506, 0.04355116, 0.06659491, 0.1059662, 
    0.06457753, 0.05334185, 0.01672283, 0.03627776, 0.0272168, 0.06836623, 
    0.04402125, 0.08111182, 0.07825907, 0.1327444, 0.08126707, 0.01182513, 
    0.06327949, 0.08072425, 0.07595791, 0.06691664, 0.01544669, 0.002505168, 
    0.05057789, 0.03179954, 0.04154234, 0.06818713, 0.04675823,
  0.004169963, -2.736528e-07, 0.06120417, 0.0005407056, 0.1458168, 
    0.02250394, 0.07236256, 0.02787085, 0.01941409, 0.04305778, 0.04109174, 
    0.01916333, 0.02143752, 0.1854071, 0.0641252, 0.01877149, 0.1566852, 
    0.08376282, 0.1424706, 0.1051547, 0.00748039, 1.990996e-06, 4.134349e-08, 
    -1.502931e-05, 0.05242588, 0.2405678, 0.06406946, 0.005779244, 0.06960644,
  0.002090645, 0.02334887, 0.02181681, 0.05676615, 0.1204527, 0.09536474, 
    0.007050158, 0.1169932, 0.001489853, 0.02560762, 0.05602635, 0.02334483, 
    0.1116157, 0.02136029, 0.06171366, 0.06926391, 0.05332044, 0.09104003, 
    0.04246231, 0.0589195, 1.002714e-07, 0.001452442, 1.955292e-07, 
    0.009403493, 0.09732907, 0.03786608, 0.001281845, 1.645956e-07, 
    2.559701e-07,
  2.839904e-06, 0.02017495, 0.242268, 0.1373494, 0.04652877, 0.05311661, 
    0.06990047, 0.06070928, 0.0731971, 0.07970616, 0.0689002, 0.0728531, 
    0.0446034, 0.0342876, 0.1045664, 0.01224273, 0.03164884, 0.007735609, 
    0.003047962, 0.0003321506, 0, 1.211181e-08, 5.32195e-05, 0.1924099, 
    0.2787393, 0.02758935, 0.006487658, 0.0004267512, 1.773707e-07,
  0.0002354082, 0.009826995, 0.003947567, 0.0007396432, 0.02370111, 
    0.03224618, 0.0484455, 0.04780617, 0.05216021, 0.1418516, 0.007841947, 
    0.01185808, 0.05562796, 0.03543484, 0.01408551, 0.005009647, 0.003568061, 
    0.01392576, 0.007492846, 0.0004833578, 0.0006848858, 1.51294e-07, 
    0.04366832, 0.03817132, 0.06961384, 0.03932967, 0.01850178, 0.002147632, 
    3.903467e-05,
  -4.973256e-07, 2.89606e-07, 7.596989e-07, 0.002796972, 0.0008178909, 
    0.001994055, 0.001171626, 0.001277198, 0.001315329, 5.369244e-05, 
    0.07426969, 0.0572823, 0.01022676, 0.04514659, 0.02968305, 0.02266561, 
    0.06622557, 0.056995, 0.02784559, 0.007203711, 0.033399, 0.002963014, 
    0.00240886, 0.0004113995, 0.01867687, 0.0508102, 0.04145262, 0.01445399, 
    0.0004046349,
  0.01977995, -1.484911e-06, 2.99539e-08, -1.880542e-07, 4.568049e-07, 
    8.472651e-06, -2.208998e-07, 2.605938e-07, 1.859447e-07, 1.372366e-07, 
    0.00100075, 0.01157991, 0.001972957, -2.612627e-05, 0.008260801, 
    0.02784623, 0.01314664, 0.001276694, 0.0005222798, 0.04445795, 
    0.007327382, 0.03795604, 0.004558052, 0.0132829, 0.01472749, 0.01152677, 
    0.0005892243, 0.03336117, 0.1010447,
  0.01790618, 0.0426212, 0.03275784, 0.02670412, 0.01564329, 0.04665937, 
    0.03154207, 0.0008103551, 0.01171777, 0.1986849, 0.2147894, 0.0915044, 
    0.08090814, 0.09300306, 0.09373606, 0.1154884, 0.1276738, 0.1485311, 
    0.1066493, 0.04488644, 0.07170977, 0.07348578, 0.04960564, 0.02801501, 
    0.05135719, 0.04953488, 0.01376994, 0.01494121, 0.01591453,
  0.066976, 0.07883254, 0.06283805, 0.06030928, 0.05143154, 0.05691547, 
    0.02090394, 0.1178527, 0.06414376, 0.04537293, 0.05613339, 0.1678612, 
    0.166627, 0.1314605, 0.1321711, 0.1623568, 0.246027, 0.2084647, 
    0.1894316, 0.2405482, 0.2133319, 0.1676116, 0.1839661, 0.181793, 
    0.1273269, 0.1736836, 0.1737223, 0.1049049, 0.1166071,
  0.1801694, 0.232406, 0.1429469, 0.1825467, 0.1708571, 0.1715154, 0.1833024, 
    0.002717014, 0.0007358745, -0.0001635334, 0.007406804, 0.07421234, 
    0.1987048, 0.1923441, 0.3092076, 0.1682602, 0.08576909, 0.0161251, 
    0.1364564, 0.1203933, 0.08801471, 0.140716, 0.2302064, 0.2121148, 
    0.2286438, 0.1669556, 0.1476021, 0.201663, 0.1941933,
  0.1738838, 0.1610279, 0.1976182, 0.187489, 0.2618354, 0.181169, 0.1017155, 
    0.06967424, 0.02932984, 0.04409829, 0.004063622, 7.358856e-05, 
    0.03684857, 0.2222618, 0.1870106, 0.02978122, 0.003144847, 0.009902904, 
    0.01848319, 0.07609348, 0.09815697, 0.1582615, 0.06764767, 0.09921743, 
    0.06931472, 0.04981911, 0.1187525, 0.2206287, 0.1653605,
  0.1045502, 0.05665819, 0.04307478, 0.1027063, 0.1018407, 0.08290793, 
    0.06400606, 0.06281241, 0.008402488, 0, -1.698282e-06, 0.007766665, 
    0.05978532, 0.1158608, 0.08616881, 0.06702265, 0.0976557, 0.1057857, 
    0.02378544, 0.000173729, -0.0006539777, 0.000107538, -0.0002947891, 
    -0.0001283548, 0.0192079, -8.927836e-05, -4.099066e-05, 0.08090495, 
    0.1171694,
  0.03617179, 0.01004141, 0.0001833533, 0, 0, -0.0002248586, 1.144446e-05, 0, 
    0, 0, 0, 0.001608144, 0.01851914, 0.02317938, 0.01971851, 0.01629338, 
    0.006965297, -0.0001771838, 0.0007364343, -4.274271e-05, 0, 
    -1.025012e-05, -7.60388e-06, -9.549662e-06, 0.0001028406, 2.04735e-05, 
    -8.052796e-05, -0.000467106, 0.03667381,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, -1.757755e-08, 0, 0, 0, 0, 0, 0, 0, 0, -3.433902e-07, -1.413205e-06, 
    2.048969e-05, 0.0421872, 0.02300395, 0.1915675, 0.2141865, 0.3430009, 
    0.2986973, 0.1656836, 0.07071453, 0.007606629, 0.1038089, 0.06626572, 
    0.05875028, 0.05475432, 0.08695397, 0.04574247, 0.0004405252,
  0.2151234, 0.269921, 0.2402902, 0.2339899, 0.01865941, 0.07975513, 
    0.2003131, 0.06197573, 0.1142687, 0.1283668, 0.1135591, 0.05095541, 
    0.1245551, 0.09253189, 0.1826625, 0.1997545, 0.2011987, 0.2017158, 
    0.2295042, 0.1614529, 0.09578709, 0.2243773, 0.3126355, 0.2323844, 
    0.3640059, 0.201765, 0.1230927, 0.1950488, 0.2265902,
  0.2133741, 0.1615339, 0.179557, 0.2433007, 0.2063577, 0.1354652, 0.1765482, 
    0.2542022, 0.2871415, 0.2759067, 0.2037904, 0.1937521, 0.1547087, 
    0.1748921, 0.1753088, 0.1129167, 0.1154087, 0.1383426, 0.1736057, 
    0.2244884, 0.2069442, 0.2467138, 0.1812218, 0.2514674, 0.2577903, 
    0.2109231, 0.2042241, 0.2109379, 0.2587253,
  0.182791, 0.2124674, 0.2353382, 0.1868324, 0.1711126, 0.1603284, 0.1339539, 
    0.1713646, 0.1327905, 0.1524341, 0.1474321, 0.1009256, 0.1674764, 
    0.1530993, 0.09775204, 0.1658054, 0.1533482, 0.09376737, 0.08722645, 
    0.1396391, 0.1239926, 0.1338921, 0.123769, 0.09663296, 0.08101726, 
    0.1440053, 0.08756877, 0.136567, 0.2004981,
  0.06470928, 0.05235833, 0.01450639, 0.05534811, 0.05421358, 0.1114989, 
    0.05496056, 0.04716803, 0.01014423, 0.02875659, 0.02632661, 0.05920485, 
    0.05483576, 0.08254404, 0.07445986, 0.1330409, 0.0616545, 0.008206017, 
    0.05017614, 0.0757615, 0.05964212, 0.06261815, 0.02564681, 0.001529576, 
    0.05629481, 0.02952621, 0.04850258, 0.06734082, 0.04178688,
  0.006935549, 1.860938e-08, 0.0414876, 0.000103014, 0.1437472, 0.01967246, 
    0.05805773, 0.02898126, 0.01561675, 0.03457706, 0.04738348, 0.05934603, 
    0.01911087, 0.1893719, 0.06620279, 0.01081383, 0.1629925, 0.0919496, 
    0.144701, 0.06821652, 0.005578088, 6.79607e-07, 4.030727e-09, 
    -1.788463e-05, 0.04920508, 0.2450734, 0.04193869, 0.003267047, 0.06942178,
  0.000633175, 0.01642795, 0.02264026, 0.07053577, 0.1130135, 0.1020948, 
    0.008707301, 0.1105705, 0.002918994, 0.01922834, 0.06144157, 0.02223236, 
    0.08805341, 0.02518836, 0.06327467, 0.06406536, 0.04691305, 0.09627555, 
    0.04598549, 0.05121763, -7.486704e-06, 0.0006931084, 1.169079e-05, 
    0.009381234, 0.09061458, 0.03503653, 0.001255272, 1.702536e-07, 
    4.042361e-07,
  0.0001283433, 0.0385258, 0.2333338, 0.1288012, 0.05373542, 0.0616334, 
    0.08403099, 0.06109494, 0.06787632, 0.07359972, 0.08409997, 0.06326193, 
    0.05191343, 0.03185792, 0.0904512, 0.00978499, 0.02700005, 0.006389771, 
    0.003753245, 0.0004517547, 0, -6.249863e-08, 0.0001767245, 0.1474497, 
    0.2731009, 0.0259013, 0.005586053, 0.0003113997, 1.424804e-07,
  0.002560376, 0.02262955, 0.005947475, 0.004655872, 0.02303814, 0.02246287, 
    0.03460074, 0.03244716, 0.06256592, 0.1605167, 0.006906612, 0.007592311, 
    0.03513877, 0.03058668, 0.0148144, 0.005913734, 0.003881682, 0.005780886, 
    0.01019469, 0.001527008, 0.0006553051, 2.240192e-07, 0.03652523, 
    0.04611384, 0.06196923, 0.03459662, 0.02395828, 0.006197058, 0.0005693203,
  8.409187e-07, 8.016574e-07, 4.276207e-07, 0.002478101, 0.0001166918, 
    0.001987296, 0.001040375, 0.000528933, 0.0007451762, 0.0009988415, 
    0.07693212, 0.05995953, 0.01256492, 0.04803791, 0.04368673, 0.03659724, 
    0.06919581, 0.0574512, 0.02776512, 0.006315291, 0.03376276, 0.01018286, 
    0.001014347, 0.0007102989, 0.04220436, 0.0441745, 0.03897399, 0.00350923, 
    0.0002164764,
  0.005077019, -2.657511e-06, 5.403599e-08, 2.863716e-08, 1.210732e-06, 
    1.974767e-05, -1.761176e-07, 4.75639e-07, 1.544722e-07, 9.18665e-08, 
    0.0005047515, 0.01614383, 0.002243003, 1.969631e-05, 0.01430645, 
    0.02825927, 0.02480115, 1.384713e-05, 0.000451568, 0.04628596, 
    0.001309513, 0.03768465, 0.004570426, 0.005201917, 0.01277079, 
    0.01914332, 0.0002924899, 0.02776267, 0.08263607,
  0.01866523, 0.03328374, 0.02967548, 0.03525678, 0.02085679, 0.05060164, 
    0.03253511, 0.002494431, 0.03355183, 0.2136873, 0.2299155, 0.09905364, 
    0.09374125, 0.08785834, 0.0993458, 0.09660178, 0.1222816, 0.1305111, 
    0.08910751, 0.02318425, 0.05684651, 0.07723653, 0.02194772, 0.02448664, 
    0.04015119, 0.04857081, 0.01288567, 0.0114758, 0.02319414,
  0.07010418, 0.07336932, 0.06510548, 0.07163819, 0.04096011, 0.04945054, 
    0.03940672, 0.1475369, 0.07671367, 0.06214475, 0.07025225, 0.1722638, 
    0.1588477, 0.1341516, 0.1549529, 0.1534905, 0.2310971, 0.2097157, 
    0.2027284, 0.2364503, 0.2157883, 0.1557935, 0.1699874, 0.1713385, 
    0.09133258, 0.1487874, 0.1351167, 0.0807824, 0.09668507,
  0.1835394, 0.2130433, 0.1293799, 0.1591703, 0.1484302, 0.1701474, 
    0.2665154, 0.02907412, 0.008109903, 0.05497883, 0.08384869, 0.1248354, 
    0.2432731, 0.2702112, 0.3191248, 0.1675619, 0.09165587, 0.01647064, 
    0.1517034, 0.1697114, 0.09204849, 0.1348113, 0.2377927, 0.2187736, 
    0.2460766, 0.1996941, 0.164239, 0.2006407, 0.1748963,
  0.2525618, 0.2008497, 0.2542256, 0.2736255, 0.3553852, 0.3112854, 
    0.1977961, 0.1345192, 0.06924415, 0.08376742, 0.04209019, 0.01686824, 
    0.06380075, 0.3056279, 0.1779628, 0.0377952, 0.006615917, 0.03442545, 
    0.0341871, 0.1103299, 0.1640647, 0.1757846, 0.07883538, 0.1142551, 
    0.08258478, 0.1128528, 0.1954261, 0.2909029, 0.2472708,
  0.2023947, 0.1568137, 0.1742151, 0.2889992, 0.2528052, 0.1853195, 
    0.1242408, 0.1314957, 0.05596213, 0.02660305, 0.02202024, 0.04755168, 
    0.105033, 0.1536707, 0.1052306, 0.08731632, 0.1208812, 0.1414386, 
    0.07654387, 0.01151527, -0.0009416354, 0.008213811, 0.0194877, 
    -0.0005298998, 0.0415182, 0.0006705488, 7.772948e-05, 0.1635636, 0.1893115,
  0.06146656, 0.04057127, 0.001789349, -0.0001420017, 0.000748553, 
    -0.0004938098, -0.001161712, 0.006456497, 0.02418028, 0.03647063, 
    0.05557673, 0.05211401, 0.04225772, 0.03860601, 0.05665386, 0.08627033, 
    0.09818044, 0.08182265, 0.04005678, 0.01985974, 0.002107505, 
    -0.0002185291, -7.618683e-05, -0.0002135098, 0.001011437, 0.0001320932, 
    -0.002313695, 0.03133681, 0.05351625,
  1.550498e-05, 5.04163e-06, -5.42172e-06, -1.588507e-05, -2.634842e-05, 
    -3.681177e-05, -4.727512e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -3.513981e-05, -2.467646e-05, -1.421311e-05, -3.749763e-06, 6.713587e-06, 
    1.717694e-05, 2.764029e-05, 2.387566e-05,
  -0.0008809567, -4.098656e-05, 0, 0, 0, -0.0001000005, 0, 0, 0, 
    0.0002197783, 0.0008141721, 0.003080346, 0.0002105071, 0.06658354, 
    0.03107659, 0.2049759, 0.2103967, 0.3579829, 0.3279741, 0.234795, 
    0.1623346, 0.1134246, 0.09237395, 0.06134141, 0.0583454, 0.06480249, 
    0.06619187, 0.06856469, 0.01905273,
  0.2330904, 0.258855, 0.2101846, 0.2398321, 0.09058601, 0.200286, 0.2456265, 
    0.1695676, 0.1725334, 0.200174, 0.1927526, 0.1165899, 0.1389408, 
    0.06017029, 0.1977188, 0.2175662, 0.1926292, 0.1975562, 0.2348717, 
    0.1179613, 0.106265, 0.2804438, 0.3167684, 0.2545166, 0.3127719, 
    0.1956841, 0.1541901, 0.2257916, 0.2151452,
  0.2316305, 0.206824, 0.18925, 0.2331384, 0.2144933, 0.1283263, 0.1791168, 
    0.2792389, 0.3132947, 0.2809776, 0.196686, 0.1899542, 0.1704008, 
    0.1884165, 0.1875777, 0.112727, 0.1114954, 0.1535107, 0.1664345, 
    0.2384158, 0.2424283, 0.2906753, 0.1967384, 0.2588841, 0.278525, 
    0.2135525, 0.1871172, 0.2230344, 0.2684733,
  0.2024372, 0.1993991, 0.2392837, 0.1851152, 0.1789595, 0.1709964, 
    0.1717296, 0.1690351, 0.1357615, 0.1496424, 0.1606176, 0.09387103, 
    0.1794195, 0.1499555, 0.1153895, 0.1467017, 0.1449818, 0.08061592, 
    0.0790531, 0.1303528, 0.09729849, 0.1298666, 0.1337793, 0.09074555, 
    0.07356565, 0.1460093, 0.1044349, 0.1265613, 0.1972371,
  0.06225768, 0.05682913, 0.01402254, 0.06972369, 0.03895816, 0.1012063, 
    0.04416339, 0.04425663, 0.01795764, 0.02732253, 0.03675374, 0.0553365, 
    0.0575172, 0.07003053, 0.07389669, 0.1276037, 0.05499319, 0.009179618, 
    0.05368725, 0.06390098, 0.07440284, 0.05940075, 0.01046091, 0.0005303111, 
    0.05606659, 0.03028966, 0.05946243, 0.07014024, 0.04277462,
  0.01090058, 3.696277e-09, 0.03276106, 2.921536e-05, 0.1334315, 0.02087674, 
    0.03938555, 0.01906092, 0.009489939, 0.02421744, 0.06012405, 0.08294199, 
    0.02113371, 0.1927341, 0.05569358, 0.0105943, 0.172038, 0.08619382, 
    0.1218178, 0.05650947, 0.005257785, 8.381892e-08, 1.613196e-09, 
    -2.313522e-05, 0.04453155, 0.2533888, 0.02377845, 0.002714083, 0.06713414,
  0.002239577, 0.01910656, 0.02679583, 0.09181517, 0.1202267, 0.1113439, 
    0.01490446, 0.1084122, 0.002240346, 0.02755668, 0.06815988, 0.02234868, 
    0.08397461, 0.02655956, 0.07684848, 0.06019475, 0.04276872, 0.106134, 
    0.05231138, 0.04895333, -3.020222e-07, -1.619934e-05, 2.346369e-05, 
    0.01799052, 0.09699926, 0.03441526, 0.001193471, -1.626968e-07, 
    1.96547e-07,
  0.006967001, 0.04909854, 0.2493435, 0.1393499, 0.05438158, 0.06570876, 
    0.09364708, 0.05243514, 0.06992967, 0.08992591, 0.1174877, 0.07060091, 
    0.07585171, 0.03106309, 0.09024833, 0.0101987, 0.0299866, 0.005540117, 
    0.003974755, 0.0004962464, 1.793784e-09, 3.59219e-08, 0.001172374, 
    0.1333788, 0.2945785, 0.02740737, 0.00557055, 0.0001031238, 1.19312e-05,
  0.03402204, 0.03644612, 0.02178689, 0.006650705, 0.02275067, 0.02061715, 
    0.03317006, 0.01711637, 0.05985873, 0.1899079, 0.01079482, 0.00727322, 
    0.02838364, 0.02987057, 0.01538704, 0.005788781, 0.004841625, 0.00290181, 
    0.009928118, 0.001164893, 0.001102127, 3.037537e-05, 0.03091678, 
    0.06345777, 0.07421365, 0.03068773, 0.02803726, 0.004980156, 0.003464169,
  -9.193112e-06, 1.509427e-06, 1.116485e-06, 0.001643263, 0.0008265662, 
    0.001491554, 0.001515674, 0.0004822973, 0.0009689292, 0.000823608, 
    0.08053897, 0.06290609, 0.0221698, 0.05239315, 0.03897629, 0.05375158, 
    0.06154918, 0.06281422, 0.03573759, 0.007962038, 0.03331334, 0.01160593, 
    0.002038323, 0.00146621, 0.05015773, 0.07360136, 0.04888855, 
    0.0002924604, 0.0001246375,
  0.00201756, -1.204852e-07, 4.82784e-09, 3.070625e-08, 1.194803e-06, 
    0.0003854641, -1.369996e-06, -1.58924e-06, 8.802437e-08, -2.457404e-07, 
    0.001797464, 0.01562988, 0.001484319, -2.209537e-05, 0.01450682, 
    0.01277947, 0.0440592, -7.198952e-06, 0.0005090923, 0.04148485, 
    -1.638928e-05, 0.04360747, 0.007905013, 0.003047975, 0.01029827, 
    0.03316272, -3.134719e-05, 0.02426545, 0.09119519,
  0.01842354, 0.02419758, 0.02640774, 0.03434175, 0.0293434, 0.05521961, 
    0.03774732, 0.001935061, 0.0689583, 0.2350329, 0.2243289, 0.1014039, 
    0.09674016, 0.1158394, 0.1023767, 0.09805258, 0.08860989, 0.1029247, 
    0.06961574, 0.01760669, 0.03503868, 0.08231499, 0.007187347, 0.02223634, 
    0.03334815, 0.0401148, 0.01488419, 0.01548143, 0.01690407,
  0.07030086, 0.06381597, 0.05304248, 0.08079134, 0.03716952, 0.03621694, 
    0.09083998, 0.1535672, 0.06322403, 0.06340148, 0.07284656, 0.1757637, 
    0.1552986, 0.1315035, 0.1671126, 0.1607169, 0.2318852, 0.2246422, 
    0.2095345, 0.2389778, 0.2132065, 0.1426758, 0.1615494, 0.1429119, 
    0.08869171, 0.1366916, 0.1224046, 0.08573838, 0.08241225,
  0.1669427, 0.1760382, 0.1125325, 0.1341772, 0.1305025, 0.1648696, 0.293779, 
    0.08742635, 0.05810387, 0.1055237, 0.09577851, 0.1735601, 0.2840653, 
    0.2659447, 0.3091487, 0.161423, 0.08981882, 0.02237419, 0.1753466, 
    0.1910865, 0.1360571, 0.1490024, 0.2339222, 0.2119278, 0.2403641, 
    0.2042627, 0.1777276, 0.2301471, 0.1631032,
  0.2311887, 0.2261318, 0.2550932, 0.2651095, 0.3637983, 0.3409184, 0.27613, 
    0.2856039, 0.1411726, 0.1648251, 0.1119803, 0.0872313, 0.16501, 
    0.2845955, 0.1470643, 0.0373689, 0.01656675, 0.04951459, 0.04686615, 
    0.237756, 0.249896, 0.2157566, 0.1100725, 0.1362398, 0.1052821, 0.201142, 
    0.2464165, 0.3089368, 0.2295725,
  0.2330714, 0.2229419, 0.3530504, 0.4216767, 0.3228486, 0.2295123, 
    0.1726154, 0.1997112, 0.136624, 0.06737393, 0.04203288, 0.08922332, 
    0.1587906, 0.1369413, 0.1051256, 0.08669633, 0.124765, 0.1589314, 
    0.09658256, 0.05539979, 0.01398555, 0.04275924, 0.03163639, 0.01718606, 
    0.07130131, 0.006350168, -0.0002630421, 0.1834183, 0.2265565,
  0.06473465, 0.08338639, 0.04543216, 0.001717469, 0.01601356, 0.07294507, 
    0.09936307, 0.1253701, 0.1814202, 0.1411793, 0.1219229, 0.09532073, 
    0.09674668, 0.1038743, 0.1328978, 0.1316984, 0.1244977, 0.1022711, 
    0.07504911, 0.04454502, 0.04415654, 0.03710376, 0.006110501, 
    -0.0007803729, 0.00503744, 0.0008367153, -0.005090198, 0.05756995, 
    0.05196874,
  0.007066551, 0.006271057, 0.005475563, 0.004680069, 0.003884576, 
    0.003089082, 0.002293588, 0.004540987, 0.004317455, 0.004093922, 
    0.003870389, 0.003646856, 0.003423324, 0.003199791, 0.003021166, 
    0.003615306, 0.004209445, 0.004803584, 0.005397724, 0.005991863, 
    0.006586002, 0.004695019, 0.005119906, 0.005544793, 0.00596968, 
    0.006394568, 0.006819455, 0.007244342, 0.007702946,
  0.006030335, 1.379079e-05, -2.198907e-05, 0, -0.0001791323, 0.001607641, 
    0.001173909, 0.004441101, 0.01242284, 0.006767021, 0.00990775, 
    0.01529142, 0.004617129, 0.08933221, 0.03413218, 0.1982674, 0.2197148, 
    0.3378011, 0.3219862, 0.2284099, 0.2427698, 0.2031515, 0.09994938, 
    0.06210057, 0.05239018, 0.06062094, 0.05786766, 0.06652031, 0.08578569,
  0.2409756, 0.2615567, 0.2087669, 0.250752, 0.2179537, 0.259281, 0.239585, 
    0.3260607, 0.2683822, 0.2752023, 0.2555777, 0.1710247, 0.1329249, 
    0.04346737, 0.2142944, 0.2189561, 0.1944305, 0.2058986, 0.2436725, 
    0.1094605, 0.1688599, 0.328003, 0.3426121, 0.3107318, 0.299437, 
    0.1871473, 0.1871826, 0.2318032, 0.2165076,
  0.2415177, 0.2158444, 0.2185411, 0.2492283, 0.2334824, 0.1382709, 
    0.2043662, 0.3180178, 0.3331425, 0.2809016, 0.2157865, 0.1860996, 
    0.1959936, 0.1819612, 0.2058613, 0.121089, 0.1223148, 0.1623331, 
    0.1645606, 0.2513215, 0.2621283, 0.347808, 0.2332298, 0.2599335, 
    0.2872894, 0.2326926, 0.1971295, 0.2510589, 0.3001504,
  0.2082491, 0.1664949, 0.2141135, 0.1630988, 0.1461385, 0.164026, 0.1956936, 
    0.161452, 0.1355759, 0.1328425, 0.1584522, 0.09807922, 0.1813764, 
    0.1518929, 0.09829438, 0.1407666, 0.1635386, 0.08889227, 0.06436104, 
    0.154434, 0.1020536, 0.123123, 0.1215098, 0.08023504, 0.06943735, 
    0.1446819, 0.1001871, 0.1110601, 0.195735,
  0.05350842, 0.0607372, 0.01632703, 0.06903841, 0.03614532, 0.09630284, 
    0.04558217, 0.04526494, 0.01715105, 0.04055925, 0.0340894, 0.0533751, 
    0.05131203, 0.06951096, 0.07973092, 0.1172966, 0.04934815, 0.02464171, 
    0.0574688, 0.06346287, 0.07163402, 0.05106783, 0.0117223, 0.0002635687, 
    0.05910723, 0.02987462, 0.07064136, 0.07429069, 0.04571652,
  0.0141528, -1.889537e-06, 0.02896562, 8.556719e-05, 0.1246148, 0.02609509, 
    0.02524025, 0.01472833, 0.01025779, 0.01975328, 0.1040733, 0.05270571, 
    0.01267737, 0.1928355, 0.06347831, 0.02856502, 0.1760379, 0.07542091, 
    0.1170085, 0.05777143, 0.007048406, 3.261596e-07, 1.464742e-07, 
    -1.968594e-05, 0.03839678, 0.2834354, 0.01990525, 0.01040359, 0.07222161,
  0.0006613826, 0.04331976, 0.03631523, 0.1131926, 0.1479625, 0.1334438, 
    0.01819058, 0.1152573, 0.003643955, 0.03043048, 0.09416011, 0.03055465, 
    0.08282793, 0.0327592, 0.09301051, 0.05716263, 0.05994811, 0.1448667, 
    0.0703326, 0.05645424, 2.62152e-07, 3.348203e-06, 1.21195e-05, 
    0.02042859, 0.1216426, 0.03416554, 0.001763726, 2.057584e-07, 6.767402e-07,
  0.004300287, 0.05576575, 0.2715443, 0.1716606, 0.06576155, 0.09307633, 
    0.1029738, 0.06331773, 0.08617754, 0.1296894, 0.1764542, 0.08676715, 
    0.127523, 0.04243237, 0.09118941, 0.01597809, 0.03626514, 0.006444725, 
    0.00484511, 0.001108381, 1.998362e-07, 2.762438e-06, 0.001261241, 
    0.1382537, 0.3301024, 0.02962423, 0.008970765, 0.0001383168, 0.0007163772,
  0.145428, 0.04505847, 0.03569039, 0.01241914, 0.02449792, 0.02054111, 
    0.03629879, 0.02001554, 0.09521551, 0.2406293, 0.01727922, 0.01428779, 
    0.03731068, 0.03183689, 0.01248188, 0.004773976, 0.01112209, 0.004478643, 
    0.008925694, 0.004250664, 0.003243896, 0.01303323, 0.04351281, 
    0.09216914, 0.1078558, 0.03649012, 0.03150556, 0.004804616, 0.08434843,
  -1.735066e-06, 1.511761e-06, 0.0001607891, 0.0185855, 0.002232106, 
    0.001717252, 0.002797651, 0.0009951205, 0.001643161, 0.001549578, 
    0.1092522, 0.07373771, 0.04109251, 0.05566581, 0.04637236, 0.05461608, 
    0.06294032, 0.06397657, 0.03284747, 0.009747488, 0.03474563, 0.008316856, 
    0.005128929, 0.002381099, 0.06338646, 0.09378466, 0.05382237, 
    0.001513129, 0.001435618,
  -5.394028e-06, 2.043443e-06, -3.45459e-08, -7.300494e-09, 8.769219e-05, 
    0.0008362463, -1.817933e-05, -9.826116e-07, 6.744892e-08, -3.123959e-06, 
    0.007124373, 0.02474883, 0.0001359381, 0.001387291, 0.02172874, 
    0.0003726334, 0.05327757, 6.458661e-05, 0.001331678, 0.03899502, 
    0.00380082, 0.05748104, 0.01862748, 0.005787199, 0.009059534, 0.04877635, 
    5.554351e-05, 0.06900089, 0.07515115,
  0.01833027, 0.02320632, 0.02191909, 0.02813601, 0.03333839, 0.05830652, 
    0.03593637, 0.0003335986, 0.1060869, 0.2531713, 0.2305728, 0.1168877, 
    0.07350604, 0.1241267, 0.08928699, 0.08565307, 0.06418031, 0.09377484, 
    0.05511733, 0.01739231, 0.02324225, 0.06941112, 0.009252778, 0.02522653, 
    0.02781522, 0.03804904, 0.01277816, 0.01119532, 0.01856496,
  0.06423624, 0.06320272, 0.04754004, 0.08570433, 0.03679864, 0.03738995, 
    0.1530155, 0.1284682, 0.04497439, 0.05584236, 0.07648219, 0.1575301, 
    0.1634464, 0.1488818, 0.1642765, 0.1686426, 0.2274259, 0.2213212, 
    0.2012015, 0.2423639, 0.2077714, 0.1271212, 0.15148, 0.1398688, 
    0.07691734, 0.1254804, 0.1084354, 0.0695351, 0.08670153,
  0.1615392, 0.1508233, 0.09345441, 0.1588061, 0.1360848, 0.1582735, 
    0.2397733, 0.1632351, 0.1231679, 0.1436033, 0.1034471, 0.1539826, 
    0.2709096, 0.2762064, 0.3046829, 0.1540205, 0.07422476, 0.0266797, 
    0.1855647, 0.2382549, 0.1483076, 0.1524111, 0.224906, 0.2208826, 
    0.2725289, 0.2195374, 0.1988995, 0.2130894, 0.1759428,
  0.2130094, 0.2266997, 0.2427702, 0.2573545, 0.3894659, 0.3549979, 
    0.2852378, 0.3163751, 0.3007298, 0.2386519, 0.1822698, 0.2019399, 
    0.2584342, 0.2611038, 0.1171097, 0.03527655, 0.01666771, 0.06446555, 
    0.05889357, 0.3234558, 0.2607878, 0.2477902, 0.1476626, 0.1702628, 
    0.1363225, 0.2793804, 0.236009, 0.3173556, 0.1932078,
  0.220433, 0.1890529, 0.350949, 0.4477133, 0.3166736, 0.215138, 0.1880649, 
    0.2636153, 0.200601, 0.1000028, 0.07673252, 0.1038749, 0.1648343, 
    0.1489048, 0.1401571, 0.1338654, 0.1763092, 0.1563416, 0.08859845, 
    0.1331972, 0.07043061, 0.07589695, 0.1144259, 0.03830785, 0.1011515, 
    0.01230906, 0.004507822, 0.1911747, 0.2265891,
  0.07447608, 0.1574955, 0.1930109, 0.1729299, 0.1977605, 0.1823275, 
    0.167058, 0.2095615, 0.2839698, 0.2368723, 0.1940706, 0.1724268, 
    0.1533466, 0.1718653, 0.2040658, 0.1860767, 0.1744693, 0.140069, 
    0.1077541, 0.05605987, 0.06941714, 0.1021301, 0.02269355, -0.004228644, 
    0.03901906, 0.007266524, 0.02573958, 0.06001282, 0.05021511,
  0.03892121, 0.03680561, 0.03469002, 0.03257442, 0.03045882, 0.02834322, 
    0.02622762, 0.03133919, 0.03141388, 0.03148855, 0.03156323, 0.03163791, 
    0.03171259, 0.03178727, 0.02689776, 0.03074053, 0.0345833, 0.03842607, 
    0.04226884, 0.04611161, 0.04995437, 0.05561877, 0.05381691, 0.05201507, 
    0.05021321, 0.04841137, 0.04660951, 0.04480767, 0.04061369,
  0.08309711, 0.01622687, 0.0003384278, 0.0009594586, -0.0006127956, 
    0.01294565, 0.02037459, 0.02995466, 0.01977169, 0.01658265, 0.02540159, 
    0.02285997, 0.03698068, 0.1042653, 0.04720467, 0.1703819, 0.239571, 
    0.3323617, 0.2762944, 0.2021932, 0.305544, 0.306895, 0.110004, 
    0.06454282, 0.04818834, 0.05755948, 0.04902716, 0.0620435, 0.1008719,
  0.2539111, 0.2565067, 0.2055427, 0.2429099, 0.2711482, 0.2863658, 
    0.2921316, 0.4204608, 0.3287989, 0.3133315, 0.2589213, 0.179548, 
    0.1390358, 0.05401222, 0.2391227, 0.2153122, 0.1952115, 0.2205218, 
    0.2780905, 0.1329079, 0.1929154, 0.2861262, 0.3035117, 0.3822623, 
    0.2956379, 0.1953825, 0.2121772, 0.2212899, 0.2624865,
  0.2671206, 0.2181845, 0.2062354, 0.263316, 0.2460653, 0.1565593, 0.2442361, 
    0.3009265, 0.3622539, 0.3157166, 0.1830407, 0.2177485, 0.2055304, 
    0.1719346, 0.198082, 0.104237, 0.1288537, 0.1571228, 0.2000865, 
    0.2736588, 0.3514607, 0.3227558, 0.2542116, 0.2501383, 0.2885199, 
    0.2440249, 0.2083781, 0.2836966, 0.3580058,
  0.199962, 0.1594033, 0.2385829, 0.156953, 0.1569054, 0.2056871, 0.166568, 
    0.182294, 0.1312874, 0.1304912, 0.1226768, 0.08058897, 0.1871113, 
    0.1569137, 0.1162415, 0.1426999, 0.1459576, 0.0837665, 0.05996143, 
    0.1517174, 0.1024059, 0.1132341, 0.1358247, 0.07772772, 0.07256842, 
    0.1297609, 0.1080019, 0.1290753, 0.1927639,
  0.05397188, 0.06304168, 0.01703256, 0.06691098, 0.0406649, 0.0948572, 
    0.05104201, 0.04489364, 0.02596985, 0.0492349, 0.03127578, 0.05609665, 
    0.0649497, 0.07232901, 0.09342174, 0.12393, 0.05124633, 0.02832753, 
    0.06851073, 0.0759029, 0.07396333, 0.04862894, 0.009899968, 0.001144365, 
    0.05063557, 0.03160544, 0.08704147, 0.08798338, 0.05456693,
  0.03221124, 1.824721e-06, 0.03095536, 0.0002457584, 0.1292012, 0.03825346, 
    0.01936892, 0.008440212, 0.01879443, 0.02053159, 0.1349901, 0.04131742, 
    0.02116911, 0.1974895, 0.07233969, 0.03414831, 0.1754065, 0.07490863, 
    0.1144834, 0.07162803, 0.01745917, 1.217445e-07, 1.904202e-07, 
    9.680261e-06, 0.03786885, 0.3110201, 0.01978093, 0.01627111, 0.07939192,
  0.0003869783, 0.09327406, 0.06038107, 0.1238471, 0.1565004, 0.147257, 
    0.02401587, 0.1193873, 0.002342776, 0.03344306, 0.1261715, 0.03428758, 
    0.0959933, 0.03093255, 0.09585709, 0.06169593, 0.0843311, 0.1712923, 
    0.08967622, 0.0700566, 1.80877e-05, 2.987045e-06, 9.045323e-06, 
    0.01333613, 0.1707414, 0.03629532, 0.004510465, 5.089458e-07, 1.053506e-06,
  0.001783663, 0.05834795, 0.3120196, 0.2219888, 0.07174867, 0.1102122, 
    0.1075159, 0.07013574, 0.1098222, 0.1467361, 0.2067869, 0.08689596, 
    0.1557147, 0.05795979, 0.09940373, 0.02053619, 0.04563355, 0.006470061, 
    0.009772812, 0.002538346, 3.478895e-06, 2.007228e-06, 0.001293295, 
    0.1503832, 0.340511, 0.04029893, 0.01171941, 0.0001840269, 4.603229e-05,
  0.177397, 0.04675724, 0.0287949, 0.02580213, 0.02140491, 0.02547562, 
    0.04730271, 0.02292319, 0.1247723, 0.2853375, 0.01940503, 0.01965147, 
    0.0426356, 0.04680109, 0.01307767, 0.005305147, 0.00783296, 0.007030458, 
    0.03606378, 0.01553662, 0.009552024, 0.03723253, 0.07248177, 0.1374288, 
    0.1477618, 0.03915949, 0.0271635, 0.003654509, 0.08835953,
  9.054509e-05, 5.06778e-06, 0.008048885, 0.07478168, 0.00477751, 
    0.002049279, 0.005103379, 0.002692056, 0.001641712, 0.005176523, 
    0.1284935, 0.09167656, 0.05304248, 0.05057956, 0.05093032, 0.05335436, 
    0.05972745, 0.07164791, 0.02517341, 0.01188417, 0.03773174, 0.007123976, 
    0.01071058, 0.004568283, 0.08068353, 0.06883129, 0.03014598, 0.008781446, 
    0.01643278,
  -5.455089e-06, 1.773056e-06, 3.121428e-07, -5.126053e-09, 0.001918479, 
    0.0002476156, -2.014909e-05, 1.604778e-06, 2.935992e-07, -7.883832e-06, 
    0.02468524, 0.0306145, 0.0001123628, 0.03641399, 0.02749651, 
    0.0006403713, 0.05837305, 7.431974e-05, 0.002384116, 0.03336682, 
    0.001215716, 0.08006456, 0.02042327, 0.008451876, 0.01205036, 0.04938828, 
    0.0001468271, 0.04311134, 0.02947906,
  0.01748583, 0.03052456, 0.02185633, 0.03079426, 0.03643799, 0.0580494, 
    0.04093909, 0.002574314, 0.1309258, 0.247436, 0.2135759, 0.1115828, 
    0.07648183, 0.1275604, 0.09521345, 0.08496955, 0.0548934, 0.08784443, 
    0.0524834, 0.01865749, 0.01664138, 0.05759046, 0.01762681, 0.03215659, 
    0.02925232, 0.04227617, 0.01278382, 0.01123465, 0.01946747,
  0.0643173, 0.05966447, 0.04230436, 0.08457296, 0.02850156, 0.03048403, 
    0.1825681, 0.07615145, 0.03646072, 0.04919112, 0.07298625, 0.1319515, 
    0.1576448, 0.188653, 0.1774489, 0.1787164, 0.2140219, 0.2269838, 
    0.1990368, 0.2441706, 0.2072953, 0.1269453, 0.1381522, 0.1368127, 
    0.07646752, 0.1089775, 0.1069301, 0.07486442, 0.08834424,
  0.1642644, 0.1429096, 0.1007568, 0.1373135, 0.1382708, 0.1662315, 
    0.2435717, 0.2115089, 0.1569725, 0.1389987, 0.09807333, 0.1486977, 
    0.2568924, 0.2920589, 0.3048832, 0.1264431, 0.05280643, 0.02759965, 
    0.1884891, 0.2972367, 0.1406799, 0.1415848, 0.2353178, 0.2171874, 
    0.2849624, 0.2329714, 0.2023427, 0.2301524, 0.2061309,
  0.2020533, 0.2243878, 0.2476468, 0.2578312, 0.3754533, 0.3435339, 
    0.2958936, 0.3414199, 0.3346535, 0.2791068, 0.2674868, 0.2018889, 
    0.268941, 0.2672496, 0.08092247, 0.03175069, 0.01728739, 0.0714001, 
    0.0991766, 0.3453771, 0.2468221, 0.247018, 0.1541059, 0.1732788, 
    0.1576745, 0.3552731, 0.2545966, 0.3313204, 0.2039506,
  0.2240983, 0.2158493, 0.3721688, 0.4282867, 0.3182288, 0.2104017, 
    0.2160203, 0.3347583, 0.3235722, 0.156593, 0.09028991, 0.1198653, 
    0.2073769, 0.1551755, 0.1473655, 0.1314836, 0.1693915, 0.1683557, 
    0.09250484, 0.1570017, 0.08640673, 0.07984154, 0.09106693, 0.05964711, 
    0.1455868, 0.0470209, 0.01403972, 0.1740142, 0.2424517,
  0.0919345, 0.2243014, 0.1891164, 0.182864, 0.2705728, 0.2673555, 0.2123418, 
    0.2186511, 0.3040703, 0.2824284, 0.2162626, 0.1943698, 0.1735059, 
    0.1805044, 0.2179065, 0.1990649, 0.1846307, 0.1695261, 0.1370003, 
    0.1274326, 0.1188894, 0.1445906, 0.1075549, 0.02083392, 0.04761821, 
    0.01125199, 0.04662936, 0.0575671, 0.05918706,
  0.07216924, 0.06890453, 0.06563983, 0.06237512, 0.05911042, 0.05584572, 
    0.05258102, 0.05666578, 0.06209864, 0.06753151, 0.07296437, 0.07839723, 
    0.0838301, 0.08926295, 0.06883302, 0.07276398, 0.07669494, 0.08062589, 
    0.08455685, 0.0884878, 0.09241876, 0.1182099, 0.1121108, 0.1060117, 
    0.09991254, 0.09381343, 0.08771431, 0.08161519, 0.074781,
  0.08641893, 0.06942788, 0.03748229, 0.01243661, 0.0226815, 0.03885707, 
    0.043913, 0.03969666, 0.02867214, 0.01482286, 0.02018958, 0.06615493, 
    0.1093268, 0.1461773, 0.03837803, 0.2421456, 0.232553, 0.3091834, 
    0.2223605, 0.1706408, 0.27057, 0.3125667, 0.1249316, 0.06168814, 
    0.07569593, 0.05235736, 0.05996509, 0.06812053, 0.09307039,
  0.2562633, 0.2560354, 0.2270401, 0.2285601, 0.2637713, 0.2742232, 
    0.3807884, 0.4441608, 0.3649922, 0.3317313, 0.2436361, 0.1752464, 
    0.1116607, 0.03656142, 0.2550505, 0.2411797, 0.2399082, 0.2557776, 
    0.3065964, 0.2231492, 0.3236714, 0.3395096, 0.2412493, 0.3018087, 
    0.3051243, 0.1851066, 0.2309477, 0.2741832, 0.2808439,
  0.2886003, 0.2375903, 0.2590035, 0.2664185, 0.2731002, 0.1829094, 
    0.2800141, 0.4137725, 0.3987319, 0.3478822, 0.1719239, 0.2300725, 
    0.2044207, 0.1934162, 0.1806833, 0.09728853, 0.1226197, 0.1777077, 
    0.2182977, 0.3316035, 0.3624534, 0.35972, 0.2837726, 0.2962286, 
    0.2896138, 0.2491499, 0.2428901, 0.2970277, 0.3601644,
  0.209914, 0.1742446, 0.2238258, 0.1624019, 0.1655442, 0.1686957, 0.1977169, 
    0.2154858, 0.1337877, 0.1383319, 0.1335285, 0.1009677, 0.1934068, 
    0.157525, 0.1060346, 0.1633665, 0.150529, 0.1042631, 0.08513848, 
    0.1573669, 0.1199463, 0.1181791, 0.1442174, 0.08322492, 0.086425, 
    0.1245103, 0.1145684, 0.1257468, 0.2099195,
  0.05323774, 0.06850329, 0.01105007, 0.07322276, 0.0522629, 0.1029533, 
    0.05295774, 0.0331411, 0.0288519, 0.05644913, 0.04077767, 0.06622549, 
    0.05742837, 0.08170112, 0.1161323, 0.1282709, 0.07602853, 0.039665, 
    0.07471289, 0.07897229, 0.08208961, 0.05281003, 0.01694238, 0.002304661, 
    0.04165861, 0.03978039, 0.104777, 0.09223521, 0.06090728,
  0.02952308, -3.272588e-06, 0.04385467, 0.0004161618, 0.1282307, 0.05877512, 
    0.01753005, 0.006901952, 0.0257421, 0.01439811, 0.1265168, 0.01786221, 
    0.02035875, 0.2032498, 0.06622342, 0.04761015, 0.1863475, 0.08398806, 
    0.1142545, 0.08818665, 0.02853745, 2.68846e-07, 3.064438e-07, 
    0.0001331465, 0.05273814, 0.3197725, 0.02535479, 0.02198713, 0.08284692,
  0.0002762091, 0.112986, 0.0777955, 0.1209322, 0.1249647, 0.1366127, 
    0.03399983, 0.1150334, 0.002621801, 0.02535872, 0.1089381, 0.03075195, 
    0.07428679, 0.03160274, 0.07868392, 0.05548101, 0.06613377, 0.1499425, 
    0.09056886, 0.07472869, 0.001726064, 1.445556e-06, 5.354911e-06, 
    0.002657317, 0.1784032, 0.04894353, 0.008466423, -3.418487e-06, 
    8.341335e-07,
  6.74418e-06, 0.04010116, 0.3391314, 0.2262206, 0.05042658, 0.09592571, 
    0.0936471, 0.06483942, 0.09518267, 0.1044459, 0.1764337, 0.06655849, 
    0.1246097, 0.04784271, 0.08735561, 0.0203873, 0.03332953, 0.006850368, 
    0.00947908, 0.003600334, 8.142059e-05, 7.451338e-07, 0.0004004244, 
    0.1724539, 0.3184941, 0.06342109, 0.0138622, 0.0001232201, 7.9942e-07,
  0.0931145, 0.03680315, 0.01282003, 0.03083546, 0.02113174, 0.02098567, 
    0.03138392, 0.01614685, 0.1178929, 0.3238049, 0.02385172, 0.0141573, 
    0.0239098, 0.04526008, 0.01169644, 0.007775143, 0.009401816, 0.02079856, 
    0.06617088, 0.01766455, 0.01603852, 0.03067266, 0.1006324, 0.1471142, 
    0.1759707, 0.03655885, 0.02833821, 0.004704195, 0.02641867,
  -0.0003419905, 5.864604e-06, 0.001508596, 0.12311, 0.004937075, 
    0.005164491, 0.006440418, 0.001849523, 0.003734761, 0.00302474, 
    0.1418082, 0.08172385, 0.04611487, 0.04327608, 0.05061589, 0.05808825, 
    0.05670912, 0.06788901, 0.0223468, 0.01715071, 0.04359753, 0.009964892, 
    0.009420138, 0.005887248, 0.06867177, 0.07278375, 0.01702308, 
    0.009288925, 0.0226834,
  1.594853e-06, 7.7291e-07, 8.708006e-07, 1.253496e-08, 0.00109385, 
    1.568987e-05, -2.886228e-06, 8.521991e-05, 2.758369e-07, -0.0002620699, 
    0.05778705, 0.03600378, 0.007189985, 0.04152862, 0.03145704, 0.001849198, 
    0.07992769, 2.731061e-05, 0.005195732, 0.02087064, 2.609463e-05, 
    0.09909576, 0.02276036, 0.01147693, 0.01954412, 0.06417655, 0.001619908, 
    0.02354542, 0.002942595,
  0.017699, 0.03437922, 0.01355497, 0.04040872, 0.04049612, 0.05559917, 
    0.04098348, 0.005580621, 0.1618315, 0.2267557, 0.2136556, 0.1057595, 
    0.0792492, 0.1229478, 0.09058608, 0.07809916, 0.05555137, 0.08957078, 
    0.05932103, 0.02683577, 0.02441332, 0.05571771, 0.02756139, 0.03776736, 
    0.03429528, 0.04185014, 0.0153633, 0.02291914, 0.01664832,
  0.04560965, 0.0509161, 0.03104996, 0.08630735, 0.011875, 0.02628792, 
    0.2029266, 0.03537759, 0.02689157, 0.05075373, 0.07352522, 0.1162757, 
    0.1488507, 0.1859296, 0.1906969, 0.1772992, 0.2069615, 0.2336946, 
    0.2100454, 0.2407291, 0.2103079, 0.09731935, 0.1187665, 0.1292838, 
    0.08600824, 0.1043677, 0.1074255, 0.07815042, 0.1023501,
  0.1605487, 0.1323955, 0.09453202, 0.1169548, 0.1253691, 0.1574334, 
    0.2203653, 0.2470537, 0.1498033, 0.138111, 0.1006887, 0.1348122, 
    0.2460132, 0.274495, 0.3437484, 0.100538, 0.04612284, 0.05850397, 
    0.2109457, 0.2899722, 0.1368405, 0.1477843, 0.2336038, 0.2148277, 
    0.2842183, 0.219161, 0.2135074, 0.2444517, 0.2056265,
  0.1967217, 0.2324076, 0.2645444, 0.3001319, 0.4213036, 0.34366, 0.3133828, 
    0.3908504, 0.3423775, 0.2593566, 0.3094043, 0.1982571, 0.2810596, 
    0.2869343, 0.05448025, 0.01578556, 0.02550196, 0.07012264, 0.131403, 
    0.3121327, 0.2560636, 0.2450834, 0.1530696, 0.156305, 0.1485758, 
    0.3532205, 0.2654705, 0.317764, 0.2191928,
  0.2345228, 0.2248889, 0.3828215, 0.4630688, 0.318345, 0.2288818, 0.2723378, 
    0.3496823, 0.3604819, 0.192202, 0.1027402, 0.1357121, 0.2138865, 
    0.1595905, 0.1455331, 0.1486783, 0.1732991, 0.1724068, 0.09019111, 
    0.1840431, 0.1144447, 0.08175828, 0.087869, 0.07543357, 0.1506365, 
    0.08992627, 0.06444033, 0.156378, 0.2356718,
  0.1438709, 0.2315473, 0.1637155, 0.1954315, 0.2731323, 0.2693679, 
    0.1999497, 0.2154295, 0.3092337, 0.2943178, 0.2259381, 0.1964825, 
    0.1736461, 0.2059451, 0.2401292, 0.2132529, 0.1813311, 0.2281439, 
    0.1995214, 0.1727503, 0.1768639, 0.198553, 0.1513969, 0.08506081, 
    0.06277253, 0.02558561, 0.05667687, 0.06144614, 0.08214775,
  0.09311233, 0.0903368, 0.08756128, 0.08478575, 0.08201023, 0.07923471, 
    0.07645918, 0.07055508, 0.07997033, 0.08938558, 0.09880082, 0.1082161, 
    0.1176313, 0.1270466, 0.1319727, 0.1313426, 0.1307126, 0.1300826, 
    0.1294526, 0.1288226, 0.1281925, 0.134755, 0.1287453, 0.1227356, 
    0.1167259, 0.1107162, 0.1047065, 0.09869678, 0.09533274,
  0.07210723, 0.06494962, 0.07636929, 0.04310196, 0.05496977, 0.1006907, 
    0.1112356, 0.07498006, 0.04154182, 0.01413643, 0.02015921, 0.1216828, 
    0.1173743, 0.1834569, 0.1372409, 0.3688265, 0.3062438, 0.2937831, 
    0.2330623, 0.2121571, 0.2720922, 0.3545289, 0.1124615, 0.06847457, 
    0.0733158, 0.08481252, 0.08909392, 0.07895438, 0.0881862,
  0.287734, 0.3210369, 0.2489739, 0.2716426, 0.2785625, 0.2840416, 0.4417733, 
    0.4502183, 0.3919989, 0.3493181, 0.2349702, 0.1648313, 0.1225284, 
    0.06020664, 0.2880555, 0.2881306, 0.2433339, 0.2622108, 0.380601, 
    0.1902235, 0.3809923, 0.3751862, 0.2918004, 0.3326467, 0.2845269, 
    0.1910034, 0.2554381, 0.3725094, 0.3948321,
  0.2979883, 0.2926904, 0.3088429, 0.2550077, 0.2913967, 0.2306682, 0.330777, 
    0.4162957, 0.4116443, 0.2875131, 0.1542294, 0.2356121, 0.1981818, 
    0.1676833, 0.1817432, 0.1378683, 0.1351151, 0.2016787, 0.2504034, 
    0.3699323, 0.3523379, 0.3001892, 0.27899, 0.2632997, 0.2660773, 
    0.2791753, 0.2845864, 0.3401302, 0.4038595,
  0.2091218, 0.1867015, 0.2232761, 0.1750807, 0.1718245, 0.1950498, 
    0.1989416, 0.213179, 0.1379775, 0.1538549, 0.1360892, 0.1125284, 
    0.2071711, 0.1648484, 0.1357728, 0.1763795, 0.1398678, 0.1016101, 
    0.08230362, 0.1743855, 0.140662, 0.1364577, 0.1587362, 0.09824156, 
    0.08431006, 0.1132231, 0.1143902, 0.103057, 0.1976383,
  0.05611994, 0.08110948, 0.006931644, 0.0730451, 0.06078425, 0.1058529, 
    0.06285886, 0.03605887, 0.04002608, 0.04928995, 0.04666444, 0.0736022, 
    0.06417905, 0.08576974, 0.1325697, 0.1339093, 0.10032, 0.05271105, 
    0.07384291, 0.08097075, 0.09448609, 0.06130591, 0.02587178, 0.00389649, 
    0.03580681, 0.03292689, 0.1138386, 0.0871396, 0.06288464,
  0.02748471, -1.97259e-05, 0.06673406, 0.001591883, 0.09196179, 0.07630891, 
    0.01832859, 0.006806951, 0.02690069, 0.02119518, 0.06713772, 0.01058384, 
    0.02729097, 0.1654916, 0.04244966, 0.04844483, 0.1960384, 0.07961194, 
    0.1175054, 0.09011207, 0.02875223, 3.986879e-06, 9.617198e-08, 
    0.0001809251, 0.04449288, 0.2445395, 0.02947484, 0.02562298, 0.08111033,
  0.001143145, 0.1072473, 0.08008242, 0.1237177, 0.1120765, 0.1197332, 
    0.03808277, 0.1043556, 0.001387799, 0.0231629, 0.09157617, 0.02098397, 
    0.04974095, 0.02977443, 0.06344865, 0.04471797, 0.04852565, 0.1113954, 
    0.08000948, 0.06694826, 0.01487517, 5.982652e-07, 3.919548e-06, 
    0.0004988473, 0.1554065, 0.05775949, 0.01433184, -1.164164e-05, 
    5.658871e-07,
  2.3566e-06, 0.01131863, 0.3585346, 0.13438, 0.03916788, 0.07756995, 
    0.07314623, 0.06099144, 0.07759922, 0.07366531, 0.147863, 0.04978237, 
    0.1084254, 0.0449481, 0.07358225, 0.02227682, 0.03198956, 0.0102292, 
    0.02054138, 0.007219659, 0.0004316939, 2.418451e-06, 0.0002597967, 
    0.1122847, 0.2106505, 0.06730842, 0.01763372, 0.000274553, 2.721424e-07,
  0.0144488, 0.02177464, 0.002962864, 0.04707643, 0.02266708, 0.01762741, 
    0.02571156, 0.0113295, 0.1000156, 0.2989001, 0.02182825, 0.01221434, 
    0.01308112, 0.0359412, 0.0138488, 0.01481924, 0.009664777, 0.01823682, 
    0.05748672, 0.01415257, 0.0281004, 0.02916269, 0.1321929, 0.1220792, 
    0.1522877, 0.03890206, 0.03285846, 0.009529753, 0.002054847,
  -0.0001740712, 4.108289e-06, 5.71556e-05, 0.194892, 0.005947795, 
    0.01711746, 0.00759086, 0.002231607, 0.00562253, 0.006789779, 0.1351365, 
    0.07391221, 0.03256254, 0.03161092, 0.04644777, 0.06010342, 0.04714703, 
    0.05667438, 0.01904852, 0.02556102, 0.03892078, 0.01050949, 0.01214379, 
    0.01057328, 0.04754313, 0.03468651, 0.004122983, 0.002385938, 0.004792666,
  2.415208e-06, 6.659269e-07, 2.984256e-07, 1.761673e-08, 0.01283476, 
    1.870227e-05, -1.624543e-06, 0.0007080014, 2.73755e-07, 6.863997e-05, 
    0.1561783, 0.04092329, 0.01554184, 0.03173289, 0.02549023, 0.003281774, 
    0.1067186, -1.752584e-05, 0.003353791, 0.009431213, 3.440566e-07, 
    0.1081461, 0.02262557, 0.01972091, 0.02629762, 0.08630881, 0.00547552, 
    0.007636759, 0.001773219,
  0.006821194, 0.04078201, 0.01454325, 0.04619715, 0.04326942, 0.05080351, 
    0.04104741, 0.00998083, 0.1741639, 0.1904455, 0.1859235, 0.1024048, 
    0.09741914, 0.1301291, 0.09576182, 0.08901484, 0.06236574, 0.09766663, 
    0.06911053, 0.03437265, 0.02773344, 0.06511854, 0.02542693, 0.03529932, 
    0.04012432, 0.04217301, 0.02249452, 0.01174417, 0.005919391,
  0.03694569, 0.05026797, 0.03017466, 0.08944388, 0.008080369, 0.03290368, 
    0.2201966, 0.02429182, 0.01566995, 0.05242636, 0.07339267, 0.1124459, 
    0.1521984, 0.1947022, 0.1726912, 0.1744064, 0.207242, 0.2308268, 
    0.2363333, 0.2456343, 0.2032211, 0.0755839, 0.1056857, 0.1400855, 
    0.1110817, 0.1084872, 0.1148359, 0.08579229, 0.1303069,
  0.1619241, 0.1261747, 0.09574487, 0.1153545, 0.1153857, 0.1316865, 
    0.2334153, 0.2747341, 0.1401534, 0.1166723, 0.09211912, 0.1297517, 
    0.2450887, 0.2967534, 0.3714899, 0.07536232, 0.03405765, 0.0853079, 
    0.2487104, 0.3010279, 0.1378293, 0.1490213, 0.2223071, 0.1937179, 
    0.2921278, 0.2195388, 0.2312306, 0.2597094, 0.2146129,
  0.1934715, 0.2519895, 0.3130422, 0.3203762, 0.4088286, 0.3761995, 
    0.3224066, 0.4061766, 0.3084012, 0.2539393, 0.3148895, 0.1819102, 
    0.2847617, 0.32204, 0.06928626, 0.01053029, 0.02746737, 0.06065656, 
    0.1556485, 0.263331, 0.2780953, 0.2317698, 0.1542755, 0.1593673, 
    0.137273, 0.3456958, 0.2759214, 0.3244097, 0.2229684,
  0.244602, 0.2146822, 0.4239365, 0.4769622, 0.3443008, 0.2429069, 0.2821089, 
    0.3698645, 0.3654446, 0.2053843, 0.109314, 0.1524202, 0.2140124, 
    0.1916029, 0.1423519, 0.1707564, 0.1878712, 0.1889794, 0.1021674, 
    0.1895662, 0.1388789, 0.09005805, 0.08715633, 0.1040287, 0.1375254, 
    0.2053523, 0.1606645, 0.161248, 0.251476,
  0.161012, 0.2479252, 0.183564, 0.1846506, 0.2710682, 0.2829908, 0.1923963, 
    0.2140244, 0.3030511, 0.2969845, 0.2480939, 0.1972884, 0.1824362, 
    0.2378329, 0.2756136, 0.2606023, 0.2312381, 0.2879857, 0.2459789, 
    0.2500345, 0.2037121, 0.2379161, 0.1606607, 0.1085368, 0.07446876, 
    0.02565337, 0.06149334, 0.05500645, 0.1052841,
  0.08248186, 0.08157716, 0.08067245, 0.07976774, 0.07886303, 0.07795832, 
    0.07705361, 0.07314065, 0.08050318, 0.08786572, 0.09522825, 0.1025908, 
    0.1099533, 0.1173159, 0.1227453, 0.1209847, 0.1192241, 0.1174635, 
    0.1157029, 0.1139423, 0.1121817, 0.1180792, 0.113382, 0.1086847, 
    0.1039875, 0.09929029, 0.09459306, 0.08989584, 0.08320563,
  0.0509961, 0.0549494, 0.07764219, 0.1011833, 0.1414639, 0.250066, 
    0.2163839, 0.1290129, 0.03882112, 0.01784473, 0.05819377, 0.1316691, 
    0.1255094, 0.1879243, 0.1186098, 0.3406695, 0.2345326, 0.2317689, 
    0.2173548, 0.2083335, 0.3109809, 0.3509712, 0.105737, 0.09328874, 
    0.09510886, 0.07820942, 0.06606144, 0.1074962, 0.0799801,
  0.3343349, 0.3331505, 0.2655874, 0.2995448, 0.3349161, 0.3352073, 
    0.4431993, 0.478391, 0.3940301, 0.349577, 0.2694143, 0.1616077, 
    0.1018224, 0.07191555, 0.3537593, 0.4442889, 0.3272014, 0.2908946, 
    0.4211237, 0.1969431, 0.2664594, 0.3200169, 0.2145871, 0.3132451, 
    0.2711383, 0.2035929, 0.3114621, 0.4467264, 0.4789094,
  0.297284, 0.3714401, 0.3368085, 0.3120336, 0.303704, 0.2585203, 0.3828246, 
    0.4914523, 0.4592167, 0.3074294, 0.2317483, 0.2494841, 0.1995706, 
    0.1681374, 0.2051379, 0.1496578, 0.155481, 0.2333023, 0.3212003, 
    0.3638441, 0.3196115, 0.2606084, 0.2432338, 0.2637378, 0.2773672, 
    0.3122094, 0.2826086, 0.261624, 0.322875,
  0.2130862, 0.1897313, 0.2397034, 0.1885832, 0.1787903, 0.2014699, 
    0.2286572, 0.2158393, 0.1531865, 0.168512, 0.15437, 0.1041631, 0.191557, 
    0.1847547, 0.1632861, 0.1910277, 0.1456546, 0.1192735, 0.1125113, 
    0.1772082, 0.1600272, 0.1600155, 0.1590766, 0.1188463, 0.09306863, 
    0.127555, 0.1282772, 0.1378687, 0.1949436,
  0.06627197, 0.08098289, 0.01256078, 0.07024311, 0.04866307, 0.1205181, 
    0.05860926, 0.05937514, 0.06861805, 0.05111345, 0.03056833, 0.08521538, 
    0.08721055, 0.09659227, 0.1490609, 0.117837, 0.09585873, 0.04945027, 
    0.06248457, 0.07665008, 0.09994003, 0.07565111, 0.02934518, 0.006181668, 
    0.02633024, 0.03565986, 0.09959237, 0.0906182, 0.05704198,
  0.03978861, -1.576975e-05, 0.08197447, 0.002882009, 0.06966291, 0.07755949, 
    0.01967263, 0.003254424, 0.02179931, 0.04964928, 0.03474075, 0.001763113, 
    0.02525341, 0.117153, 0.02904997, 0.04825393, 0.1927246, 0.08104248, 
    0.09250389, 0.08960045, 0.02294324, 0.0005794664, -2.923317e-07, 
    0.0001000967, 0.02883415, 0.2090297, 0.01779424, 0.03959096, 0.07812954,
  0.002303166, 0.09858745, 0.07687477, 0.1256144, 0.1077897, 0.1008637, 
    0.03666326, 0.1161713, 0.001989191, 0.01906406, 0.08429594, 0.02802586, 
    0.04052562, 0.02870922, 0.05717165, 0.03826984, 0.03605191, 0.08860417, 
    0.07703331, 0.064904, 0.03695969, 7.297996e-05, 3.09914e-06, 
    -1.06044e-05, 0.1475609, 0.05306505, 0.01980449, 0.001518719, 0.0001617542,
  6.998011e-07, -6.935616e-05, 0.2292746, 0.08309158, 0.0333875, 0.06538636, 
    0.07110471, 0.05462051, 0.06976555, 0.06274929, 0.1370747, 0.03843685, 
    0.09421509, 0.04314733, 0.06342249, 0.02359908, 0.05529704, 0.01641961, 
    0.02317873, 0.02451142, 0.0006715034, 0.0002195261, 4.050034e-05, 
    0.109495, 0.1752473, 0.06184047, 0.026147, 0.0003710434, 2.47165e-07,
  0.002082796, 0.02216805, 0.001750835, 0.0882555, 0.02451254, 0.01897562, 
    0.02390262, 0.01134855, 0.08444094, 0.2982176, 0.02350577, 0.01202482, 
    0.01144412, 0.03765216, 0.01818487, 0.02168848, 0.009880931, 0.0225353, 
    0.05744538, 0.01528822, 0.04022114, 0.03284364, 0.14319, 0.125271, 
    0.1437597, 0.03635746, 0.03998318, 0.01133761, 0.001698802,
  -2.172387e-05, 1.569782e-06, 4.824404e-06, 0.2251537, 0.01073316, 
    0.02278185, 0.00938121, 0.003129708, 0.01069883, 0.01465672, 0.1484721, 
    0.07051995, 0.03376347, 0.03140828, 0.05211154, 0.06548668, 0.05097855, 
    0.04310865, 0.01855324, 0.03086189, 0.0399644, 0.0143599, 0.02912456, 
    0.02116968, 0.04878686, 0.0157777, -4.55654e-05, 2.099319e-05, 0.000567553,
  1.485555e-06, 4.954414e-07, 1.393116e-07, 2.394402e-08, 0.003850028, 
    1.911212e-05, -1.516396e-06, 0.002437361, -7.848504e-06, 0.007364121, 
    0.1749427, 0.04642613, 0.02444537, 0.009977531, 0.0258748, 0.002656932, 
    0.1234621, -7.319989e-06, 0.002753596, 0.0001597381, 4.09999e-05, 
    0.1154609, 0.02723469, 0.02131979, 0.03698373, 0.09286068, 0.0157844, 
    0.005550936, 0.001360082,
  0.0128145, 0.03210969, 0.03351351, 0.04756818, 0.0455321, 0.04814875, 
    0.03610257, 0.01408373, 0.1729808, 0.1709718, 0.1697921, 0.1011583, 
    0.1069824, 0.13574, 0.1115223, 0.1057533, 0.06660139, 0.1171476, 
    0.08762801, 0.04191643, 0.03224969, 0.08311956, 0.02564379, 0.03580872, 
    0.04716417, 0.04511277, 0.03011082, 0.01630156, 0.003120321,
  0.03124668, 0.04972568, 0.03483267, 0.1024821, 0.01039501, 0.08180822, 
    0.2271882, 0.01848039, 0.009207782, 0.05238229, 0.07886104, 0.1110905, 
    0.1809341, 0.2566565, 0.1812431, 0.1742041, 0.2083215, 0.2364048, 
    0.2595223, 0.2452939, 0.2371741, 0.05488789, 0.1127354, 0.1527375, 
    0.1446712, 0.1232696, 0.1381018, 0.1657683, 0.1666044,
  0.1828123, 0.1146975, 0.1181685, 0.1509776, 0.1616672, 0.1198265, 
    0.2186019, 0.2947287, 0.1239676, 0.1041128, 0.0795896, 0.133771, 
    0.2583294, 0.3303533, 0.3581819, 0.07208347, 0.03220859, 0.1300256, 
    0.2699834, 0.3358315, 0.1431258, 0.1212955, 0.210473, 0.200123, 
    0.2972574, 0.2148612, 0.2765791, 0.2679045, 0.228768,
  0.1982588, 0.2498073, 0.3149122, 0.4042974, 0.4996332, 0.3874814, 
    0.3419002, 0.4350412, 0.3219006, 0.2675446, 0.3033203, 0.1731471, 
    0.2883592, 0.3654317, 0.08767366, 0.08628712, 0.03618971, 0.05822587, 
    0.1821202, 0.2527437, 0.2713713, 0.224657, 0.1491316, 0.1530841, 
    0.1208084, 0.3251434, 0.306201, 0.3299896, 0.2340541,
  0.270525, 0.2548918, 0.4401065, 0.4914449, 0.3312562, 0.2492597, 0.3261619, 
    0.3876334, 0.3830774, 0.2143789, 0.1102369, 0.1712605, 0.1981562, 
    0.1856163, 0.134162, 0.162634, 0.2387544, 0.2234506, 0.1174293, 
    0.2178409, 0.1827545, 0.09831313, 0.09555782, 0.1065181, 0.1228373, 
    0.2668859, 0.2237699, 0.1769792, 0.2575426,
  0.1911159, 0.3090229, 0.2195905, 0.1622817, 0.2847123, 0.3031416, 0.200727, 
    0.2252242, 0.3226224, 0.3087631, 0.2689801, 0.2092806, 0.1928792, 
    0.2418472, 0.2700053, 0.2590819, 0.2326548, 0.2763551, 0.2706693, 
    0.2862897, 0.2307798, 0.2540382, 0.1617665, 0.1100015, 0.06989891, 
    0.01807477, 0.08257736, 0.07422828, 0.1495942,
  0.08843844, 0.08719351, 0.08594857, 0.08470363, 0.0834587, 0.08221376, 
    0.08096882, 0.0651805, 0.07052325, 0.07586601, 0.08120876, 0.08655151, 
    0.09189426, 0.09723701, 0.1073903, 0.1062316, 0.105073, 0.1039143, 
    0.1027557, 0.101597, 0.1004384, 0.1032448, 0.1003056, 0.09736644, 
    0.09442727, 0.09148809, 0.08854892, 0.08560974, 0.0894344,
  0.04479598, 0.04906452, 0.05870517, 0.128722, 0.2090648, 0.3648262, 
    0.2556092, 0.1240837, 0.04532617, 0.0233638, 0.04936586, 0.1321886, 
    0.1386983, 0.2092237, 0.176049, 0.32061, 0.2127116, 0.1937839, 0.2230656, 
    0.2183435, 0.2982514, 0.3616415, 0.1188264, 0.1267353, 0.1545709, 
    0.08749637, 0.0504843, 0.09962048, 0.07376222,
  0.2888491, 0.308057, 0.2387359, 0.2656704, 0.3689359, 0.3872849, 0.4598069, 
    0.4904029, 0.3778789, 0.3359207, 0.2584246, 0.1332948, 0.05843462, 
    0.08740119, 0.2985916, 0.4437069, 0.3633221, 0.3026249, 0.3948705, 
    0.1648466, 0.2249292, 0.3524331, 0.2196576, 0.3226757, 0.2717649, 
    0.178823, 0.2395953, 0.4227592, 0.3591343,
  0.2502649, 0.3441496, 0.3477076, 0.3046366, 0.3683474, 0.2613669, 
    0.3659109, 0.3994782, 0.446438, 0.2979072, 0.230967, 0.3000569, 
    0.2346202, 0.1939851, 0.2277112, 0.1579704, 0.1685073, 0.2623177, 
    0.3364838, 0.3963286, 0.3091449, 0.2887285, 0.2621953, 0.2353777, 
    0.2930705, 0.3354774, 0.2972224, 0.2602577, 0.2508216,
  0.2378074, 0.2236953, 0.251902, 0.2048866, 0.1819215, 0.2320729, 0.243909, 
    0.23879, 0.1655221, 0.2062603, 0.1459077, 0.1249909, 0.2146858, 
    0.2070843, 0.1635296, 0.1828604, 0.1334209, 0.1076438, 0.1345115, 
    0.1996551, 0.1988919, 0.1663329, 0.167933, 0.1344667, 0.07876672, 
    0.1141595, 0.1242733, 0.1641404, 0.1836401,
  0.07486234, 0.09645024, 0.01399016, 0.07262742, 0.06002516, 0.1228044, 
    0.06220508, 0.08127683, 0.08573951, 0.07378034, 0.02311674, 0.1009115, 
    0.1179361, 0.1022751, 0.1515356, 0.106071, 0.07971197, 0.06442342, 
    0.06127666, 0.07148368, 0.1021074, 0.09798978, 0.03416737, 0.00751819, 
    0.01572603, 0.04510932, 0.09134372, 0.07412509, 0.05691675,
  0.04387777, -5.686131e-05, 0.06294043, 0.003513145, 0.07144509, 0.0779192, 
    0.03606343, 0.0005854348, 0.01544914, 0.03449672, 0.01437522, 
    0.002257025, 0.02834342, 0.09412199, 0.02980597, 0.04206511, 0.2040096, 
    0.1005753, 0.1178733, 0.08430936, 0.02872953, 0.005342792, -2.897312e-06, 
    4.874284e-05, 0.02591088, 0.1938259, 0.01828875, 0.05411567, 0.08414863,
  0.01243933, 0.05708919, 0.08308518, 0.123399, 0.105278, 0.08310989, 
    0.0537433, 0.1117528, 0.01240727, 0.02037524, 0.07020225, 0.01096578, 
    0.0391317, 0.02956877, 0.05618048, 0.03576245, 0.03298272, 0.07353652, 
    0.0711435, 0.07025407, 0.06248387, 0.01047708, 1.508946e-06, 
    -6.496641e-05, 0.1499939, 0.05237618, 0.03393082, 0.01804086, 0.007008838,
  3.696224e-07, -0.001886296, 0.1684982, 0.0539778, 0.0282909, 0.05414779, 
    0.0700255, 0.0499116, 0.06345411, 0.05817875, 0.1268852, 0.03338193, 
    0.08018728, 0.03649278, 0.05079518, 0.02480821, 0.06262594, 0.02118936, 
    0.02186991, 0.03407039, 0.003748792, 0.002625223, 1.74152e-05, 0.1152238, 
    0.1412039, 0.04893865, 0.03877473, 0.0005047058, 3.286413e-06,
  0.001037849, 0.01076266, 0.001945946, 0.05308045, 0.02458832, 0.02185818, 
    0.02382828, 0.01567338, 0.09472833, 0.2797846, 0.03022389, 0.01450043, 
    0.01217998, 0.04194349, 0.02081219, 0.02747093, 0.01257775, 0.03084859, 
    0.05637069, 0.02685546, 0.05046646, 0.0405781, 0.1152564, 0.1122497, 
    0.1312352, 0.03470423, 0.03582196, 0.01345172, 0.001431198,
  -7.911503e-06, 2.919043e-07, 1.034289e-06, 0.103919, 0.02461603, 
    0.02473252, 0.01579723, 0.004074128, 0.01772311, 0.02417877, 0.1716406, 
    0.06792118, 0.04226193, 0.0311786, 0.04569576, 0.06428158, 0.05260617, 
    0.03932155, 0.02572209, 0.03628194, 0.03905487, 0.01572667, 0.05044187, 
    0.0362176, 0.0545521, 0.01566189, 0.0001408546, 1.191453e-06, 3.965825e-05,
  5.580641e-07, 2.12881e-07, 7.065255e-08, 6.904577e-05, 0.0006471379, 
    2.190859e-05, 0.001974293, 0.002470256, 0.008027958, 0.01096701, 
    0.1314656, 0.07165575, 0.03830761, 0.01359152, 0.03084429, 0.004814246, 
    0.119329, 0.001460571, 0.0036342, 3.64606e-06, 1.632583e-05, 0.1219042, 
    0.03055819, 0.02309137, 0.03793835, 0.07923254, 0.03599187, 0.004502826, 
    0.0001524594,
  0.01630123, 0.0226472, 0.09997852, 0.06313574, 0.04922674, 0.04268254, 
    0.01820586, 0.01688899, 0.1620807, 0.1532304, 0.1619213, 0.1098676, 
    0.1171218, 0.1358303, 0.1434225, 0.1198772, 0.07614417, 0.1139457, 
    0.1125714, 0.04610926, 0.02729432, 0.1007697, 0.04015172, 0.04145893, 
    0.05293046, 0.05080296, 0.03615503, 0.04325208, 0.002386709,
  0.02074085, 0.05038906, 0.03770638, 0.1211917, 0.0165493, 0.05108213, 
    0.2221999, 0.008794966, 0.003308388, 0.05662167, 0.05358528, 0.1198506, 
    0.1982341, 0.276804, 0.1853642, 0.1741645, 0.243256, 0.2481399, 0.263345, 
    0.2647536, 0.2249021, 0.04777856, 0.1280567, 0.1831946, 0.1466986, 
    0.1543121, 0.1549657, 0.1790732, 0.1896735,
  0.1712907, 0.1355455, 0.1371267, 0.170586, 0.1186498, 0.1400089, 0.198227, 
    0.3002112, 0.1175416, 0.09093844, 0.07490257, 0.1344363, 0.2381051, 
    0.3798894, 0.4056518, 0.07333168, 0.0584601, 0.1429281, 0.3084632, 
    0.3611869, 0.1423432, 0.08259446, 0.2041016, 0.2284675, 0.3044099, 
    0.2254154, 0.3191475, 0.2862751, 0.2139034,
  0.197093, 0.2220028, 0.3089914, 0.3604081, 0.472404, 0.3812039, 0.3199414, 
    0.407173, 0.3382698, 0.2883292, 0.3361607, 0.179182, 0.2905613, 0.35882, 
    0.1296645, 0.2031655, 0.03504102, 0.05208192, 0.2545192, 0.2665234, 
    0.2556747, 0.2146563, 0.1188741, 0.1558202, 0.1085288, 0.2984463, 
    0.3243506, 0.3354799, 0.2369647,
  0.257049, 0.2865469, 0.4173175, 0.5078992, 0.315021, 0.2235123, 0.3002876, 
    0.3982845, 0.3840843, 0.2101399, 0.1183716, 0.1918975, 0.1751908, 
    0.2182485, 0.1504663, 0.1694385, 0.2625426, 0.2745574, 0.1429862, 
    0.2411242, 0.1931866, 0.09831464, 0.1104535, 0.08241992, 0.09186866, 
    0.3586361, 0.2385146, 0.2379495, 0.2764761,
  0.2853759, 0.2900118, 0.1888431, 0.1420493, 0.2849201, 0.3078047, 
    0.2110246, 0.2451435, 0.3364168, 0.3005355, 0.2778327, 0.2244118, 
    0.2034208, 0.2149004, 0.2551083, 0.2663437, 0.2220873, 0.2713538, 
    0.2981293, 0.312315, 0.2589975, 0.2820253, 0.1694055, 0.1032135, 
    0.06557978, 0.03564811, 0.08168809, 0.09500507, 0.1786184,
  0.09118559, 0.08987503, 0.08856449, 0.08725393, 0.08594338, 0.08463282, 
    0.08332227, 0.06965925, 0.07246201, 0.07526477, 0.07806753, 0.08087029, 
    0.08367305, 0.08647581, 0.09287366, 0.09208158, 0.09128951, 0.09049743, 
    0.08970535, 0.08891328, 0.0881212, 0.08893038, 0.08823025, 0.08753012, 
    0.08682999, 0.08612986, 0.08542974, 0.0847296, 0.09223403,
  0.04027409, 0.04334169, 0.05650988, 0.1508582, 0.2336529, 0.3891053, 
    0.2727906, 0.1426401, 0.07468894, 0.02408934, 0.04327344, 0.1237823, 
    0.1643531, 0.1755342, 0.1727803, 0.2048013, 0.1963442, 0.1823692, 
    0.1997122, 0.2791408, 0.2846861, 0.3269551, 0.1422261, 0.05816443, 
    0.1781408, 0.1379546, 0.1794195, 0.0909545, 0.06401623,
  0.2551487, 0.2396231, 0.2209529, 0.2203057, 0.3784409, 0.471932, 0.4167526, 
    0.4802836, 0.370283, 0.3183787, 0.2520046, 0.1008956, 0.06009563, 
    0.09434782, 0.2992194, 0.3954038, 0.388256, 0.2770758, 0.3624663, 
    0.276345, 0.2900431, 0.2925382, 0.2336935, 0.2538042, 0.3024932, 
    0.1443432, 0.2314804, 0.3462003, 0.3235843,
  0.2998962, 0.3074925, 0.329104, 0.2876815, 0.3172494, 0.2339703, 0.3138901, 
    0.3671687, 0.355803, 0.2960661, 0.2270175, 0.2287762, 0.2149514, 
    0.1720965, 0.2760347, 0.1975388, 0.1582499, 0.2677266, 0.3344387, 
    0.3939275, 0.3188615, 0.2583964, 0.2495808, 0.2412977, 0.2589414, 
    0.2796719, 0.2650612, 0.2769621, 0.2298744,
  0.25847, 0.2352134, 0.273326, 0.2166502, 0.1932415, 0.2593461, 0.247081, 
    0.2371256, 0.1735255, 0.2342592, 0.1658967, 0.1618846, 0.2589221, 
    0.2296591, 0.1508197, 0.1782013, 0.1285039, 0.1112956, 0.1715945, 
    0.2312945, 0.2478128, 0.194593, 0.1746954, 0.1515994, 0.04967188, 
    0.08691511, 0.1458797, 0.1461206, 0.1876256,
  0.07843145, 0.1033066, 0.02388946, 0.09165682, 0.07859937, 0.1314415, 
    0.0610407, 0.1094659, 0.0914437, 0.05567495, 0.02665329, 0.1168969, 
    0.1275339, 0.100501, 0.1461117, 0.1138013, 0.07921129, 0.06815511, 
    0.05544524, 0.07868306, 0.1205398, 0.09171795, 0.04762834, 0.009173157, 
    0.008962222, 0.05050151, 0.07931162, 0.0777985, 0.06499578,
  0.06387014, -6.96621e-05, 0.0769881, 0.01256856, 0.1147665, 0.08462922, 
    0.04902678, 0.01144741, 0.01817873, 0.03539021, 0.01003589, 0.0003049983, 
    0.01648135, 0.0910242, 0.03949839, 0.04400281, 0.197996, 0.1225349, 
    0.1325905, 0.08631217, 0.03868128, 0.01776902, 0.0001159056, 
    3.760951e-05, 0.01935371, 0.1852152, 0.02202058, 0.05819657, 0.1147223,
  0.01002515, 0.032872, 0.08269003, 0.1066225, 0.09007633, 0.06925799, 
    0.06422617, 0.1171943, 0.01361223, 0.03192938, 0.06183371, 0.008932303, 
    0.04336308, 0.02971943, 0.06089376, 0.03812695, 0.02862131, 0.05759399, 
    0.05736389, 0.04564242, 0.07946307, 0.07292458, 6.353773e-06, 
    5.363838e-05, 0.1410637, 0.05638767, 0.03597147, 0.06318698, 0.03953866,
  3.843707e-06, -0.0006016883, 0.133472, 0.04786322, 0.0230247, 0.04432616, 
    0.06134332, 0.04273621, 0.05485789, 0.05457224, 0.1107339, 0.02660243, 
    0.06928501, 0.03051099, 0.03919915, 0.02228478, 0.04962895, 0.02545013, 
    0.02524205, 0.0340786, 0.003374848, 0.006789654, 0.001600499, 0.1172762, 
    0.1230492, 0.0378433, 0.04501443, 0.002027922, 0.001558936,
  0.001032805, 0.008048079, 0.001836202, 0.01838357, 0.03002794, 0.02557909, 
    0.02524817, 0.01838421, 0.1103192, 0.2914012, 0.03477935, 0.01739435, 
    0.01282165, 0.03770498, 0.0216881, 0.02722785, 0.02069092, 0.04011792, 
    0.06078819, 0.04389669, 0.06308542, 0.04575051, 0.1090584, 0.09914634, 
    0.1221288, 0.03014589, 0.03326597, 0.01544773, 0.001351877,
  -2.49447e-06, 6.97207e-08, 2.039953e-07, 0.03190407, 0.03593281, 0.0221519, 
    0.02082466, 0.01233544, 0.02950376, 0.03317388, 0.1663821, 0.06491898, 
    0.04016045, 0.03514621, 0.05148336, 0.05853818, 0.05523018, 0.02595094, 
    0.0343697, 0.04036426, 0.03658883, 0.01697092, 0.06342077, 0.08181019, 
    0.05491937, 0.01630464, 0.0006160622, 1.78784e-07, 3.584796e-05,
  2.234821e-07, 1.000575e-07, 3.424909e-08, 0.001540898, -7.772825e-06, 
    3.464958e-05, 0.003825721, 0.00372188, 0.006400507, 0.01913943, 
    0.09401901, 0.1210479, 0.03210286, 0.03457585, 0.05124838, 0.01514718, 
    0.1198065, 0.005017782, 0.006434508, 7.531636e-07, 6.556765e-06, 
    0.1208968, 0.02830487, 0.03364675, 0.02882353, 0.06606584, 0.0523468, 
    0.002193939, 9.371539e-06,
  0.01678853, 0.03250438, 0.1144082, 0.0184227, 0.06108857, 0.0402919, 
    0.003661698, 0.01175433, 0.149366, 0.16287, 0.1743959, 0.1301226, 
    0.1362331, 0.1311402, 0.1567064, 0.1318363, 0.08855671, 0.1068113, 
    0.1267163, 0.04169695, 0.02500747, 0.09986972, 0.05996974, 0.05442575, 
    0.04933805, 0.05374432, 0.04621882, 0.0630117, 0.000149157,
  0.01188411, 0.05016622, 0.05015796, 0.1302632, 0.02025912, 0.03045839, 
    0.2134057, 0.001169769, 0.0004520742, 0.06167835, 0.0370895, 0.1762959, 
    0.2386857, 0.2920085, 0.1899371, 0.2128182, 0.3127543, 0.273797, 
    0.285096, 0.2868551, 0.2019773, 0.05136856, 0.1559682, 0.197755, 
    0.148607, 0.1496061, 0.16243, 0.1745203, 0.218227,
  0.1589499, 0.1576285, 0.126801, 0.172766, 0.08721273, 0.1756639, 0.2153047, 
    0.3030882, 0.09528147, 0.07443437, 0.078471, 0.1310337, 0.188372, 
    0.3434183, 0.405613, 0.08923945, 0.1129619, 0.179978, 0.3449383, 
    0.3914829, 0.131579, 0.07766776, 0.1946918, 0.2443093, 0.3138078, 
    0.291935, 0.3497066, 0.3057095, 0.2004291,
  0.2019941, 0.1960709, 0.3378057, 0.3561636, 0.460534, 0.3686596, 0.380592, 
    0.3720039, 0.3725592, 0.2847784, 0.2817042, 0.1787959, 0.2967517, 
    0.4733425, 0.2763111, 0.1845481, 0.048145, 0.04296611, 0.2680007, 
    0.2904558, 0.2352488, 0.2111532, 0.09991486, 0.1605898, 0.1102057, 
    0.3078224, 0.3066224, 0.3162267, 0.2521616,
  0.2296596, 0.2688224, 0.4196965, 0.4736513, 0.240011, 0.1649932, 0.2705265, 
    0.4030701, 0.3838364, 0.2162642, 0.1265814, 0.1997988, 0.159478, 
    0.244191, 0.1830697, 0.1905593, 0.2806341, 0.3179294, 0.1492272, 
    0.2725426, 0.2006749, 0.1137552, 0.1385742, 0.0545168, 0.06701406, 
    0.3692968, 0.2507134, 0.2362585, 0.2954391,
  0.2506896, 0.2280884, 0.1629062, 0.1436454, 0.2523761, 0.2883475, 
    0.2197733, 0.2506609, 0.3681961, 0.3707342, 0.3350815, 0.2584192, 
    0.2083505, 0.2120535, 0.2278255, 0.2467366, 0.2272598, 0.3057486, 
    0.3240972, 0.3614372, 0.3193824, 0.2970379, 0.1809572, 0.0956853, 
    0.06605098, 0.04647893, 0.08270445, 0.121914, 0.2928842,
  0.100023, 0.09964643, 0.09926987, 0.09889331, 0.09851675, 0.0981402, 
    0.09776364, 0.08646572, 0.08586926, 0.0852728, 0.08467633, 0.08407987, 
    0.08348341, 0.08288695, 0.08415243, 0.08462586, 0.08509929, 0.08557272, 
    0.08604614, 0.08651958, 0.086993, 0.08883761, 0.0893372, 0.08983679, 
    0.09033638, 0.09083597, 0.09133556, 0.09183515, 0.1003242,
  0.04200535, 0.04575753, 0.06179339, 0.1742972, 0.2569498, 0.4005759, 
    0.2840261, 0.1501332, 0.09389964, 0.0254397, 0.04178349, 0.1152478, 
    0.2264956, 0.1029549, 0.08059014, 0.1052913, 0.1838937, 0.1768435, 
    0.1751382, 0.2556693, 0.3197881, 0.3281256, 0.1655091, 0.03949178, 
    0.1561829, 0.2314585, 0.2534779, 0.08820063, 0.05477932,
  0.2752677, 0.3087711, 0.2214221, 0.1776226, 0.3530611, 0.4319065, 
    0.3271244, 0.5287579, 0.3798185, 0.3224815, 0.2377875, 0.04916936, 
    0.05128041, 0.137472, 0.4142264, 0.4085622, 0.3747586, 0.3568416, 
    0.4552749, 0.357036, 0.3278659, 0.3061751, 0.222597, 0.2695459, 
    0.3125902, 0.2064466, 0.2355679, 0.2779034, 0.3367698,
  0.3237499, 0.3319608, 0.294352, 0.3202773, 0.3274081, 0.2644821, 0.3292227, 
    0.3960322, 0.4018971, 0.3811513, 0.1981781, 0.2573231, 0.211518, 
    0.2352948, 0.3278875, 0.2383569, 0.2263046, 0.2819287, 0.3541019, 
    0.4015185, 0.3298256, 0.2540569, 0.2849914, 0.3123647, 0.2704423, 
    0.2992537, 0.2590423, 0.3126584, 0.3211403,
  0.2700753, 0.2399594, 0.2766975, 0.2456483, 0.2328067, 0.2766559, 
    0.2686855, 0.2706581, 0.2009443, 0.2820616, 0.2038522, 0.2039022, 
    0.2783531, 0.2276728, 0.1803888, 0.1892179, 0.1459602, 0.1443892, 
    0.234312, 0.3085947, 0.2611947, 0.2650968, 0.219078, 0.1574129, 
    0.03562604, 0.07745401, 0.1705504, 0.1620339, 0.2309206,
  0.09026487, 0.1276975, 0.08820157, 0.1103396, 0.1277396, 0.1576604, 
    0.0857984, 0.1361241, 0.1362193, 0.05938425, 0.07355754, 0.1692846, 
    0.1276235, 0.1144837, 0.1439279, 0.1620002, 0.1102346, 0.07636176, 
    0.08426614, 0.1084822, 0.1704225, 0.1568662, 0.07303704, 0.01234346, 
    0.02083199, 0.0764522, 0.08196247, 0.08732636, 0.09646192,
  0.08983096, -3.040843e-06, 0.0760192, 0.0574731, 0.1158589, 0.08969749, 
    0.06480998, 0.09191599, 0.01830255, 0.03484687, 0.007797674, 
    7.956944e-05, 0.0139994, 0.09635647, 0.06525181, 0.05213398, 0.2149728, 
    0.1627501, 0.1003631, 0.09256632, 0.0433423, 0.03598088, 0.004961656, 
    5.348936e-05, 0.01502582, 0.1736048, 0.0260163, 0.0606979, 0.1221109,
  0.009848047, 0.0206751, 0.08082313, 0.09638278, 0.07462321, 0.05768709, 
    0.04965215, 0.1245575, 0.02353917, 0.03549366, 0.04425849, 0.01006239, 
    0.03970081, 0.03495159, 0.06218355, 0.03678111, 0.02655273, 0.04540168, 
    0.04235478, 0.030998, 0.05783466, 0.09969164, 0.005836942, 0.0002992971, 
    0.1297733, 0.05615954, 0.02595013, 0.04358912, 0.09920389,
  0.001604791, -0.00025179, 0.109076, 0.04587843, 0.02147237, 0.03876382, 
    0.05110463, 0.03509225, 0.04753408, 0.04116999, 0.09703054, 0.02122221, 
    0.06087773, 0.02421875, 0.03330831, 0.02124571, 0.04368521, 0.02646691, 
    0.02664746, 0.03323992, 0.01176087, 0.01253296, 0.01920836, 0.1133584, 
    0.1038559, 0.03295543, 0.04791531, 0.01765056, 0.01496496,
  0.001304616, 0.0109574, 0.001726005, 0.005002949, 0.03978865, 0.05621497, 
    0.02969318, 0.01968776, 0.1271834, 0.2943813, 0.03416502, 0.01761679, 
    0.01513306, 0.03181286, 0.02225998, 0.02567099, 0.02365433, 0.03962477, 
    0.07078433, 0.05504816, 0.07650774, 0.04057835, 0.09449127, 0.09067361, 
    0.106675, 0.02770242, 0.02932716, 0.01682533, 0.001859183,
  -1.803579e-07, 2.047681e-08, 2.814716e-08, 0.01609263, 0.05684531, 
    0.01890029, 0.02300439, 0.02048281, 0.02253998, 0.03502211, 0.1694791, 
    0.06182447, 0.04233854, 0.03664884, 0.05402024, 0.04817767, 0.05870992, 
    0.02744593, 0.04548676, 0.03649851, 0.03243568, 0.01793656, 0.07846233, 
    0.1023539, 0.05409381, 0.01808462, 0.01028836, 9.153464e-08, 3.283264e-05,
  1.347257e-07, 6.069798e-08, 1.429948e-08, 0.01557652, -2.335005e-06, 
    0.0003307885, 0.00057075, 0.008092741, 0.003203506, 0.06934321, 
    0.09485666, 0.127168, 0.03163102, 0.04433415, 0.07214791, 0.03507751, 
    0.1178258, 0.01295252, 0.01632244, 7.755565e-06, 4.128849e-06, 0.1505904, 
    0.04521712, 0.0462149, 0.0305872, 0.05121153, 0.05111515, 5.154346e-07, 
    3.050098e-06,
  0.01442538, 0.0215971, 0.07528705, 0.00929517, 0.0478266, 0.0394683, 
    -0.00107847, 0.003528239, 0.1356484, 0.15294, 0.2153023, 0.2136535, 
    0.1676771, 0.1607348, 0.2060523, 0.1548595, 0.1150481, 0.1230959, 
    0.1546667, 0.05264441, 0.02260696, 0.09436445, 0.06829585, 0.09882988, 
    0.05473129, 0.05600061, 0.06966434, 0.08920903, 0.003826725,
  0.01089028, 0.04725624, 0.0870712, 0.1567504, 0.05712475, 0.03006014, 
    0.1986439, 0.0003824455, -0.0002366729, 0.04939275, 0.03857089, 
    0.2643645, 0.3574393, 0.2957404, 0.234178, 0.2587889, 0.3642296, 
    0.3114229, 0.3366709, 0.3180847, 0.2008543, 0.05300447, 0.1919615, 
    0.2186592, 0.2082738, 0.1764826, 0.2264314, 0.221071, 0.2632145,
  0.1829304, 0.1871321, 0.1048392, 0.1657723, 0.1147788, 0.1755153, 
    0.2217999, 0.3103853, 0.07172931, 0.05279712, 0.05183728, 0.1244118, 
    0.2137641, 0.2972353, 0.3962185, 0.1535503, 0.1738368, 0.2471766, 
    0.3209144, 0.4719807, 0.1239493, 0.07809551, 0.2086413, 0.2638872, 
    0.3168954, 0.4099886, 0.3417677, 0.2808988, 0.2013383,
  0.1976508, 0.2325403, 0.336736, 0.3340035, 0.4644795, 0.3751281, 0.339836, 
    0.3989518, 0.3752005, 0.294163, 0.3063573, 0.1808461, 0.3069708, 
    0.5214522, 0.2672156, 0.1240517, 0.05845525, 0.03330984, 0.2603265, 
    0.3069492, 0.2559465, 0.2367854, 0.1070339, 0.1612091, 0.1540043, 
    0.3022273, 0.3024869, 0.3051482, 0.2593916,
  0.2874358, 0.2665306, 0.3503768, 0.5056952, 0.2431239, 0.1879932, 
    0.2829689, 0.4011589, 0.3860584, 0.2178954, 0.1393568, 0.1912487, 
    0.1487926, 0.2608933, 0.2019382, 0.2203963, 0.300446, 0.3531374, 
    0.1598714, 0.2757195, 0.2216122, 0.1367253, 0.1467236, 0.04457596, 
    0.04417468, 0.3703107, 0.2584719, 0.2014568, 0.3019369,
  0.1711775, 0.1848701, 0.1638295, 0.1337517, 0.2332564, 0.2909281, 
    0.2269286, 0.2555617, 0.3993196, 0.406399, 0.3554332, 0.2573667, 
    0.2034529, 0.232041, 0.2280743, 0.2612294, 0.2586506, 0.3401496, 
    0.339174, 0.3800465, 0.33364, 0.3218206, 0.1718801, 0.0917372, 0.0732675, 
    0.03875196, 0.08018203, 0.1453098, 0.2944157,
  0.1149001, 0.1144186, 0.113937, 0.1134555, 0.1129739, 0.1124924, 0.1120108, 
    0.1093466, 0.1065991, 0.1038516, 0.1011042, 0.09835673, 0.09560928, 
    0.09286182, 0.08929513, 0.09214962, 0.09500409, 0.09785857, 0.100713, 
    0.1035675, 0.106422, 0.1150955, 0.11547, 0.1158445, 0.1162191, 0.1165936, 
    0.1169681, 0.1173426, 0.1152853,
  0.04214699, 0.04915907, 0.06771241, 0.1915519, 0.2883475, 0.403034, 
    0.2974553, 0.1556747, 0.1190485, 0.03317852, 0.03668311, 0.1115068, 
    0.2435899, 0.03724035, 0.104001, 0.09660888, 0.1500035, 0.1832702, 
    0.1829314, 0.2466075, 0.3476881, 0.3183484, 0.1916261, 0.04770934, 
    0.1642796, 0.2098632, 0.2064393, 0.05987692, 0.0461896,
  0.3226331, 0.2770357, 0.2115662, 0.142903, 0.2932619, 0.4161141, 0.2382752, 
    0.5523561, 0.3923278, 0.3189138, 0.1952017, 0.02216725, 0.03237374, 
    0.1840737, 0.5096753, 0.4322777, 0.388539, 0.4758227, 0.4643879, 
    0.5218628, 0.3933322, 0.3593136, 0.3248064, 0.2812082, 0.2952514, 
    0.3880873, 0.3488036, 0.3571884, 0.4182454,
  0.3198026, 0.3266629, 0.3066556, 0.3531379, 0.3676807, 0.326053, 0.4402603, 
    0.4282365, 0.4544357, 0.4288977, 0.2436484, 0.3319233, 0.3272269, 
    0.3734607, 0.4010633, 0.2813128, 0.2553579, 0.3006, 0.3769369, 0.4205915, 
    0.3462613, 0.2908135, 0.3620834, 0.4013567, 0.3277216, 0.3906972, 
    0.3679582, 0.3912284, 0.4342546,
  0.3385228, 0.3011148, 0.3207219, 0.2731339, 0.2781081, 0.3331638, 0.306511, 
    0.3042945, 0.2244194, 0.3456504, 0.3024223, 0.2900746, 0.2983502, 
    0.2402452, 0.1921626, 0.2669804, 0.206726, 0.1919822, 0.2876972, 
    0.3756979, 0.305012, 0.3048842, 0.2968566, 0.1806017, 0.02289465, 
    0.0978992, 0.196402, 0.2253879, 0.3198474,
  0.1562854, 0.220399, 0.1946006, 0.1757853, 0.2065354, 0.2034462, 0.1888817, 
    0.1778872, 0.1747149, 0.09587038, 0.1459082, 0.2449974, 0.189438, 
    0.134625, 0.1802768, 0.2158685, 0.1560168, 0.1228016, 0.1519607, 
    0.2206341, 0.2464896, 0.180144, 0.1628231, 0.01751116, 0.02949597, 
    0.1324847, 0.1218676, 0.09947108, 0.1440974,
  0.1252371, 0.004826966, 0.06476237, 0.0941796, 0.1117763, 0.1036397, 
    0.06770434, 0.1433187, 0.1022906, 0.0344546, 0.007166575, 0.0002034664, 
    0.009010219, 0.114281, 0.08977818, 0.07625996, 0.2102551, 0.1807538, 
    0.09036579, 0.09659221, 0.04412593, 0.09588914, 0.05703204, 0.000173695, 
    0.01866323, 0.1538161, 0.02674042, 0.05591621, 0.1211229,
  0.06864902, 0.01659989, 0.05278147, 0.0934399, 0.06513911, 0.04872595, 
    0.05238226, 0.1203752, 0.03268581, 0.02763818, 0.03469129, 0.009254703, 
    0.04088623, 0.0456804, 0.05479413, 0.03459899, 0.02617067, 0.03929722, 
    0.03325059, 0.03371878, 0.03853822, 0.1568293, 0.09033699, 0.0002556368, 
    0.1134415, 0.05832816, 0.02671052, 0.03494688, 0.1001491,
  0.02610911, 0.0004014004, 0.08539832, 0.05315197, 0.02336821, 0.03405416, 
    0.04662221, 0.03267796, 0.04228986, 0.03102533, 0.08765634, 0.01887174, 
    0.05496348, 0.02151326, 0.03030209, 0.02596416, 0.04086516, 0.02797178, 
    0.0280554, 0.03132927, 0.02344103, 0.0132924, 0.05928959, 0.1039261, 
    0.08539764, 0.03027885, 0.05347505, 0.03598607, 0.0533081,
  0.002112117, 0.01300357, 0.001244097, 0.002255955, 0.047075, 0.04563057, 
    0.03362135, 0.02097087, 0.1271635, 0.2653788, 0.03197369, 0.01962742, 
    0.0194018, 0.03144406, 0.02582506, 0.02727339, 0.02289952, 0.0354962, 
    0.06474607, 0.04789404, 0.07112996, 0.03173528, 0.07505513, 0.07881498, 
    0.09828372, 0.0280262, 0.02830185, 0.02134899, 0.003898057,
  -1.181271e-07, 6.446386e-09, 7.427078e-09, 0.005020173, 0.1143228, 
    0.02796544, 0.02814866, 0.04514031, 0.01815413, 0.03933739, 0.144938, 
    0.05979866, 0.05275824, 0.06518572, 0.05527414, 0.04858678, 0.06325916, 
    0.03703119, 0.06357908, 0.04120219, 0.03295584, 0.02266482, 0.1137405, 
    0.1443932, 0.05528695, 0.02276556, 0.02287664, 1.87494e-07, 2.979392e-05,
  8.937391e-08, 5.117648e-08, 5.942052e-09, 0.002613488, 3.340346e-08, 
    0.0353264, 0.0001405453, 0.01516073, 0.006650476, 0.1266184, 0.07534067, 
    0.1480639, 0.06964988, 0.09813377, 0.105171, 0.05029053, 0.1285678, 
    0.02359558, 0.06264763, 0.006010299, 3.371382e-05, 0.1794314, 0.04722223, 
    0.03631564, 0.04752783, 0.06609177, 0.09810924, 0.04416541, 1.407157e-06,
  0.003608972, 0.01301671, 0.05244473, 0.006247552, 0.03549311, 0.03980587, 
    -0.002002422, 0.001121283, 0.1373499, 0.1479277, 0.2657389, 0.2643915, 
    0.1776338, 0.1604812, 0.1936163, 0.1605467, 0.1672276, 0.1501289, 
    0.2409844, 0.05652084, 0.02259407, 0.1230932, 0.08202827, 0.1476415, 
    0.06024583, 0.06386974, 0.1237568, 0.08768709, 0.01074431,
  0.01356397, 0.05006199, 0.0853739, 0.1908172, 0.09695526, 0.0690869, 
    0.1813466, -1.050023e-05, -0.0003097642, 0.03746726, 0.03192912, 
    0.3158332, 0.4589159, 0.3125283, 0.2418558, 0.3089624, 0.4378864, 
    0.37463, 0.3023273, 0.3472346, 0.2238527, 0.05738277, 0.2262567, 
    0.2314456, 0.3306938, 0.3096645, 0.2934203, 0.230071, 0.2672221,
  0.1907582, 0.205135, 0.1369647, 0.1670299, 0.1395666, 0.1802251, 0.2721637, 
    0.3249124, 0.05858959, 0.04037631, 0.02924054, 0.1187722, 0.2619603, 
    0.4158901, 0.4700736, 0.3276152, 0.3413512, 0.3270948, 0.3036759, 
    0.5194068, 0.1162655, 0.09798753, 0.2396975, 0.297805, 0.3057816, 
    0.4923652, 0.3153041, 0.2389815, 0.1687595,
  0.2070597, 0.2889653, 0.3304919, 0.3540478, 0.4658744, 0.4270455, 
    0.4328003, 0.441907, 0.39054, 0.3469391, 0.3289303, 0.1963857, 0.2867834, 
    0.5528006, 0.3584691, 0.1652418, 0.05529898, 0.02652201, 0.2570076, 
    0.343994, 0.28852, 0.2646624, 0.1245658, 0.1736453, 0.3190444, 0.3015713, 
    0.2585577, 0.2929096, 0.221491,
  0.4002645, 0.2746708, 0.3773535, 0.5631998, 0.2902761, 0.2534746, 
    0.2660281, 0.4029759, 0.3940021, 0.22055, 0.150759, 0.1740884, 0.1657536, 
    0.258674, 0.2312615, 0.2375782, 0.3788523, 0.3859047, 0.1893333, 
    0.2954799, 0.2512076, 0.1600353, 0.152767, 0.03936071, 0.04094462, 
    0.3557989, 0.2669287, 0.2095712, 0.3701986,
  0.1637858, 0.1435338, 0.1556034, 0.1100181, 0.2291182, 0.3423776, 
    0.2612041, 0.2838032, 0.4290824, 0.4237525, 0.391446, 0.2531678, 
    0.2145288, 0.2353325, 0.2412855, 0.284595, 0.3120694, 0.3798205, 
    0.3422048, 0.3788858, 0.3482803, 0.3380531, 0.1769715, 0.08984216, 
    0.07835505, 0.04359968, 0.08346464, 0.1851001, 0.2534564,
  0.1242735, 0.1244703, 0.1246671, 0.1248639, 0.1250607, 0.1252574, 
    0.1254542, 0.120677, 0.1169274, 0.1131779, 0.1094283, 0.1056787, 
    0.1019291, 0.09817955, 0.09734733, 0.09991086, 0.1024744, 0.1050379, 
    0.1076014, 0.110165, 0.1127285, 0.1134094, 0.1143987, 0.1153879, 
    0.1163772, 0.1173665, 0.1183557, 0.119345, 0.1241161,
  0.03330694, 0.05728827, 0.06718411, 0.2091344, 0.3241329, 0.4250657, 
    0.3081908, 0.1708653, 0.1381964, 0.04436061, 0.02530947, 0.1239827, 
    0.2867143, -0.00239309, 0.1670047, 0.1013261, 0.09087842, 0.1593713, 
    0.2473812, 0.2343108, 0.3407246, 0.324516, 0.1922379, 0.09308981, 0.289, 
    0.275125, 0.1111645, 0.03453907, 0.04572086,
  0.3572593, 0.2772193, 0.2625612, 0.1543581, 0.2375095, 0.4040053, 
    0.1740947, 0.5400177, 0.3865286, 0.302474, 0.1532086, 0.008884742, 
    0.02385746, 0.1914372, 0.4227385, 0.4207974, 0.3533297, 0.4641509, 
    0.4829175, 0.4641355, 0.4143735, 0.4042785, 0.3541507, 0.2841522, 
    0.3355254, 0.4471653, 0.3897622, 0.4258711, 0.4891351,
  0.3727665, 0.3807476, 0.3510371, 0.369141, 0.3651358, 0.3757405, 0.5049042, 
    0.5232851, 0.5069129, 0.4782106, 0.347357, 0.4052247, 0.4459599, 
    0.4661412, 0.5118753, 0.3909208, 0.2854108, 0.3806077, 0.3876483, 
    0.4097495, 0.3347757, 0.3218212, 0.3661204, 0.3998811, 0.3762958, 
    0.4941866, 0.4837598, 0.3925433, 0.4458723,
  0.398588, 0.3902155, 0.3848299, 0.3082501, 0.3055576, 0.3877477, 0.3555827, 
    0.3648227, 0.4233282, 0.4330009, 0.4457668, 0.3730175, 0.3705218, 
    0.2282923, 0.3431812, 0.3551582, 0.3555247, 0.3819514, 0.392452, 
    0.4159988, 0.3213745, 0.2539988, 0.2896663, 0.206299, 0.01694714, 
    0.1357515, 0.2808807, 0.3003226, 0.3414797,
  0.2240227, 0.2747354, 0.2259831, 0.2504029, 0.2565355, 0.2757572, 
    0.1917724, 0.1873178, 0.3714131, 0.2046253, 0.2715831, 0.3714064, 
    0.1936682, 0.1454189, 0.1822234, 0.2692689, 0.1970426, 0.2400973, 
    0.2904457, 0.2400858, 0.2142769, 0.1885733, 0.2468054, 0.02384678, 
    0.01991535, 0.1642451, 0.1806849, 0.1672988, 0.2729656,
  0.2140594, 0.05707545, 0.05227721, 0.1137132, 0.1101732, 0.1195815, 
    0.0795579, 0.1313125, 0.2790742, 0.04038144, 0.006210847, 2.348737e-05, 
    0.003246302, 0.173108, 0.08529823, 0.09247679, 0.2032004, 0.2306527, 
    0.09262264, 0.09811724, 0.05103844, 0.2219725, 0.2234245, 0.0004194663, 
    0.02348274, 0.1459889, 0.04229156, 0.0629459, 0.1138035,
  0.2298094, 0.02117303, 0.03244296, 0.09273621, 0.06111249, 0.05092665, 
    0.06112655, 0.1248769, 0.07687178, 0.04536233, 0.0265397, 0.005891994, 
    0.03935618, 0.06083861, 0.0521281, 0.0384275, 0.0305047, 0.03527877, 
    0.05859677, 0.04500704, 0.0425212, 0.178904, 0.2287843, 0.001205563, 
    0.09198318, 0.04305496, 0.03490245, 0.03768144, 0.1073632,
  0.09329771, 0.007590664, 0.06233101, 0.06886291, 0.02871815, 0.03510724, 
    0.04553509, 0.04366944, 0.04894982, 0.02585634, 0.07734211, 0.02004846, 
    0.05177221, 0.02247601, 0.03227003, 0.02710707, 0.05291841, 0.04143091, 
    0.05878805, 0.04247303, 0.05246922, 0.02497352, 0.07918085, 0.08633556, 
    0.0676368, 0.01620668, 0.07074338, 0.05567802, 0.07457545,
  0.004467921, 0.01040143, 0.0004980002, 0.000721855, 0.05383363, 0.04592398, 
    0.05296977, 0.03393245, 0.1188668, 0.210576, 0.0305572, 0.0246323, 
    0.02744493, 0.04193601, 0.04468252, 0.03122165, 0.02324586, 0.02777107, 
    0.05414344, 0.0366191, 0.05791669, 0.03559453, 0.0774183, 0.05752249, 
    0.08271953, 0.03476116, 0.03201163, 0.03087974, 0.01067962,
  -8.582038e-08, 2.803948e-09, 1.597076e-09, 0.0003255678, 0.1092013, 
    0.1793403, 0.01726111, 0.1043404, 0.0151329, 0.0817603, 0.1338195, 
    0.0673653, 0.07596775, 0.1101511, 0.07283435, 0.05214015, 0.07152604, 
    0.05168126, 0.06766864, 0.04941222, 0.04090969, 0.03645194, 0.1462736, 
    0.1416937, 0.07752107, 0.04491248, 0.07140601, 1.972182e-07, 1.783604e-05,
  6.041262e-08, 3.472083e-08, 2.670433e-09, 0.009824004, -4.33094e-08, 
    0.01798343, 7.332465e-05, 0.01649413, 0.005691563, 0.1890402, 0.1105497, 
    0.1970885, 0.1464009, 0.1562361, 0.2036417, 0.06274402, 0.1489221, 
    0.05450071, 0.1256341, 0.1718055, 0.01388519, 0.2233302, 0.0429507, 
    0.03160054, 0.05659681, 0.09416214, 0.03865236, 0.05441255, 5.911589e-07,
  0.0002775643, 0.01064676, 0.02372606, 0.00544886, 0.03035324, 0.03884234, 
    -0.00250727, 0.0003113609, 0.1217374, 0.1256382, 0.2427084, 0.1369377, 
    0.1107418, 0.109832, 0.1465383, 0.1635984, 0.2239028, 0.1451785, 
    0.2384009, 0.07556941, 0.02615857, 0.1536027, 0.09122191, 0.160172, 
    0.06181492, 0.1099355, 0.1380769, 0.1182828, 0.006916466,
  0.01457996, 0.03075678, 0.0754601, 0.206563, 0.10306, 0.07260577, 
    0.1712498, -0.0002083114, -0.0002865233, 0.03146592, 0.03236831, 
    0.2009256, 0.3885489, 0.2286789, 0.2239032, 0.3031836, 0.4670891, 
    0.3319416, 0.2443014, 0.356489, 0.2367344, 0.1051759, 0.2423239, 
    0.261996, 0.3631781, 0.2827264, 0.2909983, 0.2269254, 0.2657282,
  0.2166201, 0.2033706, 0.158091, 0.1760339, 0.2246345, 0.2445612, 0.3361361, 
    0.3397252, 0.04805935, 0.03637889, 0.02055634, 0.1121665, 0.2762348, 
    0.55738, 0.6501589, 0.4348543, 0.2867221, 0.1810619, 0.240475, 0.5812509, 
    0.101331, 0.1255189, 0.266509, 0.3254184, 0.3102263, 0.4442475, 0.232004, 
    0.1844455, 0.1499084,
  0.1981133, 0.2489005, 0.3909888, 0.4147524, 0.5794004, 0.4536603, 
    0.4809786, 0.5421492, 0.3934398, 0.4753135, 0.3322521, 0.2239428, 
    0.3280348, 0.5126134, 0.4965953, 0.1927669, 0.06718457, 0.03575135, 
    0.2471863, 0.3812688, 0.3048882, 0.2768134, 0.1358108, 0.1629798, 
    0.6144661, 0.2186331, 0.1942635, 0.2171476, 0.1765742,
  0.311615, 0.2242671, 0.3708563, 0.6315427, 0.2837299, 0.2755882, 0.2898821, 
    0.4485556, 0.4220347, 0.234343, 0.1770553, 0.1580915, 0.1598798, 
    0.2785737, 0.2846119, 0.270859, 0.4414003, 0.4230047, 0.2135796, 
    0.310261, 0.2892998, 0.1919674, 0.1653904, 0.0423737, 0.04613018, 
    0.3260303, 0.2587974, 0.1691525, 0.4751717,
  0.1635291, 0.1107985, 0.1415538, 0.101041, 0.2039351, 0.3249015, 0.3583139, 
    0.3134254, 0.4569418, 0.4333557, 0.3927603, 0.2947724, 0.24374, 
    0.2735161, 0.2813461, 0.3234687, 0.3553835, 0.4038275, 0.339898, 
    0.4027952, 0.3738925, 0.3520757, 0.1863622, 0.08185993, 0.07239813, 
    0.05672201, 0.09666497, 0.2124695, 0.2189617,
  0.1733709, 0.1712074, 0.1690439, 0.1668805, 0.164717, 0.1625535, 0.16039, 
    0.1460796, 0.1407217, 0.1353639, 0.130006, 0.1246481, 0.1192903, 
    0.1139324, 0.1087986, 0.1131492, 0.1174997, 0.1218503, 0.1262009, 
    0.1305514, 0.134902, 0.1490037, 0.1521745, 0.1553453, 0.1585161, 
    0.1616869, 0.1648576, 0.1680284, 0.1751017,
  0.0263656, 0.05740754, 0.0641057, 0.2347944, 0.355817, 0.439402, 0.3066126, 
    0.1809052, 0.1559793, 0.06249514, 0.03841605, 0.1192729, 0.2576159, 
    -0.01605273, 0.1577315, 0.09072749, 0.05885402, 0.1803716, 0.2792928, 
    0.2412252, 0.3758957, 0.3076591, 0.1848524, 0.1431892, 0.3753284, 
    0.3492716, 0.1353357, 0.02345916, 0.04336124,
  0.3713533, 0.2732068, 0.2430187, 0.07699187, 0.1884301, 0.3634942, 
    0.1131411, 0.5107672, 0.4067125, 0.3098047, 0.1372536, 0.001886185, 
    0.02696345, 0.1503826, 0.3107078, 0.3828266, 0.352543, 0.4543166, 
    0.5054421, 0.5032915, 0.4379686, 0.4360194, 0.4092015, 0.2989175, 
    0.3973432, 0.3728839, 0.4216797, 0.4375208, 0.3892049,
  0.4289586, 0.3880864, 0.3313937, 0.3727998, 0.4191216, 0.3650913, 
    0.4749057, 0.5227812, 0.5506578, 0.4942054, 0.4287, 0.4860889, 0.4986446, 
    0.4884827, 0.4673291, 0.4177908, 0.4104175, 0.4839335, 0.4214172, 
    0.3912836, 0.3319267, 0.3331904, 0.3104183, 0.3856353, 0.4117851, 
    0.4756091, 0.4769213, 0.3897715, 0.4520651,
  0.4173492, 0.4422399, 0.415144, 0.3587652, 0.2995733, 0.403339, 0.3724199, 
    0.380621, 0.3998538, 0.4439098, 0.416819, 0.5571138, 0.4840381, 
    0.3461853, 0.3695385, 0.4008139, 0.402767, 0.5537483, 0.4297772, 
    0.3901978, 0.2681371, 0.2439184, 0.2237918, 0.2162228, 0.01046661, 
    0.1317288, 0.2862993, 0.3603695, 0.364363,
  0.2522174, 0.3239152, 0.2739986, 0.2752903, 0.2225118, 0.2006728, 0.161104, 
    0.2287149, 0.352035, 0.358858, 0.4179864, 0.3092605, 0.09915393, 
    0.1354948, 0.2114247, 0.3033196, 0.2971094, 0.3185558, 0.3804938, 
    0.2675511, 0.2460256, 0.2266955, 0.1983351, 0.02901115, 0.0243869, 
    0.1626168, 0.1918306, 0.2372127, 0.2469044,
  0.1877579, 0.1097875, 0.03976569, 0.1130452, 0.1555631, 0.1414129, 
    0.07187166, 0.1469864, 0.2226675, 0.03282486, 0.006102762, 1.377763e-06, 
    -0.001882635, 0.1128452, 0.1182309, 0.08933534, 0.2183808, 0.2523288, 
    0.1459933, 0.1137828, 0.08133363, 0.1969011, 0.3431413, 0.0003713771, 
    0.02921935, 0.147495, 0.1213073, 0.0950224, 0.1380433,
  0.2635872, 0.02659939, 0.01881583, 0.07371192, 0.05496665, 0.05143484, 
    0.05813677, 0.09736925, 0.1173668, 0.08932061, 0.01854469, 0.002245458, 
    0.05539412, 0.1443831, 0.1317958, 0.07462435, 0.0477554, 0.07514282, 
    0.04432599, 0.04395167, 0.04976218, 0.1236299, 0.3106748, 0.01434324, 
    0.07616968, 0.03147433, 0.04282676, 0.0700334, 0.09041667,
  0.1192938, 0.03067382, 0.04051395, 0.06178394, 0.03475263, 0.06188389, 
    0.08335317, 0.06649017, 0.06162635, 0.03820005, 0.06624524, 0.0355386, 
    0.05672769, 0.0966104, 0.06682882, 0.06841775, 0.06528115, 0.08882624, 
    0.07963283, 0.129518, 0.2020603, 0.1733466, 0.1339341, 0.05903261, 
    0.04778686, 0.007159375, 0.08554039, 0.1434142, 0.07979729,
  0.008408124, 0.005067637, 0.0001594075, 0.0002047239, 0.08763878, 
    0.07945023, 0.06272972, 0.0499317, 0.1132007, 0.1658273, 0.05529021, 
    0.06110092, 0.05537481, 0.07373959, 0.1271833, 0.07011516, 0.03322782, 
    0.02543564, 0.05363498, 0.03495794, 0.0697059, 0.06358698, 0.0664456, 
    0.02819455, 0.05306882, 0.04557674, 0.04393374, 0.104734, 0.03583824,
  -4.712138e-08, 1.659814e-09, 6.002077e-10, -0.00147887, 0.13452, 0.1189989, 
    0.01148809, 0.1032383, 0.02178105, 0.1378828, 0.1383039, 0.06239417, 
    0.05954507, 0.07464572, 0.09601494, 0.1095819, 0.09634095, 0.05395738, 
    0.05739323, 0.0616553, 0.05295033, 0.05616778, 0.2575766, 0.1520417, 
    0.06069321, 0.06055001, 0.101356, -0.0001590596, 8.691046e-06,
  5.341283e-08, 2.172595e-08, 1.073939e-09, 0.001351464, -2.987997e-08, 
    0.029743, -6.109063e-07, 0.01335059, 0.004358283, 0.2587926, 0.12964, 
    0.1817617, 0.08786958, 0.1331788, 0.1523874, 0.09635703, 0.2226795, 
    0.1312936, 0.1507147, 0.2344833, 0.01437489, 0.2424206, 0.05224082, 
    0.02611799, 0.01933094, 0.0274889, 0.007042442, 0.006267131, 3.499755e-07,
  -9.951505e-05, 0.003771096, 0.009274852, 0.004358581, 0.02920652, 
    0.02823096, -0.002639259, -3.782358e-06, 0.0934706, 0.1164554, 0.1752902, 
    0.07711779, 0.08322208, 0.07929981, 0.1398102, 0.1113432, 0.1352676, 
    0.1473304, 0.1575677, 0.1226097, 0.03674248, 0.196123, 0.08141244, 
    0.1877435, 0.1251895, 0.1821615, 0.07648539, 0.06558724, 0.003538969,
  0.02397095, 0.04929829, 0.08117962, 0.2105122, 0.0496008, 0.03583232, 
    0.163693, -0.0001694353, -0.0003112935, 0.0244493, 0.03336279, 0.1268512, 
    0.3241339, 0.1931097, 0.1789279, 0.2555786, 0.3993641, 0.2788896, 
    0.1944437, 0.3756956, 0.2335989, 0.1652503, 0.2501124, 0.2703638, 
    0.3011393, 0.2563506, 0.234236, 0.2417135, 0.252654,
  0.2206963, 0.2447495, 0.1636048, 0.2066888, 0.4103472, 0.3456003, 
    0.2918677, 0.3420525, 0.0448939, 0.03397222, 0.0227536, 0.1241595, 
    0.2134292, 0.5231484, 0.6769792, 0.3819951, 0.1808885, 0.08931638, 
    0.1956598, 0.6341348, 0.09094151, 0.1745875, 0.3027222, 0.3343578, 
    0.3072511, 0.3394126, 0.1701257, 0.1577319, 0.1381008,
  0.1637258, 0.2843258, 0.5286496, 0.5619869, 0.7217339, 0.4620514, 
    0.4966861, 0.6074944, 0.439003, 0.4893242, 0.3390438, 0.2511368, 
    0.3454682, 0.4867338, 0.3960177, 0.1555074, 0.09031154, 0.0560015, 
    0.2665798, 0.3846748, 0.3198008, 0.2703674, 0.1409491, 0.1640145, 
    0.8085588, 0.1447177, 0.1282873, 0.1633725, 0.1414363,
  0.2286981, 0.1634386, 0.3500775, 0.5630028, 0.2884406, 0.2844566, 
    0.3111805, 0.4596296, 0.4313796, 0.2788841, 0.2328075, 0.143337, 
    0.1575879, 0.306726, 0.2937075, 0.2736753, 0.52307, 0.4481319, 0.2599095, 
    0.3769855, 0.2952879, 0.2490596, 0.1830909, 0.04519884, 0.05189252, 
    0.3042098, 0.2455338, 0.1548925, 0.4584728,
  0.1518966, 0.08926239, 0.1056526, 0.08025394, 0.1958876, 0.359235, 
    0.3786679, 0.3373567, 0.4829276, 0.4412638, 0.4225439, 0.3204004, 
    0.2824114, 0.3121521, 0.3212235, 0.3607985, 0.3653627, 0.4380343, 
    0.4032479, 0.4399588, 0.4038422, 0.3524912, 0.2021849, 0.05990824, 
    0.07251283, 0.07212098, 0.09697191, 0.2298704, 0.2058329,
  0.2691303, 0.2681251, 0.26712, 0.2661148, 0.2651097, 0.2641045, 0.2630994, 
    0.245565, 0.2381619, 0.2307587, 0.2233555, 0.2159524, 0.2085492, 
    0.201146, 0.1862348, 0.1908867, 0.1955385, 0.2001904, 0.2048423, 
    0.2094942, 0.2141461, 0.2515167, 0.2552732, 0.2590296, 0.262786, 
    0.2665425, 0.2702989, 0.2740553, 0.2699344,
  0.02007959, 0.0535381, 0.07391515, 0.2583517, 0.4093121, 0.4412522, 
    0.3421923, 0.2176127, 0.1604077, 0.1034873, 0.05895055, 0.1066815, 
    0.2441437, -0.01523317, 0.16162, 0.1202076, 0.1161615, 0.1563628, 
    0.2010145, 0.2264544, 0.3957177, 0.2929453, 0.1813108, 0.1646704, 
    0.2435777, 0.2770143, 0.08947675, 0.009287104, 0.03809659,
  0.3264042, 0.1971909, 0.1886469, 0.02831101, 0.1293545, 0.3504365, 
    0.07033964, 0.4129967, 0.3808688, 0.3070814, 0.1318219, 0.0002589936, 
    0.03773026, 0.06165334, 0.2667477, 0.3898168, 0.3665466, 0.4284451, 
    0.5173414, 0.3487488, 0.4096923, 0.3328219, 0.3039679, 0.2911385, 
    0.3787534, 0.284645, 0.3266364, 0.3255671, 0.3071812,
  0.3766286, 0.3762782, 0.2962056, 0.3710331, 0.3823107, 0.3084033, 
    0.4560196, 0.5132326, 0.5884557, 0.4818516, 0.4628436, 0.4882224, 
    0.5410864, 0.4856303, 0.4200757, 0.4230677, 0.4078053, 0.4938234, 
    0.4144881, 0.3442631, 0.2598093, 0.3083607, 0.2790661, 0.3355077, 
    0.3940798, 0.4796662, 0.4662478, 0.3946703, 0.4503327,
  0.411968, 0.4293577, 0.4489718, 0.4132476, 0.3647097, 0.3747029, 0.3951281, 
    0.3239296, 0.319236, 0.3578898, 0.3034971, 0.4300652, 0.392128, 
    0.3196624, 0.3114938, 0.38533, 0.3771491, 0.5051622, 0.4161128, 
    0.3592626, 0.2337576, 0.2312077, 0.2022758, 0.2047154, 0.008955478, 
    0.1380709, 0.3293702, 0.3748132, 0.3915139,
  0.2338093, 0.3027816, 0.2519284, 0.2400976, 0.1907146, 0.2693407, 
    0.1808309, 0.1828719, 0.2783183, 0.2875194, 0.2477147, 0.1498242, 
    0.04910612, 0.1734684, 0.2463429, 0.2805304, 0.2754392, 0.2682729, 
    0.3591729, 0.1716393, 0.2004493, 0.175273, 0.1544869, 0.03422789, 
    0.04722885, 0.19623, 0.1684518, 0.2192034, 0.2110165,
  0.1299886, 0.1564142, 0.03164613, 0.0613187, 0.121047, 0.1362613, 
    0.04203749, 0.05135623, 0.1470928, 0.02157029, 0.004316114, 1.380389e-06, 
    -0.001744878, 0.09027307, 0.09226469, 0.09466702, 0.2287565, 0.2426716, 
    0.2091468, 0.08433516, 0.03231203, 0.05171933, 0.168837, 0.002507858, 
    0.04109756, 0.1379848, 0.0880513, 0.06907136, 0.06732647,
  0.1012937, 0.0470597, 0.01080496, 0.04629107, 0.03124241, 0.01943086, 
    0.04511674, 0.05685487, 0.05762049, 0.06186672, 0.009942862, 
    0.0007843559, 0.1109268, 0.03667679, 0.04022066, 0.05384035, 0.07342218, 
    0.05578817, 0.02884895, 0.008698775, 0.0111503, 0.04999834, 0.1699332, 
    0.4013481, 0.0594541, 0.02959151, 0.01469033, 0.01282275, 0.02656567,
  0.3599645, 0.1922603, 0.02866067, 0.04797402, 0.04964485, 0.0576709, 
    0.04711147, 0.02396375, 0.03403939, 0.04040385, 0.04956067, 0.1039106, 
    0.03867486, 0.02707404, 0.03058399, 0.02068113, 0.02159179, 0.02232165, 
    0.02484211, 0.03445739, 0.04786092, 0.09514543, 0.1340069, 0.03987583, 
    0.03555987, 0.002722357, 0.01812572, 0.02919542, 0.1150477,
  0.06606163, 0.002339833, 9.126016e-05, 0.000106776, 0.06127714, 0.07051638, 
    0.03436752, 0.02865172, 0.06856246, 0.1229221, 0.03038602, 0.1572297, 
    0.02562617, 0.03556998, 0.02467651, 0.04661319, 0.05446763, 0.03831717, 
    0.04497781, 0.03862675, 0.07410619, 0.1928654, 0.07900217, 0.01228362, 
    0.02447001, 0.0193788, 0.02594559, 0.05973894, 0.1642335,
  -1.748414e-08, 1.251455e-09, 3.518204e-10, 0.0004179799, 0.1471542, 
    0.0384883, 0.005321105, 0.0451289, 0.02114718, 0.08975018, 0.1444369, 
    0.0397227, 0.02254297, 0.05710714, 0.03856289, 0.05343071, 0.05033327, 
    0.03591929, 0.03407689, 0.02834465, 0.02708905, 0.0222473, 0.4268927, 
    0.1766146, 0.02725208, 0.02350201, 0.02532728, 0.006227265, -3.595859e-07,
  5.044441e-08, 1.536551e-08, 4.989141e-10, 0.0004426177, -1.390178e-10, 
    0.01374635, 1.048527e-07, 0.01987545, 0.004523691, 0.2697497, 0.0749531, 
    0.1104885, 0.06130865, 0.07417785, 0.06775576, 0.04748628, 0.1638052, 
    0.1195416, 0.1121681, 0.1738258, 0.002293488, 0.2118899, 0.009247915, 
    0.01611164, 0.005361522, 0.009870097, 0.001157921, 0.001603262, 
    2.917694e-07,
  -3.250931e-05, 0.01376726, 0.003268725, 0.00300887, 0.02443126, 0.02469888, 
    -0.00258886, -6.548336e-05, 0.0691465, 0.1281008, 0.1392034, 0.05693867, 
    0.0600525, 0.06871493, 0.1339144, 0.09445758, 0.09575687, 0.1145692, 
    0.1164477, 0.1349187, 0.03742777, 0.2314599, 0.06241804, 0.1093912, 
    0.0869453, 0.0952292, 0.02332543, 0.02487025, 0.002362319,
  0.02453113, 0.01321747, 0.0307399, 0.2060393, 0.01232341, 0.04975842, 
    0.1574904, -0.0001049327, -0.0002312004, 0.02088238, 0.05179368, 
    0.08875571, 0.2641296, 0.172622, 0.1661642, 0.1981886, 0.3357479, 
    0.2367148, 0.1785353, 0.4023929, 0.211092, 0.2087088, 0.2374218, 
    0.289188, 0.313545, 0.2113967, 0.1953002, 0.1833728, 0.2325805,
  0.2042028, 0.2352845, 0.1852711, 0.3446139, 0.4380237, 0.430871, 0.2624515, 
    0.3377691, 0.0360527, 0.02370032, 0.01369347, 0.1284678, 0.177407, 
    0.4968714, 0.5244744, 0.219053, 0.1285428, 0.04563241, 0.1768688, 
    0.6120599, 0.1034406, 0.1967697, 0.2965221, 0.3639761, 0.335732, 
    0.2494295, 0.1325291, 0.1480847, 0.1510849,
  0.1378112, 0.321956, 0.565405, 0.6909503, 0.7179842, 0.4372166, 0.4918676, 
    0.5830772, 0.4275239, 0.4742397, 0.3669191, 0.2831585, 0.3449602, 
    0.4845292, 0.2325907, 0.0951452, 0.1226115, 0.0463446, 0.3265247, 
    0.4114835, 0.3530976, 0.280131, 0.1586346, 0.1356145, 0.7846836, 
    0.09505767, 0.0696303, 0.1325332, 0.1110674,
  0.1611399, 0.105587, 0.3333258, 0.4614568, 0.2730687, 0.3202741, 0.3595333, 
    0.5307865, 0.4319043, 0.3119429, 0.2616765, 0.1491911, 0.1560612, 
    0.3166482, 0.2922358, 0.227303, 0.6189213, 0.4872169, 0.2919689, 
    0.454586, 0.2805835, 0.3266876, 0.2133939, 0.03725918, 0.06097921, 
    0.2867875, 0.2388347, 0.1721538, 0.374275,
  0.1636235, 0.1226316, 0.1244284, 0.07402251, 0.2124058, 0.3591227, 
    0.3944237, 0.3911984, 0.4908834, 0.462757, 0.3991872, 0.3861812, 
    0.324011, 0.3585285, 0.353085, 0.4068281, 0.389205, 0.4822732, 0.4390602, 
    0.4690733, 0.4264897, 0.3579494, 0.230499, 0.04063062, 0.06917749, 
    0.08799205, 0.08150727, 0.2583133, 0.2130434,
  0.3860271, 0.3870821, 0.3881371, 0.3891921, 0.3902471, 0.3913021, 
    0.3923571, 0.39097, 0.3807516, 0.3705331, 0.3603147, 0.3500963, 
    0.3398778, 0.3296594, 0.313884, 0.3176225, 0.3213611, 0.3250996, 
    0.3288382, 0.3325768, 0.3363153, 0.3463276, 0.3517525, 0.3571774, 
    0.3626022, 0.3680271, 0.373452, 0.3788768, 0.3851831,
  0.02894714, 0.0717443, 0.1106439, 0.2912119, 0.4655885, 0.4647427, 
    0.3727922, 0.2758813, 0.1702063, 0.1802866, 0.08545409, 0.09144655, 
    0.2363545, -0.00864206, 0.1702989, 0.1630177, 0.2778884, 0.1760699, 
    0.1072572, 0.228809, 0.3466562, 0.323308, 0.1843025, 0.1856431, 
    0.2620711, 0.1973658, 0.06231547, -0.002966183, 0.02624088,
  0.2089111, 0.1276484, 0.1393494, 0.01543579, 0.06842687, 0.3134069, 
    0.04937008, 0.2929341, 0.3282051, 0.2808698, 0.1165059, 0.001596828, 
    0.03948412, 0.03531622, 0.257746, 0.4155245, 0.3859624, 0.3911091, 
    0.4981422, 0.2822312, 0.3792706, 0.2735065, 0.2339446, 0.3004798, 
    0.3748804, 0.2328093, 0.2586116, 0.2432376, 0.2480582,
  0.3700474, 0.3401752, 0.2403591, 0.329982, 0.3169664, 0.2486878, 0.4454968, 
    0.4940414, 0.5845333, 0.4492221, 0.4553233, 0.4831367, 0.5372202, 
    0.4631938, 0.4016698, 0.3893759, 0.4010673, 0.4664224, 0.3814125, 
    0.2842026, 0.2188087, 0.2643496, 0.2560411, 0.3199541, 0.3432373, 
    0.4922071, 0.4892907, 0.393406, 0.404624,
  0.4397204, 0.4218185, 0.4729162, 0.4357835, 0.3774788, 0.3719829, 
    0.3688526, 0.267917, 0.295481, 0.319285, 0.2113912, 0.2779306, 0.3083382, 
    0.2474393, 0.245649, 0.3906616, 0.3656785, 0.4075478, 0.3688551, 
    0.3067972, 0.1900011, 0.2119723, 0.1929136, 0.184669, 0.01053474, 
    0.1988862, 0.3375145, 0.4332319, 0.4190056,
  0.1561023, 0.2268516, 0.1554374, 0.2130885, 0.2074243, 0.2807156, 
    0.1323449, 0.1356643, 0.188955, 0.208073, 0.1148882, 0.08282016, 
    0.0284736, 0.1524115, 0.2448474, 0.2601286, 0.2385838, 0.1955411, 
    0.2376457, 0.1885125, 0.1586432, 0.1278337, 0.1209682, 0.05314283, 
    0.04930862, 0.2116597, 0.1767618, 0.1526143, 0.1316836,
  0.05012555, 0.08032602, 0.01468435, 0.02567388, 0.1659225, 0.1198393, 
    0.01940587, 0.02293839, 0.08810116, 0.01027303, 0.002119492, 
    -1.509676e-08, -0.001033264, 0.06316321, 0.05708137, 0.04839575, 
    0.2107306, 0.2394828, 0.1408882, 0.06126786, 0.02452771, 0.01471187, 
    0.06548756, 0.01702619, 0.04857431, 0.1191439, 0.02411807, 0.02009723, 
    0.03441766,
  0.02512811, 0.1055441, 0.007169622, 0.02218068, 0.01461773, 0.007357465, 
    0.0099363, 0.03845066, 0.03857477, 0.02959241, 0.008368385, 0.0003045994, 
    0.04146813, 0.00846504, 0.01600723, 0.01925795, 0.01782643, 0.01959476, 
    0.005004682, 0.0008080779, 0.0003748698, 0.009615855, 0.04845425, 
    0.2333491, 0.04448353, 0.02955325, 0.001615688, 0.002081051, 0.004422429,
  0.08449968, 0.1197866, 0.01875057, 0.03541958, 0.01510654, 0.01100007, 
    0.01899058, 0.004076593, 0.01860272, 0.0127669, 0.0318507, 0.01467722, 
    0.02432396, 0.008274506, 0.01005408, 0.002612001, 0.0029436, 0.006214553, 
    0.003692396, 0.007258656, 0.01186101, 0.02167584, 0.02298653, 0.03150575, 
    0.02950438, 0.0009128833, -9.769316e-05, 0.006148781, 0.01536666,
  0.00835325, 0.001204009, 0.0001130651, -9.986923e-05, 0.02919497, 
    0.01025377, 0.009138851, 0.008548735, 0.0419343, 0.08466678, 0.01992527, 
    0.04815512, 0.004303341, 0.01027752, 0.004622989, 0.006751704, 
    0.01890359, 0.03416388, 0.04127796, 0.02609366, 0.04761433, 0.1795141, 
    0.1480793, 0.005770374, 0.01406957, 0.003926202, 0.01101019, 0.008363026, 
    0.03046935,
  -4.115511e-09, 1.09377e-09, 2.437328e-10, 0.0007861504, 0.1073497, 
    0.009762607, -0.0003365002, 0.008035549, 0.005184536, 0.03311205, 
    0.08954202, 0.01881395, 0.005294825, 0.01902929, 0.007972165, 0.01831753, 
    0.02788658, 0.01477025, 0.01215045, 0.007385393, 0.01097587, 0.002969072, 
    0.4097067, 0.1589186, 0.006687575, 0.006581375, 0.005828254, 
    0.0008236998, -4.488251e-06,
  4.777235e-08, 1.241669e-08, 2.636883e-10, 0.0002024864, 3.185285e-09, 
    0.002886973, 7.432608e-08, 0.01242997, 0.002256261, 0.2443929, 
    0.04287109, 0.05361224, 0.01330791, 0.02070587, 0.03034037, 0.0121374, 
    0.1028913, 0.04762399, 0.03523538, 0.08084777, 0.0007359875, 0.1787653, 
    0.00197995, 0.003176764, 0.002077722, 0.006090745, 0.0002684049, 
    0.0006254052, 2.609337e-07,
  -1.26805e-05, 0.01493523, 0.0005344173, 0.001528626, 0.01983771, 
    0.02189853, -0.00241107, -3.239793e-05, 0.04612251, 0.1351179, 0.1142685, 
    0.03834578, 0.04244952, 0.05844881, 0.1310955, 0.08799896, 0.08870395, 
    0.09902689, 0.09745134, 0.07842463, 0.03169775, 0.2358901, 0.05656494, 
    0.07499912, 0.03318306, 0.03489707, 0.01464777, 0.005804439, 0.002812231,
  0.01974519, 0.004324169, 0.01879599, 0.1993368, 0.00425168, 0.08721265, 
    0.1558655, -5.871857e-05, -0.0001824105, 0.01601399, 0.05271842, 
    0.06353217, 0.2161551, 0.1672192, 0.1447504, 0.1678147, 0.2773739, 
    0.2178701, 0.1608495, 0.4100241, 0.2007288, 0.1728369, 0.2478689, 
    0.2638635, 0.248792, 0.1706231, 0.1620214, 0.1194324, 0.1716623,
  0.1644798, 0.1522877, 0.2348144, 0.4958695, 0.4210683, 0.4703943, 
    0.2082877, 0.3014919, 0.02854757, 0.02079936, 0.007882424, 0.1196646, 
    0.1772406, 0.4949447, 0.4060798, 0.1199321, 0.06623099, 0.02976773, 
    0.1509232, 0.5759872, 0.1207913, 0.2167028, 0.2703215, 0.3977374, 
    0.3094192, 0.1981778, 0.1069085, 0.1291069, 0.1426005,
  0.1153993, 0.3536704, 0.5505439, 0.6906621, 0.6476927, 0.3792045, 
    0.5077519, 0.5919497, 0.4392522, 0.4696673, 0.3905207, 0.3404216, 
    0.3444954, 0.4675685, 0.1350016, 0.08961027, 0.1663299, 0.03770606, 
    0.3736171, 0.4413195, 0.4366857, 0.2766536, 0.1829919, 0.1237039, 
    0.7489128, 0.05952498, 0.04214577, 0.09370554, 0.08378502,
  0.1242563, 0.07084392, 0.3095199, 0.3724919, 0.3055858, 0.3704428, 
    0.4610389, 0.5918523, 0.3540852, 0.3273526, 0.3476776, 0.1557937, 
    0.162803, 0.3510434, 0.2795854, 0.1990981, 0.6535514, 0.4994703, 
    0.3177451, 0.5055211, 0.2167624, 0.3486908, 0.2686674, 0.04639284, 
    0.06650186, 0.2674594, 0.2386149, 0.1331453, 0.3068899,
  0.2061519, 0.2300244, 0.1855133, 0.09299625, 0.2233951, 0.3663911, 
    0.4603611, 0.4386153, 0.5129737, 0.4977932, 0.4224516, 0.4674024, 
    0.3860972, 0.4254729, 0.4297034, 0.47822, 0.4739827, 0.5379586, 
    0.4842171, 0.529183, 0.4612824, 0.3503008, 0.2774226, 0.05170401, 
    0.0907907, 0.1133153, 0.08608671, 0.2792775, 0.2439938,
  0.4845036, 0.4915984, 0.4986932, 0.505788, 0.5128828, 0.5199776, 0.5270724, 
    0.5164254, 0.5089211, 0.5014169, 0.4939126, 0.4864084, 0.4789041, 
    0.4713998, 0.4582838, 0.4561226, 0.4539614, 0.4518002, 0.449639, 
    0.4474778, 0.4453166, 0.4418329, 0.4444036, 0.4469743, 0.4495449, 
    0.4521156, 0.4546863, 0.4572569, 0.4788278,
  0.03050267, 0.08193073, 0.1442336, 0.3062599, 0.4951059, 0.4702927, 
    0.4147032, 0.3224814, 0.1556811, 0.2123251, 0.09843836, 0.04812905, 
    0.180792, -0.002826135, 0.2110785, 0.2162085, 0.4731669, 0.2256528, 
    0.08095106, 0.1856851, 0.3165065, 0.3237554, 0.1765952, 0.143805, 
    0.2687928, 0.2003759, 0.04630269, -0.004018121, 0.025371,
  0.1291817, 0.0654426, 0.07946838, 0.008285855, 0.03642352, 0.2725462, 
    0.03272865, 0.1898777, 0.2612412, 0.2259317, 0.0772041, 0.001297424, 
    0.02378581, 0.01801446, 0.2416617, 0.3911566, 0.3505315, 0.3406482, 
    0.4136806, 0.2736267, 0.3480904, 0.2740436, 0.2304755, 0.261066, 
    0.3195689, 0.208322, 0.2393045, 0.1844056, 0.2070504,
  0.3202733, 0.2867143, 0.1912733, 0.2679227, 0.2739966, 0.1945567, 
    0.4042854, 0.4151135, 0.5288936, 0.4283991, 0.4024478, 0.4650223, 
    0.5138228, 0.4325824, 0.3694817, 0.3815684, 0.4001583, 0.431887, 
    0.3462305, 0.2360593, 0.2041913, 0.2026938, 0.2074355, 0.266983, 
    0.2976235, 0.4663062, 0.47364, 0.3536146, 0.3525512,
  0.425098, 0.3913921, 0.4314358, 0.3726453, 0.3612038, 0.3463924, 0.3381361, 
    0.2122793, 0.2615395, 0.2908219, 0.181652, 0.2021892, 0.2462442, 
    0.2187778, 0.231275, 0.3554694, 0.3147044, 0.2980869, 0.3182169, 
    0.2545772, 0.1465203, 0.159973, 0.1732364, 0.1439674, 0.01998211, 
    0.2152782, 0.3084377, 0.4240928, 0.4377885,
  0.1160726, 0.1398054, 0.07971539, 0.1650001, 0.1705828, 0.2454104, 
    0.09107973, 0.09206312, 0.1501257, 0.1656542, 0.05895539, 0.04932327, 
    0.02900118, 0.1030786, 0.2277191, 0.22577, 0.1674222, 0.1592553, 0.16933, 
    0.15715, 0.1262705, 0.1014581, 0.07578506, 0.06852797, 0.04182056, 
    0.1697495, 0.1707046, 0.1051242, 0.08901558,
  0.02449811, 0.02930979, 0.00764692, 0.01023385, 0.1145675, 0.09510018, 
    0.0047349, 0.005805819, 0.03189047, 0.01195634, 0.001744286, 
    -1.179057e-08, 0.002280457, 0.04960425, 0.01592016, 0.01852174, 
    0.1841225, 0.2157876, 0.09718301, 0.03329193, 0.004434668, 0.005588389, 
    0.02355525, 0.01296251, 0.04043886, 0.07635157, 0.006646743, 0.002865546, 
    0.0181584,
  0.007688835, 0.1420855, 0.006339001, 0.008039575, 0.004697963, 0.002471614, 
    0.002820924, 0.02408475, 0.01056879, 0.008985663, 0.006892081, 
    0.0001177488, 0.01233236, 0.003588919, 0.00841273, 0.004973006, 
    0.002105531, 0.00901335, 0.0004523468, 0.0001979791, 6.034313e-05, 
    0.002679508, 0.01696863, 0.07882538, 0.03273292, 0.02827912, 
    0.0002739893, 0.0006607436, 0.001336721,
  0.03101439, 0.03689627, 0.0162865, 0.03193196, 0.002662739, 0.001451667, 
    0.01099308, 0.0007020906, 0.003869753, 0.000588687, 0.01474277, 
    0.004364657, 0.005053787, 0.0007382542, 0.005395785, 0.0004777555, 
    0.0004473061, 0.001593763, 0.001149019, 0.002210704, 0.004364405, 
    0.007574723, 0.008007474, 0.02905372, 0.02708211, 0.0004925531, 
    -0.0007646474, 0.002770826, 0.004160393,
  0.001625179, 0.0008654018, 8.021263e-05, -0.0001226374, 0.01187946, 
    0.002423661, 0.0009822547, 0.0009915301, 0.02614966, 0.08614914, 
    0.00166063, 0.008324379, 0.0004740999, 0.005851462, 0.001719688, 
    0.001271917, 0.001831158, 0.00608569, 0.01608632, 0.003872921, 
    0.01210765, 0.03895869, 0.03667891, 0.002695287, 0.007567217, 
    0.0007873236, 0.002289149, 0.002084854, 0.006782023,
  -9.452147e-09, 1.042625e-09, 1.838758e-10, -0.0001594375, 0.05583806, 
    0.003239911, -0.001845835, 0.002638106, 0.0007284108, 0.006813318, 
    0.04126031, 0.00648163, 0.001132264, 0.005991801, 0.00104364, 
    0.006756413, 0.0134053, 0.002709467, 0.001381467, 0.001061554, 
    0.003878888, 0.0004457627, 0.2978115, 0.1378578, 0.001944493, 
    0.002313232, 0.002643712, 0.0002751053, -3.198281e-05,
  4.507554e-08, 1.095261e-08, 2.555605e-10, 0.0001140829, 4.258131e-09, 
    0.0007313091, 5.302245e-08, 0.006290909, 0.001540615, 0.1682732, 
    0.01751452, 0.02465823, 0.005338082, 0.007831132, 0.01368213, 
    0.003366881, 0.05937615, 0.01469422, 0.01289588, 0.03576485, 
    0.0003707941, 0.13128, 0.0007100551, -0.0008487625, 0.0008883303, 
    0.003632467, 0.0003158081, 0.0003173668, 2.362822e-07,
  -1.648561e-05, 0.01245895, 0.0002202584, 0.000626311, 0.01699497, 
    0.0178682, -0.002118445, 0.0001129591, 0.03375974, 0.1128943, 0.0896984, 
    0.02661642, 0.02887704, 0.04159287, 0.103265, 0.06351136, 0.07299056, 
    0.08120093, 0.07952742, 0.0426406, 0.02223708, 0.2065586, 0.05228706, 
    0.05869416, 0.01963774, 0.01923826, 0.01248915, 0.002642173, 0.001871331,
  0.01147103, 0.001388201, 0.01598773, 0.1881257, 0.002216351, 0.07765226, 
    0.1509221, -2.171215e-05, -0.0001421821, 0.009135839, 0.05288602, 
    0.04426243, 0.1682507, 0.1444176, 0.1131394, 0.1409438, 0.2150234, 
    0.1707583, 0.1290425, 0.3964115, 0.1762865, 0.1501766, 0.2275774, 
    0.2637115, 0.1718467, 0.1132743, 0.113095, 0.07666617, 0.133402,
  0.1135132, 0.1023549, 0.1967857, 0.5182311, 0.4322779, 0.3935336, 
    0.1558248, 0.2512483, 0.03137355, 0.01675042, 0.004210467, 0.1162787, 
    0.1979815, 0.4391426, 0.3289435, 0.07413353, 0.04265014, 0.02123351, 
    0.1239349, 0.5402844, 0.1201569, 0.2075598, 0.240874, 0.3778263, 
    0.2698635, 0.1631691, 0.08721896, 0.1122501, 0.1016156,
  0.08636158, 0.4209322, 0.5500534, 0.612609, 0.5810673, 0.3841392, 
    0.4908966, 0.5607831, 0.4436947, 0.4550852, 0.3995676, 0.3736235, 
    0.3168263, 0.438223, 0.08057966, 0.1311407, 0.2104241, 0.0618384, 
    0.3704522, 0.4248888, 0.4466359, 0.2182003, 0.2088641, 0.1262642, 
    0.7223818, 0.03938072, 0.03030152, 0.06889516, 0.05867167,
  0.09835126, 0.04883855, 0.3174496, 0.2611145, 0.4496844, 0.4532044, 
    0.5637561, 0.5319455, 0.2856528, 0.3505586, 0.4118969, 0.1480451, 
    0.2050919, 0.3880732, 0.2648686, 0.2225999, 0.6262518, 0.4417142, 
    0.3269815, 0.5167041, 0.1793861, 0.4156992, 0.281198, 0.09499078, 
    0.07688174, 0.2508148, 0.2457834, 0.1086071, 0.2445874,
  0.2783522, 0.3712397, 0.2748137, 0.1654986, 0.2010873, 0.404709, 0.5167137, 
    0.5194448, 0.5526852, 0.566259, 0.5739563, 0.5696846, 0.5186651, 
    0.5442948, 0.5208475, 0.5376175, 0.5658721, 0.5968199, 0.5831921, 
    0.5820337, 0.5740334, 0.343907, 0.2789445, 0.1008754, 0.1197428, 
    0.1390342, 0.06823798, 0.3386467, 0.3436725,
  0.5371985, 0.5458538, 0.554509, 0.5631642, 0.5718195, 0.5804747, 0.58913, 
    0.5324047, 0.5322875, 0.5321704, 0.5320532, 0.531936, 0.5318189, 
    0.5317017, 0.5992005, 0.5927645, 0.5863284, 0.5798925, 0.5734564, 
    0.5670204, 0.5605844, 0.5415578, 0.5394558, 0.5373537, 0.5352516, 
    0.5331495, 0.5310475, 0.5289454, 0.5302743,
  0.04646148, 0.09572122, 0.1376526, 0.3691686, 0.5533315, 0.4498415, 
    0.4379828, 0.3996558, 0.1394517, 0.170126, 0.09161936, 0.02619152, 
    0.1136436, -0.0006715442, 0.1919207, 0.4007028, 0.4028789, 0.2322969, 
    0.05428539, 0.2320057, 0.2894785, 0.3297255, 0.1483977, 0.09272601, 
    0.2278516, 0.1819995, 0.05621586, -0.004159555, 0.02834377,
  0.09147774, 0.03829591, 0.04762562, 0.006133959, 0.02432139, 0.2261533, 
    0.02279793, 0.1074752, 0.1922572, 0.1741598, 0.0451789, 0.0009129225, 
    0.01564956, 0.007137131, 0.2180188, 0.3442342, 0.2867129, 0.2823976, 
    0.3474955, 0.2455337, 0.3305204, 0.2661241, 0.2446344, 0.1951361, 
    0.2363157, 0.1875317, 0.1688565, 0.1166205, 0.1551773,
  0.2460608, 0.2359106, 0.1608813, 0.2117282, 0.22216, 0.1487138, 0.3204664, 
    0.3349954, 0.4602358, 0.3891744, 0.3409862, 0.4061488, 0.4744189, 
    0.3743671, 0.3294896, 0.3305983, 0.3529122, 0.3676513, 0.3019338, 
    0.1884892, 0.1813321, 0.1561816, 0.1362553, 0.2126868, 0.2608478, 
    0.4372939, 0.4411238, 0.2970985, 0.2947073,
  0.3403804, 0.3035694, 0.3504062, 0.2942566, 0.2869754, 0.2721319, 
    0.2661874, 0.1649482, 0.2019549, 0.2411461, 0.1451331, 0.1494568, 
    0.193289, 0.16139, 0.2087511, 0.3461888, 0.281181, 0.2349038, 0.2412107, 
    0.1962687, 0.1008908, 0.1058951, 0.1344127, 0.1094715, 0.02433142, 
    0.1854129, 0.2747409, 0.3475223, 0.377124,
  0.08571146, 0.09113087, 0.05382355, 0.1222472, 0.1271591, 0.1936297, 
    0.05091228, 0.06481553, 0.1335895, 0.128325, 0.03582968, 0.02722273, 
    0.02098083, 0.06877427, 0.2031703, 0.1664369, 0.1402012, 0.1420879, 
    0.150384, 0.1092164, 0.08878107, 0.07257827, 0.04127128, 0.07353077, 
    0.04613279, 0.1137313, 0.1305933, 0.07926595, 0.05925677,
  0.01292297, 0.01071222, 0.00443637, 0.003958331, 0.05392139, 0.05641691, 
    0.001504623, 0.0029994, 0.01483534, 0.003138994, 0.000633053, 
    -3.99958e-09, 0.001392332, 0.03557823, 0.004399023, 0.005015187, 
    0.1307058, 0.1985035, 0.07524581, 0.01651108, 0.001308995, 0.003023279, 
    0.01236189, 0.007048975, 0.03085806, 0.03725079, 0.002788683, 
    0.0007811605, 0.006893198,
  0.003583042, 0.1295336, 0.004429101, 0.002951638, 0.0008798641, 
    0.0007459244, 0.0009894697, 0.01197007, 0.005087214, 0.003566635, 
    0.005779177, 6.060295e-05, 0.003996383, 0.001828933, 0.004968175, 
    0.001791138, 0.000645553, 0.002549605, 0.0001231877, 5.479857e-05, 
    2.106667e-05, 0.001147375, 0.00805446, 0.04118105, 0.02359073, 
    0.02652835, 0.0001479437, 0.0003841779, 0.0006896665,
  0.0164092, 0.01396538, 0.01614351, 0.02998704, 0.000740397, 0.000626695, 
    0.0100272, 0.0002260133, 0.001855719, -0.0009657159, 0.006581114, 
    0.002012462, 0.0006821812, 0.0001352327, 0.002347014, 0.0002364344, 
    0.000195737, 0.000838991, 0.0005795142, 0.001176658, 0.002460515, 
    0.003902792, 0.00421993, 0.02717681, 0.02489009, 0.001905683, 
    -0.0003732651, 0.00159842, 0.00214154,
  0.0007334712, 0.001600199, 2.900699e-05, -0.00010039, 0.004589475, 
    0.001031938, 0.000264567, 0.0002746245, 0.0221094, 0.09010758, 
    0.0004210453, 0.003179293, 0.000176485, 0.005053017, 0.0009687252, 
    0.0005098886, 0.0004551234, 0.0006130363, 0.006577104, 0.0005333185, 
    0.006171869, 0.01285505, 0.00876065, 0.00108571, 0.00392265, 
    0.0001902812, 0.0004858319, 0.001150963, 0.003343049,
  -5.453502e-11, 1.025405e-09, 1.481932e-10, 0.001405813, 0.03165452, 
    0.001668569, -0.002332934, 0.001438572, 0.0003177704, 0.002744251, 
    0.01774063, 0.001349928, 0.0004109926, 0.001855021, 0.0004817471, 
    0.00266372, 0.006231675, 0.0007379006, 0.0002106848, 0.0003368515, 
    0.001368202, 0.0002304662, 0.2125882, 0.1153401, 0.0004702357, 
    0.001137013, 0.001495634, 0.0001343151, -0.0001144359,
  4.159961e-08, 1.035161e-08, 2.766573e-10, 7.275087e-05, 4.333744e-09, 
    0.0003427188, 3.914656e-08, 0.00212246, 0.001485969, 0.08556604, 
    0.007544497, 0.01246869, 0.003670797, 0.004109108, 0.006375625, 
    0.001766667, 0.03443222, 0.008113004, 0.006899448, 0.01861189, 
    0.000231986, 0.09358764, 0.0004245196, -0.0009372554, 0.0002044692, 
    0.001386436, 0.0001197138, 0.0001924076, 2.197543e-07,
  -8.909644e-06, 0.007978966, 0.0001368636, 0.0001572835, 0.01390477, 
    0.01277814, -0.001842213, 0.000478307, 0.02484321, 0.08838576, 
    0.05873861, 0.01595591, 0.01674996, 0.01915969, 0.06956536, 0.03170663, 
    0.05148961, 0.06575587, 0.04988107, 0.02363023, 0.01510745, 0.1595664, 
    0.04311616, 0.03072933, 0.01060318, 0.01033712, 0.006839174, 0.001594776, 
    0.002192218,
  0.004452393, 0.0006244704, 0.01835786, 0.1770898, 0.001510591, 0.06295069, 
    0.1442657, -1.177578e-05, -0.0001086964, 0.004564394, 0.04855977, 
    0.0305907, 0.1290227, 0.1240373, 0.08503637, 0.106945, 0.1525597, 
    0.1255215, 0.08650999, 0.3716104, 0.1464444, 0.1278414, 0.1891244, 
    0.2354449, 0.1118613, 0.07674604, 0.06595853, 0.04297077, 0.08930922,
  0.06647541, 0.07829704, 0.179525, 0.4863912, 0.371421, 0.2968476, 
    0.1184198, 0.2146903, 0.03652604, 0.01876175, 0.003403716, 0.115874, 
    0.221073, 0.3555194, 0.2759763, 0.0530079, 0.03189896, 0.01574132, 
    0.1013653, 0.5084322, 0.1036686, 0.1629905, 0.2107759, 0.3719774, 
    0.2149885, 0.1402609, 0.06723499, 0.08085655, 0.06522564,
  0.06631421, 0.4382631, 0.4983663, 0.5200753, 0.5017607, 0.4174601, 
    0.4672956, 0.5120542, 0.4230927, 0.4041054, 0.3934663, 0.3957584, 
    0.2850065, 0.3905911, 0.05099615, 0.1680194, 0.2631857, 0.06353087, 
    0.3240183, 0.4272888, 0.3975172, 0.1756949, 0.2530819, 0.1129784, 
    0.7044449, 0.02924423, 0.02292951, 0.05115999, 0.04285309,
  0.07769049, 0.03068264, 0.3024552, 0.1891724, 0.5549665, 0.4595954, 
    0.6532143, 0.4770318, 0.3127836, 0.4179709, 0.5479196, 0.1647868, 
    0.3585547, 0.3935635, 0.2610861, 0.2471743, 0.5264184, 0.3657858, 
    0.3680483, 0.4861071, 0.2229098, 0.4949398, 0.3013594, 0.1421755, 
    0.08569463, 0.2129932, 0.2628835, 0.08955868, 0.1987479,
  0.4091259, 0.3588395, 0.4420874, 0.2294465, 0.2413753, 0.5005907, 
    0.6058248, 0.5343933, 0.5079973, 0.6174532, 0.6315089, 0.622656, 
    0.5677125, 0.570131, 0.5164552, 0.5725172, 0.5772026, 0.6778426, 
    0.6137011, 0.6355869, 0.6462471, 0.2634324, 0.259639, 0.1640477, 
    0.09498648, 0.1359287, 0.06174482, 0.3423166, 0.4188754,
  0.5117947, 0.5172998, 0.5228049, 0.5283099, 0.533815, 0.5393202, 0.5448253, 
    0.4297071, 0.4375994, 0.4454917, 0.453384, 0.4612762, 0.4691685, 
    0.4770608, 0.6167615, 0.609404, 0.6020465, 0.594689, 0.5873315, 0.579974, 
    0.5726165, 0.5548045, 0.5487646, 0.5427247, 0.5366848, 0.530645, 
    0.5246051, 0.5185652, 0.5073906,
  0.06510687, 0.08072527, 0.1199501, 0.3960444, 0.6094645, 0.3827694, 
    0.3891216, 0.4051474, 0.1534822, 0.08240358, 0.04940511, 0.008655882, 
    0.04442764, 0.0006497232, 0.160923, 0.3678779, 0.3326051, 0.2080527, 
    0.06822816, 0.237987, 0.2787934, 0.2934074, 0.1207107, 0.07161057, 
    0.1832455, 0.1743222, 0.0913734, -0.002720034, 0.02751747,
  0.06499991, 0.02674301, 0.03289826, 0.008063613, 0.01985449, 0.1915389, 
    0.01552176, 0.0659605, 0.1464651, 0.1418815, 0.03681027, 0.001684635, 
    0.01095071, 0.002526207, 0.1807714, 0.2790572, 0.2254624, 0.2289506, 
    0.2844551, 0.2001737, 0.2766007, 0.2237323, 0.2128663, 0.1583294, 
    0.1777339, 0.1519384, 0.1229101, 0.06999011, 0.1060641,
  0.1636906, 0.1852076, 0.1155044, 0.1688117, 0.1762937, 0.1060139, 0.227432, 
    0.2510267, 0.3698659, 0.2941131, 0.2494013, 0.2919133, 0.3884326, 
    0.3003967, 0.2584001, 0.2589627, 0.2847379, 0.3117343, 0.2527535, 
    0.1428358, 0.1282105, 0.1045664, 0.08349755, 0.1560565, 0.2167166, 
    0.3776765, 0.3594206, 0.2298647, 0.2197381,
  0.2409569, 0.2160512, 0.2599841, 0.2216781, 0.2198414, 0.2124566, 
    0.1943773, 0.1226329, 0.1345298, 0.1719522, 0.09758251, 0.0971876, 
    0.136361, 0.09415604, 0.1587657, 0.2960339, 0.2168189, 0.1779543, 
    0.1647511, 0.127888, 0.06495772, 0.07140218, 0.09435076, 0.08543493, 
    0.01996521, 0.1403899, 0.2292201, 0.2668441, 0.2932924,
  0.05735852, 0.06182492, 0.03863354, 0.08111742, 0.09269579, 0.1294726, 
    0.02762495, 0.04468101, 0.1022565, 0.08651614, 0.0229417, 0.01561305, 
    0.01116323, 0.03918685, 0.1744098, 0.0912313, 0.0982964, 0.1181967, 
    0.1257349, 0.07078997, 0.05637938, 0.04342304, 0.01989069, 0.07860538, 
    0.03580702, 0.07218052, 0.08398633, 0.04855385, 0.03397032,
  0.007253266, 0.005452028, 0.003034689, 0.001306318, 0.03106017, 0.03312524, 
    0.0007451772, 0.001980385, 0.008997508, 0.001457964, 0.0002243612, 
    2.112952e-09, -0.000367144, 0.01565249, 0.001687315, 0.0023, 0.07828706, 
    0.1459262, 0.05538193, 0.008866612, 0.0007471177, 0.002002129, 
    0.007966111, 0.002292729, 0.02224662, 0.01127646, 0.001721847, 
    0.0004078645, 0.0022612,
  0.002152827, 0.09040625, 0.001588299, 0.001005775, -0.000638479, 
    0.0002814087, 0.0005197677, 0.004471054, 0.003166538, 0.001853985, 
    0.002630898, 1.347317e-05, 0.001681912, 0.001210553, 0.002482061, 
    0.0008023405, 0.0003891108, 0.0009653817, 6.786521e-05, 2.517372e-05, 
    1.194291e-05, 0.0006413969, 0.004732446, 0.02695033, 0.0169151, 
    0.02085176, 9.710063e-05, 0.0002583001, 0.0004299892,
  0.01068372, 0.007991632, 0.01196054, 0.02745797, 0.0003437938, 
    0.0003919716, 0.006366593, 0.0001272879, 0.0005284081, -0.000684496, 
    0.001818679, 0.001153317, 0.0001900716, 7.32827e-05, 0.00101886, 
    0.000146916, 0.0001285836, 0.0005538696, 0.0003389791, 0.0007516742, 
    0.001634968, 0.002472292, 0.002720152, 0.02057392, 0.02595687, 
    0.0004182424, -0.0001346959, 0.001072657, 0.001391896,
  0.0004282452, 0.002607719, 8.355069e-06, -6.612322e-05, 0.001471123, 
    0.0005946542, 0.0001536534, 0.0001614987, 0.02554177, 0.1020819, 
    0.0002100483, 0.001844705, 9.349026e-05, 0.002766703, 0.0006380974, 
    0.0002845852, 0.0002575873, 0.0002097995, 0.002099707, 0.0001799336, 
    0.002757357, 0.006334252, 0.003105469, 0.001350686, 0.001709882, 
    9.019819e-05, 0.0001812529, 0.0007758065, 0.002088695,
  6.084833e-10, 1.017061e-09, 1.227962e-10, 0.00321248, 0.02017236, 
    0.001103547, -0.001771552, 0.0009580046, 0.0001867539, 0.001656899, 
    0.006553105, 0.0003512561, 0.0002526677, 0.001022456, 0.0003235119, 
    0.001252748, 0.00294071, 0.0002393763, 9.701019e-05, 0.0002049324, 
    0.0004866086, 0.0001499906, 0.1785986, 0.09303821, 0.0001054736, 
    0.0005735603, 0.0009875082, 8.049132e-05, -0.0003303105,
  3.994141e-08, 1.014119e-08, 2.960232e-10, 5.342119e-05, 3.692774e-09, 
    0.0002220362, 3.347838e-08, 0.0007718491, 0.0006823684, 0.0413421, 
    0.003336982, 0.006143405, 0.002683514, 0.002742474, 0.003529635, 
    0.001195972, 0.01713042, 0.005434422, 0.004504478, 0.01224776, 
    0.0001655888, 0.07418834, 0.0002948004, -0.0008406007, 4.810726e-05, 
    0.0005473222, 8.626641e-05, 0.000132742, 2.117339e-07,
  -4.706567e-06, 0.005244996, 0.0001189618, 4.293166e-05, 0.01109284, 
    0.008938954, -0.001577136, 0.003038231, 0.02192892, 0.07187518, 
    0.03721338, 0.0101236, 0.008338107, 0.008927954, 0.0354857, 0.01791714, 
    0.03265167, 0.05014638, 0.02561486, 0.01117708, 0.01044585, 0.1178227, 
    0.03524737, 0.01167453, 0.006154537, 0.005996724, 0.002517011, 
    0.001119217, 0.002375551,
  0.001761073, 4.270059e-05, 0.01465117, 0.1699234, 0.001153517, 0.0519482, 
    0.1404958, -8.471307e-06, -8.907866e-05, 0.002363287, 0.03707331, 
    0.02343349, 0.1003653, 0.0943702, 0.05505799, 0.07180791, 0.1021585, 
    0.08603638, 0.05138674, 0.3395455, 0.1199728, 0.09864713, 0.1572262, 
    0.2152185, 0.07779067, 0.05015587, 0.03990552, 0.02143379, 0.05618985,
  0.04164111, 0.06734905, 0.1495351, 0.4320817, 0.3085915, 0.2175246, 
    0.09439423, 0.1815743, 0.04197256, 0.02246591, 0.004685518, 0.1168257, 
    0.2165826, 0.2740526, 0.2270475, 0.04176418, 0.02619355, 0.01236511, 
    0.07472555, 0.4629199, 0.07819714, 0.123572, 0.1546098, 0.3414105, 
    0.1758286, 0.1243939, 0.04807257, 0.05533979, 0.0393948,
  0.05106748, 0.4202489, 0.4201061, 0.4305539, 0.4246987, 0.390386, 0.420171, 
    0.450166, 0.3675624, 0.3465371, 0.3620558, 0.428795, 0.2756364, 
    0.3281356, 0.03672677, 0.17723, 0.337781, 0.08101919, 0.3102009, 
    0.4001821, 0.3587036, 0.1788361, 0.2335468, 0.1279634, 0.69186, 
    0.0230476, 0.0178158, 0.03883694, 0.03127185,
  0.05718439, 0.01848512, 0.2986531, 0.1465436, 0.5371091, 0.4353926, 
    0.6268629, 0.4430509, 0.3789765, 0.507486, 0.5624866, 0.1869203, 
    0.5821015, 0.335324, 0.2517098, 0.2969781, 0.4499902, 0.2913772, 
    0.4229794, 0.405728, 0.2156609, 0.4444909, 0.3526841, 0.1799395, 
    0.07415411, 0.1616495, 0.2878918, 0.07818433, 0.164937,
  0.5342334, 0.4079553, 0.516954, 0.2324981, 0.2636838, 0.5386238, 0.5313917, 
    0.5226991, 0.5358839, 0.5275622, 0.5408044, 0.5305387, 0.5163396, 
    0.5274541, 0.487445, 0.5062773, 0.5771651, 0.5952985, 0.5633867, 
    0.6117243, 0.6319178, 0.2208048, 0.1901314, 0.213399, 0.09074648, 
    0.09370547, 0.04979284, 0.3224613, 0.4182394,
  0.386596, 0.3897896, 0.3929832, 0.3961768, 0.3993704, 0.402564, 0.4057576, 
    0.3077431, 0.3142216, 0.3207001, 0.3271786, 0.3336571, 0.3401357, 
    0.3466142, 0.4816582, 0.4784112, 0.4751643, 0.4719173, 0.4686704, 
    0.4654234, 0.4621765, 0.4506526, 0.4442274, 0.4378022, 0.4313771, 
    0.4249519, 0.4185267, 0.4121015, 0.3840411,
  0.07288758, 0.06823067, 0.1062184, 0.3677313, 0.5298533, 0.3171964, 
    0.3132456, 0.3041272, 0.1111896, 0.04768471, 0.02712584, 0.005578279, 
    0.02704852, 0.0005743635, 0.1399866, 0.325976, 0.2759046, 0.1810381, 
    0.05210954, 0.2255513, 0.2473972, 0.2607353, 0.1001348, 0.06948552, 
    0.1517487, 0.1685592, 0.1076785, -0.000664375, 0.0346065,
  0.05671597, 0.02101732, 0.02587279, 0.006964793, 0.01877914, 0.1686557, 
    0.01074364, 0.05215422, 0.1245323, 0.1248199, 0.03081212, 0.002552196, 
    0.009520159, 0.001516472, 0.131419, 0.230621, 0.1832315, 0.1855771, 
    0.2174556, 0.1628889, 0.2168178, 0.1739931, 0.1862067, 0.1345712, 
    0.1496132, 0.1176232, 0.09806084, 0.04854487, 0.075229,
  0.1220254, 0.148994, 0.08523498, 0.1426146, 0.1377538, 0.0810255, 
    0.1740681, 0.195488, 0.2985444, 0.2315714, 0.1820545, 0.2117306, 
    0.3075694, 0.2454488, 0.2040428, 0.2062194, 0.2349868, 0.2617361, 
    0.214333, 0.109811, 0.09442194, 0.0711253, 0.05721257, 0.1141545, 
    0.1764317, 0.3070251, 0.2829388, 0.1865537, 0.1753246,
  0.1816717, 0.165812, 0.1976249, 0.1739244, 0.1782408, 0.17681, 0.1535172, 
    0.09374442, 0.09486899, 0.1255694, 0.06889682, 0.06506903, 0.08573499, 
    0.06089296, 0.1239887, 0.2243451, 0.1541337, 0.1319819, 0.1172463, 
    0.08776883, 0.04485859, 0.05038123, 0.07106341, 0.07284967, 0.01623886, 
    0.1013396, 0.1957748, 0.2098975, 0.2338382,
  0.03855342, 0.04129455, 0.02561819, 0.04705258, 0.0673543, 0.08195808, 
    0.01755747, 0.0306119, 0.05916679, 0.05494142, 0.01630829, 0.009771611, 
    0.006995718, 0.02028236, 0.1458399, 0.04898638, 0.05690049, 0.08951213, 
    0.08830424, 0.04744433, 0.03798033, 0.02581941, 0.01037469, 0.07930715, 
    0.02425339, 0.05569953, 0.05171228, 0.02825928, 0.02052109,
  0.004788512, 0.003517591, 0.003190843, 0.0008869623, 0.01807862, 
    0.01819338, 0.0005262185, 0.001495071, 0.006481255, 0.0008998598, 
    0.0001206678, 3.281452e-09, 0.0003033035, 0.008639716, 0.001023592, 
    0.001367739, 0.04113967, 0.09141756, 0.03947593, 0.005082086, 
    0.0005310729, 0.001501004, 0.005873038, 0.001304098, 0.01730247, 
    0.00431473, 0.001259358, 0.0002811132, 0.001069533,
  0.001480469, 0.06604081, 0.0008001218, 0.0004934845, -0.0009618911, 
    0.0001621212, 0.0003486232, 0.001952056, 0.002301761, 0.001245669, 
    0.001193484, 3.611308e-05, 0.001110741, 0.0008484183, 0.001132962, 
    0.0004706332, 0.0002871535, 0.0005398047, 4.922785e-05, 1.763481e-05, 
    8.363835e-06, 0.0004278946, 0.003287056, 0.02013034, 0.01099188, 
    0.0166304, 7.248938e-05, 0.0001927208, 0.0003071374,
  0.007907866, 0.005645988, 0.01336321, 0.03334, 0.0001975357, 0.0002691066, 
    0.003354966, 9.329423e-05, 0.0002679915, -0.0002569481, 0.0007649624, 
    0.0008061821, 9.451402e-05, 5.206522e-05, 0.0006035923, 0.000105007, 
    9.583506e-05, 0.0004123213, 0.000268629, 0.0005473201, 0.001223681, 
    0.001795659, 0.001995908, 0.01232845, 0.0188964, 0.004087465, 
    -9.828615e-05, 0.0008079501, 0.001031658,
  0.000296061, 0.01214136, 8.66923e-06, -4.489831e-05, 0.0005705243, 
    0.000413163, 0.0001143205, 0.0001187606, 0.0322169, 0.09460495, 
    0.0001353685, 0.0012808, 7.393505e-05, 0.001566403, 0.0004721849, 
    0.0001920967, 0.0001824077, 0.000119127, 0.0009010352, 8.992468e-05, 
    0.001261687, 0.004016054, 0.001829502, 0.004678078, 0.002000232, 
    6.712683e-05, 0.0001068001, 0.0005900264, 0.001503113,
  6.869575e-10, 1.011054e-09, 1.011104e-10, 0.005204222, 0.01295946, 
    0.0008250187, -0.001245196, 0.0007215376, 5.681026e-05, 0.001167899, 
    0.002992517, 0.0001701836, 0.0001831464, 0.0007108313, 0.0002367081, 
    0.0007589842, 0.001298276, 0.0001220598, 6.071241e-05, 0.0001484622, 
    0.0002439432, 0.0001103309, 0.135855, 0.0689836, 6.250237e-05, 
    0.0003247689, 0.00073717, 5.645867e-05, -0.0005055568,
  3.836048e-08, 1.008263e-08, 3.100982e-10, 4.412844e-05, 3.084216e-09, 
    0.0001669215, 2.96848e-08, 0.0004394533, 0.0004868499, 0.02411592, 
    0.001149138, 0.00345828, 0.001910607, 0.002076733, 0.002469613, 
    0.0009209265, 0.008134655, 0.004094147, 0.003347159, 0.0092736, 
    0.0001303459, 0.06030396, 0.0002270903, -0.0007824529, 2.151172e-05, 
    0.0003273241, 6.855644e-05, 0.0001021903, 2.077599e-07,
  -3.522223e-06, 0.004670959, 0.0003240836, 2.065133e-05, 0.009125284, 
    0.006207794, -0.001348268, 0.03097375, 0.02066795, 0.06013951, 0.0238599, 
    0.007199388, 0.003813427, 0.004656784, 0.0180204, 0.01031279, 0.01991124, 
    0.0313344, 0.01268239, 0.005700512, 0.00804366, 0.08934659, 0.03227424, 
    0.006972148, 0.004211078, 0.004163253, 0.001536043, 0.0008677834, 
    0.001538424,
  0.0009660558, 2.947427e-05, 0.01299227, 0.1571725, 0.0009397435, 
    0.04384622, 0.1476085, -4.486062e-06, -7.451187e-05, 0.006522106, 
    0.03309425, 0.01992634, 0.081108, 0.07192273, 0.03480353, 0.0450688, 
    0.06894931, 0.06185931, 0.03064646, 0.310191, 0.112644, 0.08391824, 
    0.141265, 0.2017177, 0.05652791, 0.03552279, 0.02477768, 0.01137559, 
    0.03883401,
  0.02949165, 0.06167202, 0.1355352, 0.3967859, 0.2745158, 0.1934142, 
    0.08489073, 0.1780912, 0.07988545, 0.02709701, 0.008686594, 0.1146079, 
    0.2081677, 0.2279857, 0.190147, 0.03548493, 0.02276753, 0.01043368, 
    0.05574274, 0.4244316, 0.06402552, 0.09646226, 0.12864, 0.2956716, 
    0.1509386, 0.1100293, 0.03726469, 0.04014356, 0.02715908,
  0.04108439, 0.417692, 0.3642964, 0.3853824, 0.3708858, 0.3459798, 
    0.3637522, 0.3952959, 0.3095108, 0.3090249, 0.3551847, 0.4533459, 
    0.2932473, 0.2905489, 0.03016529, 0.2029028, 0.3847562, 0.1698502, 
    0.3523257, 0.3487311, 0.3135686, 0.1877351, 0.1460199, 0.1639623, 
    0.6828968, 0.02133868, 0.01505303, 0.03255501, 0.02536668,
  0.04730824, 0.01344143, 0.2944883, 0.1209958, 0.5273039, 0.3461092, 
    0.5355926, 0.4316363, 0.4357288, 0.533584, 0.5415366, 0.2491749, 
    0.6208915, 0.2886924, 0.2165936, 0.2737266, 0.3950646, 0.236746, 
    0.3939789, 0.2266315, 0.2309241, 0.3617877, 0.2868079, 0.1843019, 
    0.07468988, 0.1355006, 0.356108, 0.06441324, 0.1447967,
  0.4975726, 0.4457644, 0.4828103, 0.1649455, 0.2313176, 0.3727833, 
    0.3971488, 0.3917612, 0.4086324, 0.3897488, 0.3654096, 0.3550597, 
    0.3573433, 0.3533494, 0.3676161, 0.4100894, 0.4385992, 0.389422, 
    0.4067966, 0.4442968, 0.3765961, 0.1897815, 0.1437549, 0.2980211, 
    0.109664, 0.05599199, 0.04984264, 0.3342996, 0.3140314,
  0.2883959, 0.2918073, 0.2952187, 0.2986301, 0.3020416, 0.305453, 0.3088644, 
    0.2362673, 0.2422458, 0.2482244, 0.2542029, 0.2601815, 0.26616, 
    0.2721386, 0.381089, 0.3782961, 0.3755032, 0.3727104, 0.3699175, 
    0.3671246, 0.3643318, 0.3336031, 0.327006, 0.3204089, 0.3138117, 
    0.3072146, 0.3006175, 0.2940204, 0.2856668,
  0.08649805, 0.07038835, 0.1029289, 0.3049729, 0.4461772, 0.2990713, 
    0.2775388, 0.2937875, 0.1040758, 0.03964844, 0.02548351, 0.006344243, 
    0.02229742, 0.0002103375, 0.1375307, 0.3150665, 0.2540108, 0.1834893, 
    0.04225731, 0.2005241, 0.2199944, 0.2520149, 0.09068266, 0.07637249, 
    0.1319198, 0.1616234, 0.1088124, 0.007258618, 0.03657698,
  0.0509786, 0.01837038, 0.02246274, 0.007214512, 0.02317568, 0.1546872, 
    0.007921846, 0.0445127, 0.1168815, 0.1253299, 0.04174445, 0.008294237, 
    0.01211664, 0.001399026, 0.101842, 0.1886306, 0.1525273, 0.1539526, 
    0.1710662, 0.1378399, 0.1801106, 0.1487832, 0.1619197, 0.1192263, 
    0.1387693, 0.1029849, 0.08465309, 0.0381264, 0.06288171,
  0.101471, 0.1230223, 0.07165128, 0.1234592, 0.1161713, 0.06751924, 
    0.1416951, 0.1640203, 0.2565148, 0.1850284, 0.144776, 0.1666776, 
    0.2514343, 0.1971565, 0.1609704, 0.1730687, 0.1985545, 0.2320586, 
    0.1804224, 0.09176061, 0.07906107, 0.05661417, 0.0449825, 0.09459096, 
    0.1346493, 0.2416478, 0.2245768, 0.1585304, 0.1496144,
  0.1505391, 0.1401177, 0.1590939, 0.1485808, 0.1521284, 0.1485002, 
    0.1284396, 0.0783225, 0.0771096, 0.1020187, 0.05584188, 0.0490117, 
    0.0596014, 0.04782403, 0.09678578, 0.1701424, 0.1175408, 0.1024481, 
    0.09013198, 0.06740481, 0.03469681, 0.04113876, 0.05842061, 0.07687696, 
    0.01425136, 0.07986314, 0.1615734, 0.1762352, 0.1974209,
  0.0278907, 0.02865359, 0.01631643, 0.03070284, 0.04817159, 0.05651623, 
    0.01283066, 0.02162121, 0.03863429, 0.0376993, 0.01316855, 0.007435487, 
    0.005312834, 0.01110819, 0.1380858, 0.02819659, 0.03426408, 0.06622399, 
    0.06006492, 0.03554776, 0.02661896, 0.01790402, 0.007233029, 0.0841499, 
    0.01830726, 0.04205443, 0.0351437, 0.01859684, 0.01505109,
  0.003699299, 0.002762658, 0.01072316, 0.0006931161, 0.01043026, 0.01131811, 
    0.000424372, 0.001255134, 0.005322515, 0.0006991376, 8.375633e-05, 
    6.152053e-09, 0.008869923, 0.006095232, 0.0008104793, 0.00100202, 
    0.02367132, 0.05494905, 0.02446278, 0.00350861, 0.0004311876, 
    0.001245894, 0.004882995, 0.0009345773, 0.01848941, 0.002629191, 
    0.001049644, 0.0002249522, 0.0007760784,
  0.001198224, 0.0536439, 0.0007378936, 0.0003406284, -0.001131842, 
    0.0001307034, 0.000276437, 0.001306729, 0.001891186, 0.0009834298, 
    0.002294083, 1.821422e-05, 0.0008868277, 0.0006634085, 0.0007336724, 
    0.000344764, 0.0002339065, 0.0004151419, 4.134986e-05, 1.49197e-05, 
    6.732344e-06, 0.0003335501, 0.002624674, 0.01623788, 0.01702151, 
    0.02755209, 6.020107e-05, 0.0001589044, 0.0002488587,
  0.006487844, 0.004474102, 0.05181159, 0.1219953, 0.0001504658, 
    0.0002137518, 0.002144448, 7.741088e-05, 0.0001894516, -0.0001901056, 
    0.0005306251, 0.0006488895, 7.531946e-05, 4.037057e-05, 0.0004362519, 
    8.426767e-05, 7.702944e-05, 0.0003407446, 0.0002319377, 0.000450354, 
    0.001024971, 0.001465211, 0.001635795, 0.04205901, 0.03262954, 
    0.03997837, -0.0001647074, 0.0006759421, 0.0008509936,
  0.0002339579, 0.07100427, 0.0002202215, -4.604274e-05, 0.000372994, 
    0.000331682, 9.482639e-05, 9.888915e-05, 0.05235461, 0.09219306, 
    0.000106564, 0.001019371, 6.32513e-05, 0.00107146, 0.0003866341, 
    0.000153046, 0.0001490314, 8.734959e-05, 0.0005075336, 6.183262e-05, 
    0.0007324233, 0.0030854, 0.001368677, 0.1010441, 0.05176282, 
    5.373512e-05, 7.634955e-05, 0.0004949199, 0.00121314,
  7.858534e-10, 1.008171e-09, 8.624347e-11, 0.006766953, 0.009066936, 
    0.0007277055, -0.001003015, 0.0006072439, -0.0004694685, 0.0009581277, 
    0.001911174, 0.0001192147, 0.0001528758, 0.0005828708, 0.0001975746, 
    0.0006029414, 0.0007791466, 8.886122e-05, 4.774164e-05, 0.0001243826, 
    0.0001725748, 9.309634e-05, 0.1660594, 0.06250599, 4.794988e-05, 
    0.0002496788, 0.0006241738, 4.581614e-05, -0.001247516,
  3.791493e-08, 1.006241e-08, 3.151003e-10, 3.953811e-05, 2.860264e-09, 
    0.0001409772, 2.76508e-08, 0.0003128187, 0.0007159355, 0.01716492, 
    0.0007638871, 0.002388202, 0.001528263, 0.001749085, 0.002048213, 
    0.0007843822, 0.004844881, 0.003423422, 0.002778686, 0.00781503, 
    0.0001123832, 0.0530377, 0.0001933874, -0.001199369, 1.480395e-05, 
    0.0002460747, 6.116534e-05, 8.90991e-05, 2.082578e-07,
  -5.324461e-06, 0.004427525, 0.001173568, 1.293268e-05, 0.008761679, 
    0.004834773, -0.001335701, 0.1293188, 0.02532726, 0.05218972, 0.01650933, 
    0.005924221, 0.002403504, 0.003245356, 0.01033112, 0.006988476, 
    0.01404573, 0.02030465, 0.007145264, 0.003817086, 0.006853843, 
    0.08760978, 0.04270152, 0.005215785, 0.003368737, 0.003346058, 
    0.001167565, 0.0007449098, 0.001292118,
  0.0009603078, -2.443693e-05, 0.01369661, 0.1519816, 0.0007449108, 
    0.03821911, 0.1786131, -2.544309e-06, -6.626239e-05, 0.009399982, 
    0.03554361, 0.01837162, 0.07141757, 0.05710109, 0.02494475, 0.030612, 
    0.05291188, 0.04598786, 0.02121735, 0.2995988, 0.1095227, 0.08546414, 
    0.1578082, 0.1769401, 0.0470773, 0.02748073, 0.01672639, 0.007208412, 
    0.03289286,
  0.02421998, 0.06246754, 0.1357216, 0.4076743, 0.2620339, 0.1740237, 
    0.08370686, 0.2199686, 0.170855, 0.03775978, 0.03256478, 0.1386172, 
    0.2005087, 0.2023412, 0.1653875, 0.03223503, 0.02089628, 0.00948994, 
    0.04565731, 0.4202752, 0.06511096, 0.09396205, 0.1411833, 0.2898442, 
    0.1388597, 0.1004707, 0.03228775, 0.03319972, 0.02171705,
  0.03584177, 0.5021887, 0.3664314, 0.3784012, 0.3699349, 0.3445821, 
    0.3513713, 0.3786767, 0.3164305, 0.3247389, 0.3960572, 0.6012184, 
    0.3361197, 0.2984585, 0.02674935, 0.1911092, 0.4803934, 0.215085, 
    0.4102632, 0.3482638, 0.2987822, 0.2039907, 0.1149854, 0.227889, 
    0.6806852, 0.02423797, 0.0139314, 0.03047268, 0.02242172,
  0.03906835, 0.01143244, 0.3445905, 0.1076844, 0.5240797, 0.3150688, 
    0.3516525, 0.3764647, 0.4634033, 0.5148143, 0.6032502, 0.4529405, 
    0.5067208, 0.3221563, 0.2098135, 0.2387497, 0.369696, 0.2660057, 
    0.3317767, 0.1575713, 0.207701, 0.3204229, 0.2093219, 0.1871427, 
    0.06169198, 0.1284634, 0.4982703, 0.06341492, 0.1362304,
  0.5009972, 0.4840122, 0.4160277, 0.1582409, 0.189665, 0.2719016, 0.2880238, 
    0.2838203, 0.2953075, 0.2975776, 0.2851962, 0.2438913, 0.2788351, 
    0.2584619, 0.2832715, 0.324168, 0.2995856, 0.2633533, 0.293368, 
    0.3244486, 0.2716142, 0.1793309, 0.1853205, 0.3102144, 0.11243, 
    0.008155422, 0.0546088, 0.3494411, 0.2158951,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -2.335356e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, -9.313262e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -8.040414e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -6.227616e-06, 0, 0, 0, 0, 0, 0, 0, 
    1.409831e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, -4.280618e-05, 0, 0, 0, 0, 2.453809e-05, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, -3.450561e-07, 0, -2.445523e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -5.62829e-05, 6.820949e-05, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.000463355, 0, 0, 0.0005854152, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.254842e-05, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -1.678706e-05, 0, 0, 0, 0, 0, -1.459644e-05, 0, 
    0.0002973337, 0, 0, 0, 0, 0, 0, 0, 0.0002698145, 0, 0, 0,
  0, 0, 0, -6.166923e-05, 0, 0, 0, 0, 0.002809059, 0, 0, -4.632199e-05, 0, 0, 
    0, 0, 8.026962e-05, -3.936612e-06, 0, 0, 0, 0, 0, -2.537607e-05, 
    -1.493722e-05, -4.000093e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -2.53783e-05, 0, -0.0001459226, 1.22146e-05, 0, 
    0, -4.431267e-07, -2.769684e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.004062513, 0, 0, 0.001421171, 0, 0, 0, 0, 0, 0, 0, 
    0, -1.828724e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3.265659e-05, 0, 0, 
    -1.270975e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, -2.582577e-05, 0, 0, -9.972743e-06, 0, 0, -3.730685e-06, -3.141208e-06, 
    -1.912241e-05, 8.020307e-06, 0, 0, -2.802402e-06, -1.570318e-05, 
    -6.286265e-05, -1.396269e-05, 0.0005391266, 0, 0, 0, 0, 0, 0, 0, 
    0.002196083, -0.0001602824, 0, 0,
  0, 0, -5.761411e-05, -7.264893e-05, -5.889182e-06, 0, 0.001165387, 0, 
    0.007415161, 0, 0, 0.0003847737, 0, 0, 0, 0.001100721, 0.002052249, 
    0.0001978549, 0, 0, 0, 0, 0, 0.001364515, 0.001552849, 0.0006526422, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, -1.046252e-05, 0.000252384, 1.538837e-05, 
    -0.0001547595, -5.684474e-05, 0, -4.978395e-07, -3.99232e-06, 
    -3.719049e-05, -2.395295e-05, 0, 0, 0, 0, 0, 2.873803e-05, 4.190023e-05, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.01018702, 0, 0, 0.001649412, -5.1528e-05, 
    -8.756555e-06, -3.142144e-06, 0, 0, 0, 0, 0, -9.357285e-05, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3.698343e-08, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, -8.889494e-06, 0, 0, 0, 0,
  0, 0, 0, 0, 4.167712e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0001381861, 
    0, 0, -4.289313e-05, 0, 0, 0, 0, 0, 0, 0.0005933797, 0, 0,
  0, -8.114467e-05, 0, 0, 0.002689954, 0, -3.431074e-05, -4.864709e-05, 
    -6.428449e-05, -3.123876e-05, 5.85377e-05, 0, 0, -8.732959e-05, 
    -4.82574e-05, 0.0002456452, -0.0001191414, 0.0006372653, -8.212277e-06, 
    0, 0, 0, 0, 0, 0.0005671489, 0.00427305, -0.0002584062, 0, 0,
  0, 0.0005820931, 0.0003409697, -8.289535e-05, 1.118888e-06, -2.885475e-06, 
    0.00354047, -5.128809e-06, 0.01683659, 0, 0.0009143973, 0.0004599465, 
    0.0001025511, 0, 0, 0.008758157, 0.005161304, 0.0008853762, 
    -0.0001495645, 0, 0, -4.21457e-05, 0, 0.004481512, 0.004406955, 
    0.000885699, 0, 0, 0,
  0, 0, 0, 0, -6.794214e-06, 0, 0, 0, 0.0004752009, 0.001089847, 
    0.0003308885, 8.314686e-05, -0.0001082555, 2.482497e-06, -4.981568e-06, 
    -1.011854e-05, -8.420695e-05, -8.287052e-05, 0, 0, 0, 0, 0, 4.539554e-05, 
    0.001252136, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.01160482, -1.797585e-05, 0, 0.002066019, 
    -0.000156059, 0.0003437364, -6.822954e-05, -3.109172e-06, 0, 0, 0, 
    -1.135622e-08, -0.0001898321, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.410352e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -4.844347e-06, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, -5.653981e-07,
  0, 0, 0, -4.81223e-06, -6.505548e-06, 0, -1.178216e-05, 0, 0, 0, 
    0.0005943868, 0, 0, -1.08256e-05, 0, 0, 0, 1.091555e-06, 0, 0, 0, 
    0.0002969374, 0, 0, -2.116259e-05, -2.082306e-06, 0, 0, 0,
  0, 0, 0, 0, 0.001060565, 8.42608e-05, 0, 0, 0, 0, 0, 0, -2.018034e-05, 
    -2.699561e-05, 0, 0, 0.000259442, 0, -6.655608e-06, 0.0002672286, 0, 0, 
    0, 0, 0, 0, 0.001822453, 0, 0,
  0, -0.0001718279, 0, 0, 0.01761856, 0, 0.001952016, -0.0003744988, 
    -0.0001759421, -9.941705e-05, 0.0002103203, 0, 0, -0.0003389492, 
    -0.0001082352, 0.008537478, -9.387164e-05, 0.002290814, -7.391049e-05, 0, 
    0, 0, 0, 0, 0.002107452, 0.008329534, -0.0004726992, 0, 0,
  0, 0.001803023, 0.001642029, -7.217868e-05, 0.000218323, -4.838814e-05, 
    0.006689023, 0.0005673894, 0.02500561, 0, 0.003140739, 0.002281768, 
    0.0004202856, 0, -5.457245e-05, 0.01259147, 0.008389702, 0.001607857, 
    0.0003289182, 0, 0, -0.0001883438, 0, 0.01053006, 0.006963173, 
    0.002894592, -8.918571e-06, 0, 0,
  0, 0, 0, 0, -1.899817e-05, 0, 0, 0, 0.001020904, 0.001877123, 0.0008515723, 
    0.001204497, -9.960175e-06, 0.0001395609, -1.734789e-05, 0.0004365567, 
    0.0001110869, -0.0001579013, 0, 2.843211e-05, 0, -2.859041e-05, 0, 
    5.779613e-05, 0.001921355, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.01256158, -8.74055e-05, 1.38214e-05, 0.004563197, 
    -0.0001311586, 0.001273911, -0.0001703238, -4.559563e-05, -0.0001189246, 
    -2.261607e-05, 0, 0.000325765, 0.002151018, 0, -2.894903e-05, 0, 0, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.140715e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.423838e-06, 0, 0, 0, 0, 0, 
    0.0003652426, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -7.737015e-05, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.765183e-05, 0, 0, 0, 0, 0, 0, 0, 
    -8.898014e-05, 0, 0, 0, 0, 0, -1.563804e-05, 0.0003841702, 0, 
    -1.130796e-06,
  0, 0, 0, -5.903518e-05, 8.873785e-06, -4.037114e-05, -8.221459e-05, 
    -2.709496e-05, 0, -7.893641e-05, 0.001767881, 0, 0, 0.001095355, 0, 0, 
    -2.493565e-05, 0.0008250833, 0, -8.188878e-05, -5.942813e-06, 
    0.004382767, 0, 0, -6.805457e-05, 0.003181561, -8.151837e-05, 0, 
    5.935756e-05,
  0, 0, 0, 0, 0.004172366, 0.0001697741, 0, 0, -3.921684e-05, 0, 
    0.0006659069, 0, -0.0001744469, 0.001246389, 0, -8.019309e-05, 
    0.00329428, -7.567519e-05, -9.374202e-05, 0.003478464, 0.000175259, 
    -5.099984e-05, 0, 0, 0.0008551415, 0, 0.01002776, 0, 0,
  0, -0.0003104544, 1.248406e-05, 0, 0.032918, 0, 0.009623791, -0.0006643012, 
    0.0001143471, -0.0001954392, 0.005122287, -6.890402e-08, 0, 
    -0.0006348079, 0.002345926, 0.02120587, 0.0007614034, 0.005291422, 
    -0.0001741325, 0, 0, 0, 0, 0, 0.004781248, 0.01112992, 0.0006366638, 0, 0,
  0, 0.003242043, 0.005801374, -4.693164e-05, 0.0004049309, -0.0001044809, 
    0.01474375, 0.00257914, 0.03838715, 0, 0.004897753, 0.007123843, 
    0.0005771547, -7.021592e-05, -8.742698e-05, 0.021698, 0.01122982, 
    0.003138578, 0.003428553, 0, 0, 0.001103289, 0, 0.01493301, 0.01478174, 
    0.004389155, -8.918571e-06, 0, 0,
  0, 0, -2.0341e-05, -4.395229e-06, -4.895217e-05, 0, 0, -3.027052e-05, 
    0.00256068, 0.002400136, 0.003764184, 0.007532208, 0.008342364, 
    0.000165426, -7.350981e-05, 0.005004602, 0.000412927, 0.00157912, 0, 
    5.961089e-05, 0, -3.891748e-05, 0, 0.0004788623, 0.003511478, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.0137184, -0.0003022415, 0.003844063, 0.006307898, 
    0.004754033, 0.002223938, -0.0002865917, -0.0001058163, -0.0003910966, 
    -0.0002156617, -1.724475e-05, 0.001003474, 0.01120372, -1.444379e-05, 
    -0.0001210628, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.008634e-05, 0, 0, 0, 0, 0, 0, 0, 
    -2.711834e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -9.769531e-06, 8.075364e-06, 0.0002530128, 0, 0, 
    0, 0, 0, 0.006227547, 0, 0, 0, 0, -1.66428e-05, 0, -5.941625e-05, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0002810417, -1.128948e-07, 0.0001503697, -1.044859e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 5.695336e-06, 0, 0, -6.486355e-05, 0.000500498, 0, 0, 
    0.002006322, 0, 0, 0.0007898954, 0, 0, 0, -1.809837e-06, 0.00202912, 0, 
    0, -8.741973e-07, -1.130064e-06, -5.684772e-06, 0.001911762, 0.002202004, 
    -1.922738e-05, 4.347125e-06,
  0, 0, 0, 0.000824509, 0.005856973, 0.000190466, 0.0045063, 0.002483142, 0, 
    -0.0001298383, 0.004313005, 0, -1.936764e-05, 0.002840663, -6.378564e-05, 
    0, 0.006483181, 0.005998397, 0, 0.0001993304, 0.0004852222, 0.007852416, 
    0, 0, 0.0004023692, 0.008207927, 0.001322949, -5.276098e-06, 0.0001488314,
  0, 0, 0, 0.0009290656, 0.007738167, 0.001331562, -8.364316e-05, 
    -0.0001172162, 0.000578702, 1.518092e-08, 0.006388732, 7.624155e-07, 
    0.001352304, 0.006979762, 0, -0.0002094331, 0.01706533, 0.0005827738, 
    0.004832467, 0.006809401, 0.004021934, -0.0002717854, 0, 0, 0.004106374, 
    0.0007368538, 0.02015253, 0, 0,
  0, 0.0002155479, 0.0005932311, 0, 0.05392312, -3.208794e-05, 0.02631178, 
    0.003841294, 0.005761172, -0.0002008824, 0.01278374, -1.202487e-07, 0, 
    0.0009437226, 0.01201984, 0.04352557, 0.009420968, 0.0196569, 
    -0.0004347601, 0.0001182105, 0, 0, 0, 0.0003823758, 0.01092499, 0.016253, 
    0.007397687, 0, 0,
  0, 0.007321548, 0.0143812, 0.001150119, 0.00140352, 0.0002739744, 
    0.02760853, 0.004110309, 0.05055393, 9.672603e-05, 0.005645758, 
    0.01558453, 0.0009961857, 0.002272435, -0.0001128786, 0.02965497, 
    0.0173559, 0.02203657, 0.007008143, 0, 0, 0.001370079, 0, 0.02265034, 
    0.02555113, 0.009478202, -3.640856e-05, 0, 0,
  0, 0.0007954382, 5.377723e-05, 0.0005202718, -0.0001365747, 0.001654958, 
    0.0006895232, -2.676623e-05, 0.006219078, 0.0111867, 0.009459273, 
    0.02741534, 0.02013341, 0.0006151285, 0.001598098, 0.01014523, 
    0.0008510635, 0.008770447, 0, 0.001272696, 0, 0.0006729207, 0, 
    0.01411626, 0.01054153, -2.059356e-06, -1.446014e-05, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.01823676, 0.001239303, 0.007741528, 0.01479653, 
    0.01620638, 0.005270582, 0.0003374981, -0.0002619672, 0.001689697, 
    0.004006298, 0.001448311, 0.007829576, 0.02089011, -5.788642e-05, 
    -0.0002929013, -5.813177e-06, 0, 0, 0, -3.335452e-07, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0006154258, 0, 0, 0, 0, 1.135156e-05, 
    0.006573939, 0.001699281, -5.072313e-05, 6.188312e-06, 0, -1.167734e-05, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0003602626, 0.003090318, 0.003063297, 
    -1.925472e-05, 0, 0, 0, -9.525336e-05, 0.01557611, 3.592995e-06, 0, 0, 
    -2.26325e-05, -6.912314e-05, -1.964966e-05, 8.862129e-05, -6.755534e-06, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.948811e-05, -5.122118e-05, 0, 
    0.001147269, 0, 4.015659e-05, 0, 0, -9.408275e-06, 0.003273922, 
    0.0001879636, 0.001861375, 0.0005368275, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -6.630714e-05, 0, 0, 0, 0, 0, 0, -5.608098e-06, 0, 0, 0, 
    -7.869857e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.001754463, -4.820906e-05, 0, -8.202715e-06, 0.001759687, 0, 0, 
    0.002143819, 0.006158287, 0, 0.0004392668, 0.003445985, 2.358007e-05, 
    -5.277465e-05, 0.002759519, -6.09583e-06, 0, 0.001498776, 0.004435879, 
    0.007728452, -1.852637e-05, 0, 0.0001899102, 0.0008741998, 7.247323e-05, 
    0.006293999, 0.004909399, 0.0007542581, 0.001090796,
  0.002727364, -0.0001982952, 0, 0.002549183, 0.008683086, 0.009599346, 
    0.01097172, 0.004897724, 0, 0.004225944, 0.008555977, 0, -6.720112e-05, 
    0.009709909, 0.001939553, -0.0001824542, 0.01453151, 0.0113296, 
    0.0002715531, 0.003305857, 0.006817734, 0.0152292, 1.491482e-05, 0, 
    0.003527207, 0.01731586, 0.004149782, 0.0004684434, 0.002701775,
  0, 0, 1.033026e-05, 0.005221358, 0.01066126, 0.006255471, 0.00299532, 
    0.002378633, 0.008683286, 6.894306e-05, 0.01990247, 2.854424e-05, 
    0.00742464, 0.01489007, -5.531318e-07, 0.001817959, 0.04529428, 
    0.008006796, 0.01786037, 0.009973298, 0.02040471, -1.841541e-05, 0, 0, 
    0.006188521, 0.005054099, 0.03602865, -2.455427e-05, 1.614858e-06,
  0, 0.005084841, 0.001565443, 0, 0.07808634, -0.0002379089, 0.03743846, 
    0.01075602, 0.01697677, 0.0004532121, 0.03385331, 0.0001402944, 
    -2.956093e-07, 0.005653086, 0.01968505, 0.08302154, 0.02635185, 
    0.04117011, 0.002054421, 0.001462691, 0, 0, 0, 0.003906577, 0.01738579, 
    0.03259693, 0.02478114, -2.713816e-06, 0,
  0, 0.02100038, 0.03017059, 0.006123586, 0.01075047, 0.00791521, 0.04977937, 
    0.01902547, 0.08444695, 6.629415e-05, 0.008676979, 0.05186484, 
    0.003012397, 0.005593315, 0.0003521098, 0.04710446, 0.03739682, 
    0.04262539, 0.01069693, -4.802329e-06, -1.375228e-05, 0.003467433, 0, 
    0.06713528, 0.07123335, 0.02666419, 0.0005480803, 0, 0,
  0, 0.001375526, 0.0003884757, 0.0005237838, 0.0002405261, 0.002046886, 
    0.01110326, 0.0005830958, 0.02254345, 0.04823983, 0.0157925, 0.04489825, 
    0.0435545, 0.01582767, 0.02009735, 0.02221661, 0.003648027, 0.02364125, 
    -4.406787e-06, 0.004611049, 4.552657e-07, 0.004724899, 9.645274e-07, 
    0.033155, 0.02302014, 4.646073e-05, 1.840339e-05, 0, 0,
  -9.108402e-10, 0, 0, 0, 0, 0, 2.600553e-05, 0.0295427, 0.004259333, 
    0.009889224, 0.03895234, 0.02467306, 0.01173511, 0.006486055, 
    0.001113281, 0.01296047, 0.01037459, 0.003445749, 0.01941826, 0.02901155, 
    -0.0001822683, -0.0001596339, -2.959152e-05, 0, -1.736812e-10, 
    -1.673987e-09, -2.022963e-08, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.004290997, -1.51163e-05, -9.566052e-10, 
    0, -1.494382e-05, 0.0008247469, 0.01637721, 0.01938927, 0.0119423, 
    0.01064412, 0.0005070549, 0.0003644387, 5.949381e-08, 0, 0, 0, 
    -1.743194e-10, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002015918, 0.008096869, 0.005292714, 
    0.001408698, -1.519918e-05, 0, -4.160748e-05, -9.850697e-05, 0.01699685, 
    0.002271865, -0.0001299314, -4.985908e-05, 1.725915e-05, 0.001181217, 
    -7.192413e-05, 0.001485733, 0.002331617, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0.00013307, 8.743785e-05, 0.002300709, 
    -7.987111e-05, 0.002542057, 0, 0.001439425, 0, 0, 0.004323561, 
    0.006677403, 0.005508939, 0.00879578, 0.002335947, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -7.93905e-06, 0, 0, 0, 0, 0, 0, 
    0, 0.0002351513, 0, 0, 0.003712556, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, -1.983617e-06, 0.0003375594, 0, 0, -6.045975e-07, 0, 0, 0, 
    0.001360465, 0, 0, 0, 0.001100283, 0, 3.266842e-05, 0, 0, 0, 0, 0, 0, 
    -5.915153e-05, 0, 0,
  0.005887319, 0.003228403, 0, 0.003034719, 0.01028473, -0.0001521688, 
    0.0008955277, 0.005550893, 0.01607847, 0.002821093, 0.00317377, 
    0.003522434, 0.002197961, 0.00423161, 0.005193838, -1.05654e-05, 
    0.002722406, 0.009804692, 0.009245683, 0.01408101, 0.001801572, 
    -1.634841e-05, 0.01173772, 0.005986978, 0.00184626, 0.01296296, 
    0.01471684, 0.00718856, 0.0008767928,
  0.01352763, 0.002702255, 0.0003450209, 0.006118081, 0.01683733, 0.02922256, 
    0.02995938, 0.009948919, 0.0003389628, 0.01645547, 0.01569401, 
    -2.398836e-07, 0.001770679, 0.02477246, 0.01219805, 0.001335973, 
    0.01933433, 0.01833657, 0.006349931, 0.01102113, 0.0282768, 0.02185894, 
    0.0009478347, -2.631657e-05, 0.008136263, 0.03034225, 0.02054037, 
    0.004888111, 0.02581088,
  -6.932417e-05, -1.567533e-08, 0.001426803, 0.01161555, 0.01463603, 
    0.02271468, 0.05767476, 0.01663634, 0.02865042, 0.002682331, 0.03318124, 
    0.002196264, 0.01027227, 0.02931841, 0.0003734207, 0.009942993, 
    0.0834097, 0.04564498, 0.03602907, 0.03035147, 0.04064426, 0.003708369, 
    -2.478087e-05, 6.964344e-05, 0.007119195, 0.01487123, 0.06356557, 
    0.001443716, 0.0003479375,
  0, 0.02772128, 0.002934141, 0.0003086268, 0.1296883, 0.01715207, 0.0485881, 
    0.02206505, 0.1332988, 0.02266474, 0.1050318, 0.01774458, 0.003032101, 
    0.07736141, 0.1039461, 0.1647027, 0.0709237, 0.1386097, 0.009100166, 
    0.006398967, -1.855828e-06, -2.020416e-10, -0.0002133089, 0.03768311, 
    0.07836348, 0.04746311, 0.04611684, -9.000398e-05, 0,
  7.065025e-09, 0.03890875, 0.09463982, 0.0298023, 0.07593734, 0.0611061, 
    0.1335375, 0.09640361, 0.2599619, 0.02658661, 0.02875988, 0.2656009, 
    0.05642072, 0.06886808, 0.01699993, 0.1276071, 0.1460941, 0.1025308, 
    0.03294499, -4.127426e-05, -7.554093e-05, 0.0111476, 0.003182924, 
    0.1925954, 0.2664786, 0.09306287, 0.01014088, 1.884582e-05, -1.664204e-10,
  -2.483116e-06, 0.007118235, 0.009745685, 0.006074591, 0.002590413, 
    0.01209608, 0.04076969, 0.05062003, 0.07489646, 0.1291551, 0.08037556, 
    0.1409176, 0.1716086, 0.1422792, 0.1390623, 0.09568989, 0.05288696, 
    0.04690654, -4.071503e-05, 0.01486558, -0.0002090026, 0.02015883, 
    0.0002498244, 0.1506872, 0.07450594, 0.002365949, 0.0003960612, 
    -3.34029e-05, -2.532757e-07,
  -4.184404e-05, -1.359394e-05, 0.0008400036, 0, -1.237648e-09, 1.146762e-07, 
    0.001091758, 0.07659981, 0.0324182, 0.04714723, 0.1060265, 0.07992266, 
    0.09625687, 0.04423138, 0.04085005, 0.05352641, 0.02625814, 0.009680414, 
    0.03518683, 0.04099017, 0.0007466214, 0.001460997, 0.001549807, 
    -3.503012e-07, 4.818255e-06, 6.19345e-05, 0.0001151404, 4.573091e-05, 
    -3.588626e-05,
  0, -2.089132e-08, -4.284561e-08, 1.435693e-06, 0, 0, 0, 0.0008857516, 
    3.172167e-05, 4.887344e-05, 1.672023e-05, 0.008718207, 0.0009584764, 
    8.074839e-06, -6.191028e-09, -0.0001612486, 0.007204247, 0.03342731, 
    0.06492604, 0.03036638, 0.04301459, 0.01099891, 0.0008137271, 
    5.404496e-05, 0.0002644465, -5.885504e-13, 0, 0.000121488, -2.771033e-05,
  0, 0, 0, 0, -2.001465e-05, 0, 0, 0, 0, 0.01212697, 0.02007575, 0.01091784, 
    0.004037409, 0.000571252, 0.0001024557, -0.0001633024, 0.003070803, 
    0.02089636, 0.01341654, 0.001409065, -0.0002150831, 0.01570556, 
    0.00311407, 0.008506307, 0.005413406, 0.01243295, 0, -3.972774e-09, 0,
  0, 0, 0, 0, -3.387943e-05, 0, 0, 0, 0, 0, 0, 0, 0.001191813, 0.004058597, 
    0.004992638, 0.0005778131, 0.01029026, 0.001924669, 0.003128588, 
    -2.000095e-05, 0, 0.01148518, 0.01705467, 0.01723919, 0.01594573, 
    0.02784251, -3.86289e-06, -8.797464e-06, 1.288975e-05,
  0, 0, 3.900434e-05, 0, 0, 6.499092e-05, 0, 0, 0, 0, 0, 0, 0, 0, 
    -2.059957e-05, 0, 0, 0, 2.793443e-05, 0.0001522149, 0, 0, 0.001112517, 0, 
    5.278671e-05, 0.006514114, 9.287911e-05, 0.0001185209, 6.8351e-06,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, -1.969745e-05, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0004895544, 1.760836e-05, 0, 
    0.00255983, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, -8.966484e-07, 0.0006049295, 0, -1.215159e-05, -2.912676e-05, 
    0.0004882906, 7.103125e-06, 0, -1.82875e-05, -3.720301e-05, 8.938008e-05, 
    -2.528482e-05, 0.004640026, 0.0002105376, -1.038115e-06, -2.074653e-05, 
    0.005081286, -0.0001265105, 0.004716099, 0, 0, -3.66196e-05, 
    -1.349623e-06, 0, -3.143305e-05, -0.0001358723, 5.486679e-05, 0.0005056512,
  0.02304611, 0.009023225, -1.029655e-06, 0.006045876, 0.02999425, 
    0.003339804, 0.0008867735, 0.00996604, 0.02140085, 0.004035119, 
    0.01102009, 0.004876521, 0.004287153, 0.008283739, 0.01388836, 
    -4.470756e-05, 0.00799296, 0.02410845, 0.01751298, 0.02213939, 
    0.007523383, 0.001150418, 0.0264377, 0.01621747, 0.005200746, 0.02669081, 
    0.02530159, 0.01342681, 0.005535908,
  0.01833264, 0.008772608, 0.001974312, 0.01282929, 0.02982913, 0.05520506, 
    0.05015833, 0.0197395, 0.00196958, 0.02390954, 0.02770516, 0.0008241177, 
    0.003037147, 0.0378353, 0.02549409, 0.007322043, 0.03619183, 0.03168094, 
    0.02708622, 0.02994964, 0.04877362, 0.05104155, 0.002570009, 
    0.0004575352, 0.02273898, 0.04021307, 0.0539953, 0.05880985, 0.05840598,
  0.007730673, 0.0005217675, 0.01087942, 0.03830522, 0.1012734, 0.0970233, 
    0.1509889, 0.0863331, 0.07604107, 0.06473431, 0.09155712, 0.0536189, 
    0.02138251, 0.08694163, 0.09254133, 0.07032249, 0.164227, 0.2183758, 
    0.1575712, 0.07970686, 0.07457671, 0.06640555, 0.0007971223, 0.02056324, 
    0.05694234, 0.05158108, 0.1741549, 0.08545129, 0.04015093,
  1.012737e-06, 0.0830169, 0.04269587, 0.004615622, 0.1924221, 0.01913268, 
    0.04835261, 0.03238389, 0.2122987, 0.03052856, 0.162584, 0.0406093, 
    0.0066363, 0.08131174, 0.1737995, 0.1933667, 0.1074224, 0.1536939, 
    0.07648818, 0.1295163, 0.002263788, 0.0002964173, 0.01587726, 0.04229106, 
    0.1330774, 0.2007529, 0.1303014, 0.05243509, -3.343893e-05,
  0.01204125, 0.08588955, 0.2772055, 0.2083569, 0.1656136, 0.089967, 
    0.1519621, 0.1372419, 0.2474801, 0.02494534, 0.03831411, 0.207432, 
    0.03546986, 0.05593611, 0.01636674, 0.1204972, 0.1235496, 0.09854943, 
    0.08892302, 0.008331232, 0.0002058306, 0.008272303, 0.01402608, 0.355793, 
    0.3502289, 0.3367234, 0.09989679, 0.005977073, 0.0003400933,
  0.002277873, 0.1831145, 0.2580124, 0.06467691, 0.03945375, 0.0404526, 
    0.1437608, 0.2101066, 0.2483823, 0.3472684, 0.08438856, 0.1195991, 
    0.1475364, 0.122322, 0.09060945, 0.05452449, 0.02508318, 0.05769511, 
    0.0003791209, 0.01785038, 0.0006741887, 0.02103984, 0.06471392, 
    0.4082085, 0.1894163, 0.07109237, 0.1007543, 0.03944334, 0.0006866052,
  0.001652498, 0.002981255, 0.0003067018, 0, -0.0002449887, -1.855085e-05, 
    0.02035919, 0.1050759, 0.04091734, 0.03512688, 0.09122565, 0.05500562, 
    0.06850819, 0.02865042, 0.01464855, 0.05407245, 0.02634242, 0.0244203, 
    0.04522871, 0.1208204, 0.07661381, 0.009161979, 0.02365344, 0.000185792, 
    0.001165189, 0.006405198, -0.0003257009, 0.06026909, 0.01873564,
  0.0008461254, -5.53242e-06, 2.603949e-05, 2.486392e-05, 4.149144e-07, 
    -8.951909e-10, 4.34209e-09, 0.002472327, 0.0005291426, 0.001157076, 
    0.0001158301, 0.0146042, 0.002938705, 0.0009158615, 4.348128e-07, 
    -0.0002242082, 0.0447658, 0.07771508, 0.1253917, 0.09229188, 0.2460568, 
    0.06435524, 0.002078811, 0.0047602, 0.003496376, -7.62538e-05, 
    -3.108966e-06, 0.001364028, 0.0008141874,
  -3.456384e-08, 0, 2.316341e-05, 8.18116e-09, 2.220236e-05, -5.134673e-07, 
    0, 0, -1.147667e-07, 0.03998287, 0.04754119, 0.03315292, 0.01073301, 
    0.02459226, 0.01540809, 0.01069051, 0.02376698, 0.03006389, 0.02620918, 
    0.01295797, 0.003096019, 0.05360246, 0.03441906, 0.02360384, 0.02023033, 
    0.02351288, -4.876306e-05, 0.004082184, 0,
  0, 0, 0, 0, 0.00121051, -3.437906e-08, 0, 0, -2.392344e-06, 0, 
    0.0005675842, -6.499564e-05, 0.009549658, 0.01865028, 0.01261219, 
    0.01329451, 0.02379312, 0.008596428, 0.01159335, 0.0007439959, 0, 
    0.01812182, 0.02880481, 0.03557123, 0.02915177, 0.05681143, 0.001236972, 
    0.006887202, 0.0004944588,
  0, 0, 0.0003817929, 0, 0, 0.0003181329, 0, 0, 0, 0, 0, 0, 0, -1.247366e-06, 
    0.0019411, 9.652421e-06, -1.148965e-08, -3.063192e-05, 0.002584964, 
    0.0008612595, 0, 0, 0.007723955, 0, 0.002461725, 0.01888097, 0.003070506, 
    0.003546441, 0.001886543,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.001900185, 0.0004054466, -0.0003147657, 0.0003601061,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.343349e-05, 
    -7.009164e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.005082101, 0.002319823, 
    6.657663e-07, 0.004712995, -2.191128e-09, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.001333778, 0.006819994, 0.0007283444, -1.152738e-05, 0.002159987, 
    0.000101119, 0.00205214, 0.0007272801, -4.481624e-06, 0.003899003, 
    0.0005379696, 0.002238383, 0.002639315, 0.01217104, 0.005446749, 
    0.0001734477, 0.002362532, 0.009646809, 0.00251194, 0.006982668, 
    0.000597153, 0.0001474927, -0.0001093591, 0.000341924, 0.00329614, 
    0.0001288525, 0.0007364712, 0.001375657, 0.0009722176,
  0.09261853, 0.07027228, 0.02008805, 0.02573128, 0.05506564, 0.02039831, 
    0.01592216, 0.04169425, 0.06396046, 0.05424792, 0.01558742, 0.01984121, 
    0.008722323, 0.01736752, 0.0374558, 0.005996791, 0.0259247, 0.03020831, 
    0.04040803, 0.05134102, 0.06693523, 0.02347602, 0.05043, 0.03720779, 
    0.03035246, 0.08436463, 0.0420392, 0.02488001, 0.05068971,
  0.1295635, 0.06057729, 0.08949104, 0.1448, 0.09015624, 0.09871041, 
    0.1459903, 0.07060906, 0.05306114, 0.06145236, 0.0764716, 0.03947056, 
    0.03778602, 0.1030413, 0.0664095, 0.09563506, 0.04670362, 0.0775272, 
    0.07593452, 0.110341, 0.1256964, 0.1024633, 0.07017322, 0.01241658, 
    0.07681831, 0.07528166, 0.0537467, 0.1440451, 0.1421998,
  0.007704683, 0.02180598, 0.1039645, 0.05623059, 0.1052455, 0.1101024, 
    0.1796323, 0.0897026, 0.06855017, 0.08465275, 0.1800816, 0.08905288, 
    0.04709731, 0.1479441, 0.09798307, 0.07119209, 0.1591458, 0.2190967, 
    0.1618171, 0.1357055, 0.1776306, 0.08778794, 0.01652968, 0.0339994, 
    0.04801542, 0.05155944, 0.1705709, 0.1148093, 0.04807729,
  -5.966932e-07, 0.08222848, 0.04042024, 0.005574928, 0.1691927, 0.01599616, 
    0.04204609, 0.01835646, 0.1812061, 0.02694, 0.1513724, 0.02225732, 
    0.006484168, 0.0598126, 0.1330767, 0.1728571, 0.08792947, 0.1260384, 
    0.06867414, 0.07326124, 0.004175543, 8.64656e-05, 0.005970604, 
    0.03015301, 0.1064103, 0.1911451, 0.1022399, 0.03079532, 2.406234e-05,
  0.001956608, 0.06348445, 0.2606071, 0.1673709, 0.1019915, 0.06713378, 
    0.126711, 0.1151508, 0.2122619, 0.01503027, 0.03591328, 0.1675414, 
    0.02602078, 0.03144624, 0.01557163, 0.1013428, 0.09530567, 0.09044696, 
    0.06883945, -0.000707276, -6.035412e-05, 0.00393768, 0.008259444, 
    0.3105042, 0.3154652, 0.2879836, 0.07919062, 0.00364824, 8.342519e-05,
  0.000729915, 0.1307944, 0.1667675, 0.059967, 0.00693243, 0.03160059, 
    0.105095, 0.1425978, 0.1985882, 0.2929212, 0.04465896, 0.09536701, 
    0.1088342, 0.08880446, 0.07645731, 0.03037405, 0.007185667, 0.04159878, 
    0.0005866715, 0.01694337, 0.0005686359, 0.008570691, 0.01928789, 
    0.3035261, 0.1469174, 0.0453576, 0.05707644, 0.008113433, 0.002387338,
  8.515729e-06, 0.0003499339, 2.035562e-05, 4.651984e-05, 2.551018e-06, 
    -2.59902e-05, 0.01508558, 0.08871152, 0.02501645, 0.02342979, 0.0745856, 
    0.03884133, 0.05863268, 0.02268575, 0.005705706, 0.04806773, 0.01833505, 
    0.02414736, 0.03780567, 0.07868306, 0.05348271, 0.002821939, 0.00386054, 
    1.824361e-05, 0.0002781115, 9.744315e-05, -0.0003716199, 0.01893876, 
    0.01667673,
  0.08861357, 0.008003902, 1.840592e-05, 8.77077e-06, 2.271573e-06, 
    -1.0608e-08, -3.998825e-08, -0.0003893641, 0.0001166682, 0.0009362079, 
    0.003465074, 0.01713845, 0.001005401, 0.000336492, 0.01121859, 
    -7.314205e-05, 0.04334005, 0.07303848, 0.1455391, 0.1395438, 0.2371623, 
    0.05283152, 0.001348225, 0.001145819, 0.01533762, 0.02190769, 
    0.005455059, 0.005047487, 0.08154844,
  0.003024929, -0.0006958433, 0.009272939, 7.627672e-05, 0.003610233, 
    -1.856256e-05, 1.433496e-05, 0, 0.000669309, 0.07714686, 0.09441894, 
    0.09619146, 0.06755748, 0.08219893, 0.0518849, 0.02165837, 0.08424595, 
    0.08389654, 0.06137365, 0.04637014, 0.0342483, 0.1408544, 0.1092086, 
    0.1322186, 0.1724413, 0.1490689, 0.05374636, 0.01109355, -0.0003170852,
  0.0001434083, 0, 2.183423e-06, -1.091027e-09, 0.006731443, -4.094127e-06, 
    2.013024e-05, 0, -9.925268e-06, 0, 0.002559216, 0.0001018472, 0.0186756, 
    0.03367006, 0.02489715, 0.02669748, 0.04834674, 0.0300466, 0.01843396, 
    0.003088239, 0, 0.0286331, 0.05071215, 0.07541571, 0.05318831, 0.1021552, 
    0.02433546, 0.01895208, 0.001916188,
  0.007812834, 1.741212e-07, 0.001558282, 0, 0, 0.000486283, -2.175424e-06, 
    0, 0, 0, 0, 0, 0, -0.000113209, 0.006726997, 0.006327717, 0.001198724, 
    0.0003129331, 0.01027991, 0.0008934521, -4.190249e-05, -4.113371e-05, 
    0.01161701, 0, 0.009155825, 0.03412036, 0.01473124, 0.01544536, 0.01285785,
  -0.0001151537, 0, 0, 0, 0, -1.681652e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.004054538, 0.003374678, 0.003922597, 0.001267447,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3.134092e-05, 
    -1.530855e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -3.77987e-05, -7.577186e-09, 0, -2.328643e-06, 
    0.0006884785, 0.007194984, 0.005923891, -4.201184e-05, 0.005117086, 
    -0.000152172, -0.0001307096, -0.0002328124, 0, 4.970401e-07, 
    -1.911106e-05, 0, 0, 0.0003013099, -1.978528e-05, 0,
  0.01054377, 0.01255133, 0.01053421, 2.517866e-05, 0.00436506, 0.007255782, 
    0.01531883, 0.01088549, 0.006088921, 0.02743909, 0.03725724, 0.02152634, 
    0.02734052, 0.06442815, 0.072518, 0.03802558, 0.01884076, 0.02142785, 
    0.01220437, 0.03489451, 0.02250835, 0.01043821, 0.004533296, 0.004507254, 
    0.0255445, 0.03113951, 0.02342223, 0.0244144, 0.011841,
  0.1361732, 0.1189898, 0.09589224, 0.1520857, 0.1445363, 0.1450878, 
    0.1112693, 0.1018277, 0.118005, 0.123562, 0.09723046, 0.07458951, 
    0.06211818, 0.0981006, 0.1022675, 0.03194462, 0.05362475, 0.07497526, 
    0.0933803, 0.09183243, 0.11341, 0.06315237, 0.09700496, 0.07029575, 
    0.1028281, 0.1677135, 0.1144333, 0.06233552, 0.115772,
  0.1547907, 0.09395837, 0.08629036, 0.1226222, 0.1087925, 0.09546483, 
    0.1160287, 0.08725016, 0.06910261, 0.07328502, 0.12225, 0.1179392, 
    0.1257501, 0.1418796, 0.1162303, 0.08674931, 0.08573281, 0.08234397, 
    0.08738571, 0.1111785, 0.1633949, 0.1338431, 0.09559842, 0.04216562, 
    0.08799436, 0.0838604, 0.04945497, 0.1309746, 0.1492285,
  0.008840998, 0.01573167, 0.1219013, 0.04803178, 0.08106605, 0.109358, 
    0.1599648, 0.09352575, 0.07038657, 0.0945301, 0.1965408, 0.08271087, 
    0.05079457, 0.1366613, 0.08021675, 0.04915352, 0.1502532, 0.2025601, 
    0.1394055, 0.1057375, 0.1666866, 0.09704401, 0.02005243, 0.01897644, 
    0.02851077, 0.04397813, 0.1578021, 0.1042332, 0.03833899,
  4.241255e-08, 0.07960749, 0.03191708, 0.004474858, 0.1584834, 0.01636583, 
    0.04050016, 0.01334617, 0.153863, 0.02963747, 0.148495, 0.01514613, 
    0.00665947, 0.04579335, 0.1211722, 0.1728979, 0.07945968, 0.1166061, 
    0.06900599, 0.04127178, 0.0002937, 0.0005218865, 4.484907e-06, 
    0.02283197, 0.08414207, 0.1690756, 0.07918119, 0.01359835, 1.214401e-06,
  0.0002051491, 0.07239349, 0.2472029, 0.1556077, 0.0763919, 0.06001025, 
    0.1146067, 0.1078687, 0.1884877, 0.01329613, 0.04457844, 0.1520925, 
    0.02130477, 0.02888901, 0.01914768, 0.1039008, 0.08980895, 0.08526254, 
    0.05203448, -0.0003004706, -1.038762e-05, 0.001609102, 0.001262747, 
    0.2911616, 0.2981136, 0.2516782, 0.06611884, 0.002319428, 0.0001268298,
  0.0005044658, 0.1189246, 0.1138945, 0.03656818, 0.003020549, 0.02866563, 
    0.06473482, 0.08794569, 0.1815598, 0.2566408, 0.03415915, 0.08102579, 
    0.1010631, 0.075409, 0.0625049, 0.02906073, 0.005701729, 0.03276236, 
    0.0002874228, 0.007698514, 0.001618469, 0.006944121, 0.01700483, 
    0.2136061, 0.1275916, 0.03457292, 0.036937, 0.006355955, 0.0008928952,
  -8.351429e-08, 1.723979e-05, 5.981846e-06, 7.006874e-06, -7.871337e-06, 
    -4.057891e-05, 0.009092314, 0.06921134, 0.03442682, 0.02724577, 
    0.05801972, 0.03551751, 0.04466055, 0.02321168, 0.002556034, 0.04762501, 
    0.02576163, 0.02437942, 0.0406552, 0.05680955, 0.04195246, 0.001871306, 
    4.423634e-05, 6.548819e-06, 7.193295e-05, 4.013887e-05, -3.367568e-05, 
    0.007551556, 0.01089135,
  0.08346448, 0.008942672, 2.051223e-06, 2.325721e-06, 1.552075e-06, 
    8.187888e-08, -9.222304e-07, -3.638643e-05, 3.371043e-05, 0.0005430349, 
    0.01026653, 0.01865957, 0.004147481, 0.0003919503, 0.009487135, 
    -3.698968e-05, 0.04513576, 0.05975069, 0.1314943, 0.1251025, 0.1616768, 
    0.02414301, 0.002213722, 0.0001569699, 0.009323921, 0.01267107, 
    0.002704563, 0.02582755, 0.06919952,
  0.05729013, 0.00737836, 0.01566676, 0.00473843, 0.0114663, 0.006666366, 
    0.009376157, 0, 0.003221741, 0.1732283, 0.1861654, 0.135499, 0.08939728, 
    0.1088004, 0.09788324, 0.1042359, 0.1242252, 0.08736724, 0.1532828, 
    0.1095914, 0.08359318, 0.1573022, 0.1592797, 0.142834, 0.1812814, 
    0.2026291, 0.1266774, 0.05576769, 0.08650527,
  0.05154253, 0.005957974, 0.002042636, 0.001064476, 0.03794205, 0.0353317, 
    0.0002009046, -1.228651e-05, -1.372239e-05, -7.122309e-09, 0.003433, 
    0.009708589, 0.05141761, 0.07738892, 0.07148259, 0.1041174, 0.1250321, 
    0.1487858, 0.1240833, 0.0066655, 0.0001959384, 0.04727053, 0.1146558, 
    0.1431006, 0.09421905, 0.254465, 0.1436114, 0.1153478, 0.07913662,
  0.02727652, -9.371149e-06, 0.01134877, 0, -7.920264e-05, 0.009254524, 
    0.003426773, 0, 0, 0, 0, 0, 0.0002974235, 0.003863036, 0.01990152, 
    0.01940816, 0.005472351, 0.01111115, 0.02492118, 0.003160358, 
    0.0002944495, 0.006429521, 0.02150915, 0.001199628, 0.01240629, 
    0.09327116, 0.1337689, 0.0633821, 0.03428813,
  -0.0002335157, 5.752026e-05, 0.0005112641, 0, 0.001371543, 0.0002728411, 0, 
    0, 0, 0, 0, 0, 0, -1.927545e-05, -6.548889e-05, -2.38921e-07, 0, 0, 0, 
    1.333508e-05, 0, -1.312821e-05, 0, 0, -2.495388e-05, 0.00488623, 
    0.009462967, 0.01510437, 0.009128491,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0002973057, 
    0.001911585, 0.0002226441, -2.254577e-05, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 5.628267e-06, 0, 0, -5.959131e-05, -9.356146e-06, 
    -2.028833e-08, 2.917859e-05, 0.005810048, 0.01520088, 0.01598867, 
    0.01815038, 0.00999971, 0.06203574, 0.02904853, 0.01833347, 0.008968187, 
    0.009015494, 0.0003445187, 0.002770289, -1.74143e-05, 0.0005219741, 
    0.001215248, -1.485607e-05,
  0.09162809, 0.04851909, 0.02972445, 0.03589598, 0.0314098, 0.0442394, 
    0.03016124, 0.04279868, 0.04720816, 0.07432658, 0.06705378, 0.107808, 
    0.1236393, 0.1534183, 0.160246, 0.1414033, 0.08708156, 0.1120904, 
    0.08587739, 0.08577283, 0.08712751, 0.07809675, 0.0927626, 0.07354038, 
    0.08161675, 0.09585706, 0.04532281, 0.03693885, 0.03637382,
  0.1595311, 0.1297658, 0.1501368, 0.1872026, 0.1892481, 0.1870304, 
    0.1517308, 0.1494137, 0.1326593, 0.1534155, 0.1395082, 0.1299876, 
    0.1368873, 0.1235585, 0.1158801, 0.04551412, 0.1036525, 0.1314643, 
    0.1258439, 0.1147462, 0.1475816, 0.1042824, 0.1420923, 0.1021801, 
    0.1356227, 0.2056028, 0.1633856, 0.06716803, 0.152956,
  0.1440908, 0.07717282, 0.07701971, 0.09692907, 0.1052276, 0.07265296, 
    0.09715687, 0.06903227, 0.05326509, 0.06552006, 0.1137329, 0.08898811, 
    0.109008, 0.1332597, 0.1155504, 0.0712136, 0.0993723, 0.06804539, 
    0.06680393, 0.1107819, 0.1564374, 0.1363711, 0.08937106, 0.06587878, 
    0.05860536, 0.08531082, 0.04582021, 0.117481, 0.1348534,
  0.009122218, 0.01261929, 0.08685956, 0.04218198, 0.05491088, 0.1202644, 
    0.1534769, 0.09325569, 0.05934308, 0.09511028, 0.1951783, 0.09486397, 
    0.04518882, 0.1303084, 0.06280199, 0.04022329, 0.1346549, 0.1981747, 
    0.1572939, 0.07798891, 0.1260181, 0.0724153, 0.008979359, 0.01702724, 
    0.02511027, 0.03063191, 0.1684556, 0.08715994, 0.03383205,
  -7.588152e-08, 0.07030655, 0.02578493, 0.003506229, 0.1481361, 0.01265012, 
    0.03863328, 0.009831387, 0.1315015, 0.01397675, 0.1409764, 0.006939468, 
    0.002138689, 0.03469658, 0.1093245, 0.1570253, 0.07015471, 0.1005531, 
    0.07004076, 0.03314076, 0.00460227, 0.001682524, 2.996887e-05, 
    0.02005554, 0.09451938, 0.1674943, 0.07201348, 0.002537799, 1.5363e-06,
  7.693829e-05, 0.09738703, 0.2342358, 0.1321048, 0.063928, 0.04940997, 
    0.09720431, 0.09535098, 0.1504441, 0.01084356, 0.04504543, 0.1270092, 
    0.01554773, 0.02181588, 0.01954526, 0.09343784, 0.0827406, 0.07262764, 
    0.03943192, 0.0002237431, 2.542544e-05, -7.768527e-05, 0.0001336918, 
    0.2414922, 0.2698641, 0.2039098, 0.06000005, 0.001752942, 0.0001335394,
  0.0003606769, 0.09918008, 0.08183313, 0.02736733, 0.005660782, 0.02630974, 
    0.04400714, 0.07488874, 0.1616303, 0.2141074, 0.03021154, 0.06679806, 
    0.08264195, 0.05305695, 0.04796904, 0.03125319, 0.005560043, 0.01707173, 
    0.0006038492, 0.006632096, 0.00381979, 0.007419873, 0.02112412, 
    0.1479711, 0.1189493, 0.03096403, 0.02284043, 0.005798942, 0.0004593242,
  2.199733e-06, 7.492208e-06, 2.049346e-06, 3.082477e-06, -1.020562e-06, 
    -1.475553e-05, 0.004659412, 0.06483602, 0.02932482, 0.02534513, 
    0.05662676, 0.03452456, 0.03406054, 0.01998422, 0.003281748, 0.04147898, 
    0.02536513, 0.03815126, 0.05681975, 0.04534635, 0.03236067, 0.001081859, 
    7.542834e-05, 3.81739e-06, 0.0003284287, 0.005484198, 2.344587e-06, 
    0.03000265, 0.006948249,
  0.05429136, 0.008553312, 5.178119e-07, 5.679248e-07, 1.322345e-06, 
    -2.900416e-08, -3.53595e-06, 6.554386e-05, 0.0002279576, 0.0005699193, 
    0.01184871, 0.0305035, 0.01251931, 0.0001991528, 0.003457064, 
    7.343165e-05, 0.05202623, 0.05264796, 0.1202688, 0.08450023, 0.1241612, 
    0.009493185, 0.0018652, 0.0001239728, 0.0008678613, 0.007647097, 
    0.003221781, 0.02052677, 0.05969771,
  0.07787439, 0.02656502, 0.01881054, 0.008966393, 0.01647023, 0.01415056, 
    0.01970033, -5.870282e-05, 0.007834687, 0.22575, 0.2132199, 0.1328603, 
    0.0767718, 0.09406277, 0.102816, 0.1083308, 0.1002186, 0.08670397, 
    0.1135185, 0.07890947, 0.1237865, 0.1412606, 0.1515256, 0.1354438, 
    0.1553885, 0.1611582, 0.09943507, 0.05357489, 0.07456514,
  0.09258075, 0.05698989, 0.0412509, 0.00538319, 0.07621567, 0.09432444, 
    0.002931464, 0.01546633, 0.0005847987, -2.927639e-05, 0.01714369, 
    0.04455334, 0.1090947, 0.1380873, 0.14926, 0.1723674, 0.2075424, 
    0.2669199, 0.2108119, 0.08032437, 0.002839569, 0.100205, 0.187679, 
    0.1998441, 0.1428527, 0.3025054, 0.1662962, 0.1448931, 0.1379015,
  0.1886636, 0.0665381, 0.02667261, 0.006961029, 0.003868421, 0.04722891, 
    0.01164646, 0, 0, 0, 0, 0, 0.006174964, 0.02429248, 0.05086676, 
    0.06604834, 0.05246081, 0.05925252, 0.07087403, 0.0119523, 0.000529122, 
    0.01502049, 0.05225613, 0.02840759, 0.03738954, 0.2233134, 0.2211998, 
    0.1475729, 0.1645571,
  0.07055132, 0.001473007, 0.009209073, 4.788928e-05, 0.002465428, 
    0.00356931, -8.499858e-05, 1.009352e-05, 0, 0, 0, 0, 0, 0.01172244, 
    0.01475889, 0.003217363, 0.004045772, -1.984056e-06, 0, 0.001708568, 
    -0.0001595321, 0.001293514, 0, -2.752174e-05, 0.004805361, 0.02256662, 
    0.07221226, 0.1004751, 0.08964948,
  -8.857766e-07, 0, -4.325601e-05, 0.0003561744, 0.002776852, 4.773053e-05, 
    0, 0, 0, 0.000164203, 0, 0, 0.0003898411, 0.002587389, 4.805306e-06, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.103471e-06, 0.006984655, -4.715697e-06,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.109561e-07, -0.0005349985, 
    0.005563525, 0.007676336, 0.002057848, -0.0001594036, 0, 0.0005068555, 
    0.0002336695, 0, 0, 0, 0.0001051321, 0,
  0, 0, -6.565633e-07, 0.0005198282, 0, 0, 0.007215379, 0, -0.00018208, 
    -0.000599506, -1.420827e-05, -0.0001177481, 0.001662754, 0.07122345, 
    0.06538624, 0.05472649, 0.04993953, 0.1019207, 0.08773462, 0.06367716, 
    0.05423563, 0.06390901, 0.07500461, 0.02905913, 0.04090725, 0.018261, 
    0.01917916, 0.01532115, 0.0002973862,
  0.1268365, 0.07831793, 0.05228009, 0.05932375, 0.06306335, 0.0859572, 
    0.1060404, 0.1424673, 0.1500459, 0.1283512, 0.1143722, 0.2064547, 
    0.2186844, 0.2202814, 0.1852479, 0.165001, 0.1578566, 0.1599836, 
    0.1308988, 0.1479383, 0.1410263, 0.1476358, 0.1607736, 0.147844, 
    0.1553178, 0.1736861, 0.1426691, 0.1242725, 0.1074402,
  0.1620168, 0.1434729, 0.1562103, 0.1949476, 0.1968782, 0.1815207, 0.158781, 
    0.1405306, 0.142336, 0.1616894, 0.1520293, 0.1574547, 0.1514853, 
    0.1239302, 0.1277829, 0.06280583, 0.1002514, 0.1453532, 0.1458263, 
    0.150849, 0.15266, 0.1041977, 0.1517238, 0.1474717, 0.1298658, 0.2130566, 
    0.1655955, 0.07270782, 0.1494038,
  0.1367621, 0.07218526, 0.062378, 0.083888, 0.0947312, 0.05849976, 0.10767, 
    0.08986481, 0.05315868, 0.05670121, 0.1026148, 0.07879502, 0.104118, 
    0.1363961, 0.09616677, 0.07019823, 0.1133835, 0.05064476, 0.06319734, 
    0.0986582, 0.1367133, 0.1187746, 0.08376507, 0.07652074, 0.04772423, 
    0.0750219, 0.03976529, 0.1105671, 0.1337577,
  0.009523837, 0.008833677, 0.05307214, 0.03668455, 0.03903632, 0.1028054, 
    0.1517102, 0.06586071, 0.06086651, 0.0949514, 0.198134, 0.101285, 
    0.03923753, 0.1260862, 0.0547933, 0.03754782, 0.1159157, 0.2057553, 
    0.177069, 0.06669523, 0.1125629, 0.04351759, 0.004257297, 0.003052169, 
    0.02822731, 0.02635237, 0.1512118, 0.09016486, 0.03118876,
  -5.949903e-10, 0.06940407, 0.01768701, 0.00230369, 0.1394733, 0.008060592, 
    0.04047447, 0.00813218, 0.09297605, 0.01074633, 0.1224659, 0.003559606, 
    0.0004248744, 0.02750932, 0.0877833, 0.1483905, 0.06299522, 0.0868787, 
    0.0626104, 0.02297106, 0.013724, 1.192663e-06, 0.0001186268, 0.01552612, 
    0.1015508, 0.1499557, 0.06087128, 0.0001311574, 2.079118e-06,
  0.001682134, 0.09400956, 0.2329773, 0.1250221, 0.06207051, 0.03343629, 
    0.07297256, 0.0688051, 0.1167971, 0.007975833, 0.04728494, 0.08587511, 
    0.01139716, 0.0161106, 0.01344847, 0.08134638, 0.07033496, 0.05408608, 
    0.03067495, 0.0002891175, 1.783075e-05, -0.000644512, 1.469875e-05, 
    0.2061833, 0.2371191, 0.1482999, 0.05652446, 0.001372939, 0.0002296514,
  0.0006736213, 0.07524328, 0.05997291, 0.01791, 0.00654248, 0.02062444, 
    0.02179126, 0.05808856, 0.1457324, 0.1842661, 0.02445213, 0.04651667, 
    0.0686147, 0.03962412, 0.02387453, 0.03021501, 0.003575519, 0.006445933, 
    0.0006758365, 0.006351107, 0.001632705, 0.007765623, 0.0417325, 
    0.1148894, 0.0942249, 0.02855527, 0.01682642, 0.005444942, 0.000640548,
  2.484944e-05, 2.680807e-06, 5.754569e-07, 1.316349e-06, 4.455035e-06, 
    -1.177437e-05, 0.002863123, 0.05714488, 0.03440544, 0.02665237, 
    0.0541922, 0.02829709, 0.02639625, 0.03306222, 0.004286089, 0.02799166, 
    0.02529964, 0.03656905, 0.07992828, 0.04225424, 0.02342299, 0.001026138, 
    4.448961e-05, 1.294885e-05, 0.0006495361, 4.23053e-05, -5.886036e-06, 
    0.04504821, 0.00978163,
  0.04362016, 0.002378343, 6.247969e-08, 2.274882e-07, 2.157219e-06, 
    -8.718424e-08, 6.762809e-05, 0.0005657263, 0.002123693, 0.002965989, 
    0.01993552, 0.02986786, 0.01260329, 9.71501e-05, 7.788648e-05, 
    5.046323e-05, 0.03638427, 0.02299756, 0.09616529, 0.08487108, 0.1039796, 
    0.003688244, 0.002966262, 2.82073e-05, 0.0001540481, 0.02013953, 
    0.01054394, 0.008084993, 0.04272924,
  0.05521829, 0.02757932, 0.01348415, 0.01261382, 0.01963044, 0.01079822, 
    0.02136595, 2.687205e-06, 0.0153564, 0.2284162, 0.2030903, 0.1174288, 
    0.06705164, 0.08923162, 0.1028987, 0.08995937, 0.08460761, 0.08450451, 
    0.06991053, 0.06139408, 0.09535451, 0.1040189, 0.1143641, 0.1166374, 
    0.1157248, 0.1183204, 0.04843853, 0.05198862, 0.0436422,
  0.07501687, 0.05313412, 0.07608466, 0.0221469, 0.1484589, 0.1254316, 
    0.01401683, 0.1254532, 0.03965753, 0.002699401, 0.06669912, 0.121803, 
    0.1645585, 0.1640262, 0.1621191, 0.174246, 0.2169179, 0.2551647, 
    0.2122984, 0.1637589, 0.02824613, 0.1621215, 0.1887626, 0.2122417, 
    0.1560447, 0.3012254, 0.154422, 0.1461938, 0.1370149,
  0.1848248, 0.1344489, 0.10319, 0.05232534, 0.07097515, 0.09496713, 
    0.0763658, -0.0001251582, -1.042739e-05, 0, 0, -0.0001868402, 0.01702832, 
    0.07069025, 0.07197998, 0.09913173, 0.08614817, 0.1092479, 0.1752295, 
    0.04455892, 0.02295459, 0.1201785, 0.1685383, 0.04070227, 0.09349455, 
    0.2343356, 0.2315927, 0.1495, 0.188728,
  0.2236471, 0.08250702, 0.0733854, 0.1045567, 0.07322922, 0.03553927, 
    0.02603316, 0.02313406, 0.002700355, 0.0001844383, -3.116584e-06, 0, 
    -0.0006030213, 0.02945713, 0.0192969, 0.02104197, 0.0169631, 0.02502345, 
    -1.719493e-05, 0.01301679, 0.007563121, 0.02756838, 0.02270176, 
    0.02064118, 0.03469797, 0.03742076, 0.145394, 0.2045876, 0.2222195,
  0.01415304, 0.0121376, 0.002816386, 0.02572886, 0.03744284, 0.03283599, 
    0.0006934325, 0.008904354, 0.004335454, 0.009549985, 0.001878318, 
    0.006145351, 0.009565561, 0.009220291, 0.001473513, 0.003742177, 
    -9.100726e-05, 0.003457833, 0.0004508143, 0.001081874, -9.808647e-07, 0, 
    0, 0, 0.0002730702, -2.620036e-05, -9.962131e-06, 0.0205836, 0.01132727,
  0, -1.367022e-08, 0, -5.493536e-05, 0.005416658, 0.005485533, 0.000855128, 
    5.566158e-07, -1.595216e-05, -3.775807e-06, 2.447483e-05, 0.0008799206, 
    0.002366296, 0.00289181, 0.002189178, 0.002955036, 0.001029831, 
    3.371897e-06, -4.209764e-07, 0, 0, 0, 0, 0, 0, 0, 0, -6.60419e-08, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -4.972138e-07, 0, -0.0004186435, 
    0.007416308, 0.01545327, 0.0150112, 0.01214856, 0.001490397, 
    -0.0001252976, 0.00269403, 0.01335828, 0.002333659, -0.0009459196, 
    -4.213156e-07, 0.0008383312, 0.0001500256,
  0.03631589, 0.004429294, 0.0578675, 0.02328676, -0.0006644217, 
    -0.0007522067, 0.02382023, -3.885572e-05, -0.0003619998, 0.0005127808, 
    -0.0003803931, 0.0009929343, 0.04283682, 0.1608125, 0.1561727, 0.1481695, 
    0.1647275, 0.1984081, 0.1535047, 0.161489, 0.116374, 0.1278917, 
    0.1101249, 0.1366499, 0.2308004, 0.1309754, 0.1521754, 0.2026181, 0.10896,
  0.1734954, 0.1211342, 0.1182264, 0.1162341, 0.1214621, 0.1513876, 0.14957, 
    0.1973278, 0.1722647, 0.1549687, 0.1838967, 0.2814431, 0.248221, 
    0.2193399, 0.1864432, 0.1920739, 0.1692777, 0.1546307, 0.1618389, 
    0.1639542, 0.1926977, 0.2112488, 0.2051269, 0.1824289, 0.1964273, 
    0.2112918, 0.1699804, 0.1586948, 0.1622759,
  0.152193, 0.1525524, 0.1460565, 0.2059664, 0.2162959, 0.1812015, 0.1578589, 
    0.1467829, 0.1531126, 0.1548418, 0.140362, 0.1553009, 0.1656684, 
    0.1261743, 0.1211912, 0.06316893, 0.09782496, 0.143487, 0.1383937, 
    0.1614525, 0.1441626, 0.1056625, 0.1742298, 0.1667749, 0.1327849, 
    0.2117072, 0.1473373, 0.08164325, 0.1507258,
  0.1322736, 0.07715711, 0.05946827, 0.07964066, 0.08713371, 0.05866279, 
    0.1096393, 0.08318871, 0.04602249, 0.04780303, 0.1091064, 0.08041574, 
    0.09895632, 0.1400592, 0.083519, 0.05447828, 0.09454538, 0.05788369, 
    0.04618646, 0.08931664, 0.1284852, 0.1028943, 0.0984512, 0.04380945, 
    0.04752539, 0.0687369, 0.03503748, 0.1092085, 0.1393141,
  0.008626875, 0.005876921, 0.03819688, 0.0331878, 0.03277786, 0.1058448, 
    0.1148535, 0.06897411, 0.07337353, 0.07913864, 0.154644, 0.1022431, 
    0.04488682, 0.1171267, 0.04586993, 0.02984924, 0.08226456, 0.1801664, 
    0.1737457, 0.06730147, 0.09497833, 0.0267437, 0.001863359, 0.0006716725, 
    0.03277329, 0.01501093, 0.1314203, 0.08478399, 0.02625286,
  6.011414e-09, 0.06479003, 0.006564463, 0.001816932, 0.123307, 0.005387727, 
    0.03708375, 0.009749335, 0.07234367, 0.02877181, 0.09091415, 0.002957781, 
    0.001890322, 0.02320034, 0.06494261, 0.1545239, 0.05019879, 0.08115284, 
    0.06112469, 0.0164391, 0.002952403, 4.656896e-07, 4.274412e-05, 
    0.009419207, 0.09296567, 0.1208783, 0.0687094, 0.0005727626, 8.573617e-07,
  0.0002293692, 0.1246732, 0.2079934, 0.08858129, 0.06411942, 0.02755201, 
    0.05850511, 0.05167063, 0.09929649, 0.006255745, 0.05889004, 0.06762954, 
    0.01349925, 0.01319207, 0.01144474, 0.06360203, 0.06879136, 0.05330161, 
    0.02541198, 0.0001495376, -1.371184e-05, -0.0004096796, -2.969009e-05, 
    0.1825071, 0.2283136, 0.106507, 0.04573057, 0.001221676, 0.0002585946,
  0.001817882, 0.06309301, 0.04655583, 0.01462017, 0.002104179, 0.01627543, 
    0.01095106, 0.0394878, 0.1273135, 0.1526067, 0.02183871, 0.03321988, 
    0.06611506, 0.035614, 0.0106779, 0.03549957, 0.004695519, 0.01118526, 
    0.001015456, 0.002000686, 0.002872381, 0.005024645, 0.0355735, 
    0.08434585, 0.0977485, 0.0354988, 0.01060645, 0.004374909, 0.0006144797,
  0.0005692743, 1.082024e-06, 2.882619e-07, 9.975887e-07, 1.080378e-07, 
    -1.329724e-05, 0.001852406, 0.05754071, 0.03207348, 0.04039254, 
    0.05426772, 0.02553031, 0.01863056, 0.0396203, 0.002499539, 0.02223078, 
    0.03547567, 0.03563303, 0.09816451, 0.04469281, 0.017062, 0.0005545422, 
    6.551221e-05, 5.193441e-06, 0.0007078608, 1.402878e-06, 5.045803e-07, 
    0.06114135, 0.007901697,
  0.03953215, 3.026056e-05, 4.945351e-09, -4.710716e-09, 2.813854e-06, 
    2.385926e-08, 0.0004610183, 0.0001667979, 1.237578e-05, 0.002767218, 
    0.02603759, 0.02665519, 0.002313704, 0.0002990958, 1.664293e-05, 
    1.982586e-05, 0.02735138, 0.01442186, 0.0737403, 0.07074179, 0.07622916, 
    0.002533933, 0.00347999, 8.224139e-05, 0.000299672, 0.01022128, 
    0.01155075, -3.353785e-05, 0.03533639,
  0.038446, 0.02471596, 0.01179261, 0.01053366, 0.02078023, 0.00818091, 
    0.02387451, 0.001751564, 0.0433625, 0.2146974, 0.187594, 0.1099568, 
    0.06994539, 0.09490994, 0.08073776, 0.06894644, 0.07133101, 0.05014944, 
    0.05136993, 0.05446025, 0.07115572, 0.07668946, 0.1025742, 0.1026429, 
    0.09578437, 0.07818113, 0.03615178, 0.05057731, 0.02990649,
  0.04848887, 0.05192518, 0.09513637, 0.05893246, 0.1659243, 0.1451975, 
    0.04480233, 0.1760332, 0.1217687, 0.06150063, 0.1038482, 0.1318905, 
    0.1863395, 0.1734594, 0.1750721, 0.1507932, 0.2259774, 0.2392806, 
    0.216362, 0.1509636, 0.08640275, 0.190291, 0.1832579, 0.2108255, 
    0.1670917, 0.3016, 0.1400142, 0.1252614, 0.1240167,
  0.1750822, 0.1244585, 0.1726193, 0.1647131, 0.1883982, 0.1684177, 
    0.1586929, 0.002834307, -0.0001625301, 0.0001393329, 7.632592e-05, 
    0.01164004, 0.04445042, 0.08737356, 0.1069083, 0.1208638, 0.1472922, 
    0.1607531, 0.2082061, 0.09379404, 0.07878891, 0.1660618, 0.1743592, 
    0.08541695, 0.1202189, 0.2316342, 0.2289313, 0.1461034, 0.1871367,
  0.2520818, 0.1802518, 0.1368213, 0.1650911, 0.1763639, 0.1580894, 
    0.08722843, 0.06391622, 0.01425949, 0.02957608, 0.01376941, 
    -0.0002077517, 0.02604698, 0.0525474, 0.06994533, 0.05691708, 0.04564493, 
    0.0810907, 0.03737903, 0.09137531, 0.04544736, 0.1008084, 0.09165485, 
    0.05154728, 0.07876992, 0.05558737, 0.1467859, 0.2588074, 0.2489607,
  0.1035054, 0.1030702, 0.09487373, 0.09868694, 0.1117982, 0.09876538, 
    0.05446194, 0.04584074, 0.02354377, 0.05351913, 0.04250415, 0.0397755, 
    0.01546946, 0.01702213, 0.03955706, 0.03847516, 0.01943398, 0.02112254, 
    0.04899087, 0.02223059, 0.0110043, 0.0003819202, 1.056339e-06, 0, 
    0.04125594, 0.0003169793, -4.704254e-06, 0.0641026, 0.07933919,
  0.03592335, 0.02829186, 0.02594912, 0.05187328, 0.03750421, 0.009487191, 
    0.001673497, -0.0001449748, 0.003030723, 0.01239593, 0.01386914, 
    0.02186263, 0.01843769, 0.01324108, 0.02097016, 0.04037658, 0.05863695, 
    0.03228422, 0.01156769, -8.901126e-05, 0, 0, 0, -5.860018e-05, 
    -0.0006300208, 4.353211e-05, -4.122499e-06, -0.008222936, 0.04110883,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.845309e-06, 0.004904991, 
    0.01648903, 0.1249077, 0.07936574, 0.02997178, 0.03190847, 0.01633864, 
    -0.0009101309, 0.009730941, 0.02646612, 0.03263073, 0.03521268, 
    0.08191504, 0.005431994, 0.0008995752,
  0.053935, 0.024503, 0.1262007, 0.07177985, -0.001497462, -5.245718e-05, 
    0.06704126, -0.002416088, 0.001206026, 0.004147786, 0.007697622, 
    0.009946799, 0.09910651, 0.2094031, 0.1832929, 0.1858729, 0.2527196, 
    0.3113391, 0.1868379, 0.2196107, 0.1988663, 0.1974441, 0.215195, 
    0.2258787, 0.3848273, 0.2579023, 0.2694056, 0.3094664, 0.1759887,
  0.2462845, 0.1464034, 0.1772246, 0.1700211, 0.1761357, 0.227033, 0.1713442, 
    0.2368707, 0.2224715, 0.226159, 0.2267686, 0.3178732, 0.2651521, 
    0.2373053, 0.1891186, 0.1804682, 0.1684377, 0.1478282, 0.2233281, 
    0.2182846, 0.2147931, 0.259529, 0.2579094, 0.2256453, 0.2717795, 
    0.2523753, 0.2202484, 0.1868045, 0.1766297,
  0.1386846, 0.1558774, 0.1398616, 0.2173966, 0.2088225, 0.1754605, 
    0.1431328, 0.1466053, 0.154438, 0.1533356, 0.1448701, 0.166902, 0.189039, 
    0.1234048, 0.1155957, 0.05465302, 0.09151206, 0.1314822, 0.1376742, 
    0.1808929, 0.157659, 0.1004667, 0.2016308, 0.1727165, 0.121345, 0.182058, 
    0.1397965, 0.09716867, 0.1455659,
  0.1168215, 0.08333548, 0.04382545, 0.0741405, 0.08002009, 0.04425626, 
    0.101578, 0.05213257, 0.03584544, 0.04168148, 0.09178474, 0.06217274, 
    0.1047171, 0.1348003, 0.0672525, 0.03623179, 0.08830626, 0.0590794, 
    0.05594856, 0.06605384, 0.116532, 0.1047475, 0.0931837, 0.0384398, 
    0.04989123, 0.05530075, 0.03602108, 0.1142187, 0.1219706,
  0.01075177, 0.001156882, 0.02644739, 0.02622552, 0.03294556, 0.1032638, 
    0.08799292, 0.0687844, 0.08336724, 0.06428077, 0.1487866, 0.11729, 
    0.05273073, 0.1274143, 0.04374896, 0.004345914, 0.06758384, 0.1749714, 
    0.1486541, 0.07277001, 0.07606709, 0.03322455, 0.006832967, 5.161534e-05, 
    0.02988628, 0.009400578, 0.121339, 0.07629906, 0.02870824,
  1.013098e-05, 0.05677976, 0.002489528, 0.001648, 0.1136352, 0.004619107, 
    0.03108581, 0.02198697, 0.05196208, 0.01463563, 0.08202057, 0.004854649, 
    0.001050988, 0.02391938, 0.04482662, 0.1445629, 0.04860046, 0.07132596, 
    0.06158882, 0.01920598, 0.001110549, -6.446497e-07, -4.616557e-06, 
    0.005470765, 0.08082393, 0.1051018, 0.07181823, 0.009439106, 2.039716e-07,
  0.00363825, 0.1216577, 0.1945952, 0.07410535, 0.05702522, 0.02848034, 
    0.05715698, 0.04804237, 0.09059292, 0.005936549, 0.06005442, 0.06033149, 
    0.01269981, 0.01153977, 0.01216629, 0.05419279, 0.05428352, 0.04953753, 
    0.02092628, 9.587045e-05, -4.13791e-05, -0.0003408287, -3.934893e-05, 
    0.1871348, 0.2068211, 0.08119836, 0.02448628, 0.00102376, 0.0002732271,
  0.009005216, 0.05306378, 0.04400095, 0.01058707, 0.001275435, 0.01069694, 
    0.005982571, 0.02151329, 0.09646358, 0.1448858, 0.03477431, 0.01986685, 
    0.06319486, 0.03578547, 0.008811668, 0.03942883, 0.006281834, 
    0.005073812, 0.001210565, 0.002056457, 0.01066677, 0.002179612, 
    0.03687448, 0.06445298, 0.1140618, 0.04541909, 0.01050939, 0.005661725, 
    0.001914268,
  0.0001403677, 1.346327e-06, -1.102652e-05, 5.273083e-07, 4.940157e-05, 
    1.026157e-05, 0.002140725, 0.05545232, 0.03505911, 0.0390629, 0.05096358, 
    0.03313948, 0.01536227, 0.03051405, 0.008608162, 0.02507954, 0.04279531, 
    0.03579579, 0.1097466, 0.06217054, 0.01886719, 0.001047918, 4.132932e-05, 
    1.296701e-05, 0.0006353027, 3.179476e-06, -1.789287e-05, 0.02510873, 
    0.005433939,
  0.02111534, -1.491347e-06, 4.317375e-08, 9.117634e-07, 1.203478e-06, 
    2.202373e-09, 0.0003171983, 5.027501e-05, 1.006708e-05, 0.001620309, 
    0.01594759, 0.0249849, 0.0009137575, 0.005090741, 6.287601e-06, 
    2.83739e-06, 0.02238215, 0.002716957, 0.06817935, 0.05602272, 0.05266815, 
    0.002459623, 0.004234502, -7.597644e-05, 0.0001842693, 0.0007835591, 
    0.01362905, -2.480929e-06, 0.02142958,
  0.02807442, 0.01261162, 0.00769984, 0.006005406, 0.03231307, 0.009100826, 
    0.02405463, 0.003650774, 0.08738896, 0.212586, 0.1754317, 0.1072564, 
    0.09160227, 0.09576324, 0.0629442, 0.05517181, 0.06049274, 0.04217957, 
    0.05916586, 0.04732001, 0.05187383, 0.06478389, 0.09087403, 0.08460858, 
    0.08728186, 0.05555411, 0.03589042, 0.0493366, 0.02628459,
  0.02939791, 0.05077996, 0.1046012, 0.1075993, 0.1616559, 0.1299294, 
    0.1092963, 0.1723308, 0.1295056, 0.1104522, 0.1263776, 0.1065369, 
    0.1778825, 0.1644703, 0.1683385, 0.1488233, 0.2236244, 0.2373667, 
    0.2162331, 0.152789, 0.1147458, 0.1906211, 0.1699015, 0.2147636, 
    0.1800365, 0.2832814, 0.1179587, 0.1206341, 0.08264139,
  0.1734837, 0.1692704, 0.1927686, 0.1732839, 0.1800114, 0.1741965, 
    0.2295816, 0.03906786, 0.01411073, 0.02363323, 0.004768687, 0.02545786, 
    0.06601593, 0.1109786, 0.1634167, 0.1521269, 0.193552, 0.2014836, 
    0.2843984, 0.1488608, 0.1722848, 0.1778128, 0.164958, 0.1086359, 
    0.1400988, 0.2257935, 0.2296447, 0.1498892, 0.1724285,
  0.2668476, 0.2415635, 0.1620299, 0.2082049, 0.2095967, 0.1899126, 0.178465, 
    0.1447314, 0.1246786, 0.08619472, 0.04391237, 0.01232872, 0.04524069, 
    0.1160497, 0.1427963, 0.1212233, 0.08091932, 0.1655044, 0.1005654, 
    0.1804566, 0.1127168, 0.1068525, 0.1289733, 0.09207607, 0.1236528, 
    0.0988685, 0.1848625, 0.2795263, 0.2478672,
  0.1263942, 0.1448808, 0.135179, 0.1497413, 0.1440646, 0.1266254, 0.119293, 
    0.09570803, 0.06191124, 0.0988678, 0.07722793, 0.05771567, 0.06321276, 
    0.1130498, 0.07237422, 0.1126071, 0.03677557, 0.05709708, 0.05056011, 
    0.0899232, 0.04819961, 0.01490784, 0.000159785, -2.519565e-05, 
    0.07699014, 0.003708216, 0.002309317, 0.1037147, 0.1160702,
  0.07053594, 0.07224813, 0.04568749, 0.05700543, 0.04450022, 0.01872399, 
    0.02017697, 0.01052555, 0.008911035, 0.02330993, 0.02719059, 0.02624199, 
    0.02637007, 0.08876489, 0.1298948, 0.1387284, 0.1642797, 0.1804072, 
    0.1063293, 0.05185395, 0.009154158, 0.009696773, -6.518014e-05, 
    -0.002770687, 0.0143023, -0.0001248134, -0.0047064, 0.04667779, 0.07546994,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  -0.001269084, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0325904, 0.05471871, 
    0.1069118, 0.1915177, 0.2501342, 0.105567, 0.03630913, 0.02646646, 
    0.006982566, 0.02254699, 0.1942772, 0.2219457, 0.2490025, 0.3248174, 
    0.07715755, 0.008866895,
  0.108266, 0.124116, 0.3161928, 0.191208, 0.004496641, 0.004366315, 
    0.140945, 0.01691477, 0.01260325, 0.02366883, 0.03939407, 0.05267863, 
    0.141919, 0.241601, 0.1961507, 0.2035764, 0.2568076, 0.2911331, 
    0.1815943, 0.2164596, 0.242208, 0.2600053, 0.2616479, 0.390164, 
    0.4535018, 0.3157557, 0.2922, 0.3429928, 0.2103969,
  0.2453438, 0.1661202, 0.2276508, 0.2613709, 0.2876479, 0.2581531, 
    0.2020477, 0.2536774, 0.2402027, 0.2680594, 0.2561098, 0.353526, 
    0.2752993, 0.2556339, 0.2214939, 0.1848864, 0.1648732, 0.1648662, 
    0.2920208, 0.2422159, 0.2475156, 0.2561141, 0.271877, 0.233102, 
    0.2747432, 0.269543, 0.2308708, 0.1893765, 0.1824242,
  0.134334, 0.1872649, 0.1638501, 0.227325, 0.2075251, 0.150926, 0.1361611, 
    0.1440991, 0.1511523, 0.1749063, 0.1724856, 0.1726411, 0.176623, 
    0.1335319, 0.106299, 0.0518816, 0.1128103, 0.148595, 0.1450441, 
    0.1708118, 0.1277008, 0.09737916, 0.2138461, 0.1684782, 0.09969514, 
    0.1780198, 0.1580793, 0.1100373, 0.1377423,
  0.1112109, 0.0818409, 0.03672468, 0.07653658, 0.08498497, 0.05148805, 
    0.0952739, 0.03927405, 0.03521969, 0.03971694, 0.08746649, 0.05076332, 
    0.1024092, 0.1361394, 0.05581288, 0.03246282, 0.09409317, 0.06275804, 
    0.06881969, 0.06209202, 0.1240041, 0.1248896, 0.07484648, 0.0274834, 
    0.04925005, 0.05972425, 0.03155583, 0.1095615, 0.1165355,
  0.01392566, 0.0001287293, 0.01935929, 0.02565861, 0.03072063, 0.0966931, 
    0.06597563, 0.05561176, 0.07026798, 0.06590848, 0.1345057, 0.1264359, 
    0.05468822, 0.1365795, 0.03497847, -7.574945e-05, 0.06122421, 0.1582478, 
    0.1481237, 0.07808778, 0.06747494, 0.03246915, 0.01066934, -4.79047e-05, 
    0.0248716, 0.01162393, 0.1128677, 0.07117133, 0.02187768,
  4.302886e-08, 0.06422896, 0.001489692, 0.001728127, 0.1159148, 0.005022449, 
    0.03455264, 0.04301434, 0.03693825, 0.004889144, 0.06667117, 0.00262671, 
    0.001302525, 0.0326676, 0.0336463, 0.13652, 0.05178648, 0.06631535, 
    0.06183729, 0.01928755, 0.001148276, -2.012029e-06, 3.900847e-06, 
    0.002385541, 0.06680308, 0.08796585, 0.08140103, 0.01074645, 5.222435e-06,
  0.0007608028, 0.1091029, 0.2219166, 0.08148564, 0.05205185, 0.04166448, 
    0.052857, 0.04790825, 0.09401407, 0.006053952, 0.06489798, 0.05239, 
    0.01251357, 0.01293296, 0.01504089, 0.05148818, 0.05665643, 0.05103363, 
    0.01711978, 9.24386e-05, -2.589282e-05, -0.0007955044, 0.002177689, 
    0.1833322, 0.1996623, 0.07452396, 0.008802294, 0.0009082409, 0.0001754143,
  0.01854313, 0.04754297, 0.04024702, 0.01495999, 0.002471821, 0.005829607, 
    0.003893572, 0.01240096, 0.07874964, 0.1459479, 0.0308589, 0.02152123, 
    0.06266301, 0.0320287, 0.00856986, 0.03919441, 0.01603061, 0.001184594, 
    0.00133299, 0.01965235, 0.02235832, 0.001641563, 0.05604263, 0.05918258, 
    0.11756, 0.0388003, 0.01103293, 0.008538456, 0.007455437,
  4.291654e-06, 1.483254e-06, -0.0001588041, 3.935832e-06, 3.611476e-05, 
    5.254303e-05, 0.0034766, 0.05603127, 0.03015961, 0.02875779, 0.0503455, 
    0.03348035, 0.0204374, 0.03751342, 0.01194837, 0.01917282, 0.04422741, 
    0.04516427, 0.1261402, 0.0893229, 0.01709902, 0.00259558, 4.284207e-05, 
    2.275491e-05, 0.0009711864, 1.563135e-05, -3.470905e-08, 0.004164274, 
    0.005582953,
  0.01038913, 0.002107987, 7.291847e-08, 1.007952e-05, 9.272513e-07, 
    -1.50349e-09, 0.0005125473, 7.529284e-08, -4.227355e-06, 0.01093873, 
    0.02848705, 0.02567155, 0.002400507, 0.01019267, 1.047666e-05, 
    2.602693e-05, 0.02440171, 1.70265e-05, 0.05953383, 0.0359421, 0.03050994, 
    0.002370867, 0.007169027, -0.0002081829, 0.0001399132, 0.002316722, 
    0.00104178, -1.24747e-07, 0.006473916,
  0.02210115, 0.004360073, 0.008766428, 0.002349803, 0.05169709, 0.0154279, 
    0.03039152, 0.01555112, 0.1624094, 0.2045348, 0.1608534, 0.1084231, 
    0.09170949, 0.09688969, 0.04543543, 0.033369, 0.05032099, 0.03179588, 
    0.03648221, 0.04228274, 0.03937515, 0.06247654, 0.08953779, 0.07349072, 
    0.0757817, 0.05189043, 0.04335125, 0.04598562, 0.01586498,
  0.02512675, 0.04958803, 0.101805, 0.112078, 0.1541288, 0.1172153, 
    0.1640214, 0.133202, 0.1097189, 0.1127403, 0.1111782, 0.08051939, 
    0.1684144, 0.1582178, 0.1731237, 0.1525063, 0.2117814, 0.2038135, 
    0.1860454, 0.1634626, 0.1326706, 0.1712562, 0.1619181, 0.2129519, 
    0.1971086, 0.2818461, 0.09804876, 0.09730078, 0.07896965,
  0.1653739, 0.2037759, 0.1985307, 0.182831, 0.1618992, 0.1534682, 0.2221593, 
    0.08830103, 0.05162296, 0.0874353, 0.03030842, 0.09587143, 0.1129689, 
    0.1318062, 0.1780802, 0.2091195, 0.2296697, 0.2142964, 0.2841121, 
    0.2181701, 0.1691477, 0.1811859, 0.1692865, 0.1225583, 0.1342912, 
    0.2341504, 0.1873699, 0.1645339, 0.1727533,
  0.2857755, 0.3234228, 0.2489054, 0.243868, 0.2222811, 0.1928296, 0.2113607, 
    0.1946833, 0.1791055, 0.1714783, 0.1018032, 0.05414629, 0.1303456, 
    0.1708336, 0.2586584, 0.1664193, 0.1257454, 0.2371673, 0.1904889, 
    0.2202812, 0.1159982, 0.1378036, 0.1492534, 0.1471303, 0.1488737, 
    0.1137348, 0.1824951, 0.3071115, 0.267532,
  0.1589585, 0.1721978, 0.2185102, 0.2131511, 0.1900628, 0.1551542, 
    0.1716841, 0.1490316, 0.08984232, 0.1411758, 0.100613, 0.09446091, 
    0.1369758, 0.1551632, 0.1682839, 0.1446182, 0.07273484, 0.1179843, 
    0.06991621, 0.1151465, 0.1450779, 0.08336501, 0.004468965, -0.003986569, 
    0.09018067, 0.0157683, 0.008974343, 0.1672901, 0.1664867,
  0.07187435, 0.07398171, 0.04529598, 0.06062654, 0.0681209, 0.04746723, 
    0.07182143, 0.09375455, 0.06085463, 0.06435271, 0.08637487, 0.1087235, 
    0.1243927, 0.1979306, 0.1994854, 0.2262674, 0.2978244, 0.3013889, 
    0.2010458, 0.1217211, 0.06539584, 0.02110592, -0.0007703258, 
    -0.001571066, 0.0571497, 0.004696163, 0.001829125, 0.0821768, 0.08604014,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.978006e-05, -1.978006e-05, 
    -1.978006e-05, -1.978006e-05, -1.978006e-05, -1.978006e-05, 
    -1.978006e-05, 0, 0, 0, 0, 0, 0, 0, 0,
  0.003174752, -0.0001079531, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.03632e-06, 
    0.1109582, 0.1305692, 0.1541451, 0.2151949, 0.2857336, 0.146537, 
    0.07753736, 0.0362121, 0.009358718, 0.04952151, 0.2751441, 0.3258459, 
    0.4289711, 0.4978973, 0.2387217, 0.04011058,
  0.1233394, 0.1847206, 0.3342774, 0.3367856, 0.02663539, 0.0127869, 
    0.1678161, 0.04974532, 0.02576246, 0.1045813, 0.1326906, 0.1005256, 
    0.172234, 0.2773394, 0.2353706, 0.2444555, 0.2694797, 0.2919672, 
    0.1989834, 0.1975564, 0.2483975, 0.2882877, 0.2824339, 0.3857767, 
    0.4580833, 0.3072991, 0.2984512, 0.3323848, 0.2086897,
  0.2184386, 0.1846534, 0.2291329, 0.2706696, 0.2996799, 0.2455661, 
    0.2212718, 0.2533418, 0.250248, 0.2827241, 0.2590635, 0.3485661, 
    0.2758884, 0.2506564, 0.2001531, 0.1855762, 0.1548436, 0.1573946, 
    0.2929458, 0.285426, 0.2464312, 0.2568657, 0.2853295, 0.234463, 
    0.2704909, 0.2869177, 0.2001566, 0.1961888, 0.1937331,
  0.1430075, 0.2004386, 0.1728249, 0.2003585, 0.1949562, 0.1512608, 
    0.1472641, 0.1217028, 0.1503063, 0.1799455, 0.1912163, 0.1903815, 
    0.1809084, 0.1309131, 0.1139976, 0.05258586, 0.09794775, 0.1628564, 
    0.1452207, 0.1591126, 0.1394798, 0.1051022, 0.1857306, 0.1560854, 
    0.08035456, 0.1563981, 0.1840834, 0.1216239, 0.1240777,
  0.104819, 0.08409165, 0.03369055, 0.06326726, 0.07918368, 0.04125302, 
    0.09530428, 0.04110284, 0.02878767, 0.03927721, 0.09598016, 0.04402427, 
    0.1047456, 0.1304492, 0.04728427, 0.02623342, 0.09287498, 0.07252747, 
    0.06501308, 0.0515413, 0.099545, 0.1079891, 0.07991005, 0.02831087, 
    0.04950959, 0.05128009, 0.02747748, 0.1019036, 0.1104387,
  0.01541789, 2.25543e-05, 0.01763719, 0.0177457, 0.03260352, 0.1016925, 
    0.04642441, 0.05418766, 0.05621541, 0.03970829, 0.1163517, 0.1316987, 
    0.05420655, 0.1446856, 0.02467978, -0.0008773311, 0.06275624, 0.1421601, 
    0.1278076, 0.08011622, 0.06400584, 0.02661245, 0.01063297, -1.955462e-05, 
    0.03533896, 0.01259807, 0.1040657, 0.0611303, 0.01911567,
  9.364791e-05, 0.06582959, 0.001370305, 0.002316339, 0.127186, 0.005138619, 
    0.03614394, 0.05750129, 0.03534669, 0.003438555, 0.06486759, 0.003337307, 
    0.002136439, 0.04722091, 0.03228639, 0.1357843, 0.04953671, 0.06858429, 
    0.07234782, 0.01449676, 0.002383011, 2.22129e-07, 1.031843e-05, 
    0.001705588, 0.05517373, 0.0867996, 0.08814654, 0.008092673, 8.986814e-06,
  0.0009783014, 0.1007139, 0.2305064, 0.1044027, 0.05778808, 0.05035357, 
    0.0602209, 0.06195235, 0.09314561, 0.006216214, 0.06168811, 0.05319056, 
    0.01536149, 0.01792737, 0.02562246, 0.04619635, 0.07465473, 0.05847396, 
    0.01897478, 0.0002642294, -6.053529e-05, -0.0006518161, 0.001987532, 
    0.19374, 0.2050625, 0.08331908, 0.01566939, 0.0009533071, 0.0001493166,
  0.05486132, 0.05028482, 0.06212031, 0.01486837, 0.002052502, 0.00442143, 
    0.00337044, 0.01034122, 0.08486514, 0.1521252, 0.02071545, 0.03847194, 
    0.06223975, 0.03228099, 0.009335616, 0.03934116, 0.0194839, 0.001000248, 
    0.0009700335, 0.01257458, 0.01916155, 0.003823192, 0.08175361, 
    0.06011469, 0.129322, 0.04029198, 0.01036263, 0.01024264, 0.01487442,
  5.330937e-06, 4.933286e-06, 0.01470954, 0.0004367497, 1.457546e-06, 
    5.037545e-05, 0.003107115, 0.0613885, 0.02840264, 0.02914389, 0.05877312, 
    0.03787823, 0.01793937, 0.03176496, 0.01216364, 0.04694978, 0.05964658, 
    0.05663877, 0.1242588, 0.1058798, 0.02051346, 0.005990009, 0.0001487989, 
    4.147461e-05, 0.001789285, 3.894556e-06, 2.268611e-07, 1.904074e-05, 
    0.006371276,
  0.0003187194, 0.0189513, -9.285785e-08, 2.110309e-05, -6.554773e-07, 
    1.065685e-09, 0.0009224805, -1.326938e-06, 4.703705e-05, 0.02591814, 
    0.02333063, 0.02716659, 0.001493055, 0.01228173, -0.0002705722, 
    0.0001276892, 0.01699708, 2.873635e-05, 0.05694715, 0.02654117, 
    0.03461749, 0.00326667, 0.008356951, 0.001027091, 0.0006154088, 
    0.008367249, 0.0003365608, -3.167075e-07, 0.001571773,
  0.01010693, 0.002132725, 0.01076514, 0.004496007, 0.08011734, 0.02038613, 
    0.04168829, 0.03437632, 0.2103346, 0.1871076, 0.1585593, 0.1043034, 
    0.09872341, 0.09206693, 0.043775, 0.02636163, 0.03992866, 0.02123983, 
    0.02433679, 0.03344723, 0.0282281, 0.06057199, 0.09355919, 0.05883084, 
    0.06688141, 0.0521094, 0.05881943, 0.04360712, 0.008549011,
  0.02065019, 0.05017276, 0.09874084, 0.1157847, 0.1353728, 0.1032536, 
    0.1822949, 0.09589001, 0.08693701, 0.08056295, 0.1111319, 0.07393309, 
    0.1508658, 0.1598615, 0.1791403, 0.1251859, 0.1933173, 0.169553, 
    0.1526469, 0.1658972, 0.1709078, 0.1501337, 0.1601353, 0.2146472, 
    0.1880517, 0.2670515, 0.07725026, 0.08691514, 0.0554451,
  0.1455474, 0.2085387, 0.2194413, 0.1676466, 0.1460484, 0.1396877, 
    0.2042619, 0.1347405, 0.1048692, 0.08467738, 0.06990557, 0.1199083, 
    0.1252557, 0.1435071, 0.194676, 0.2123648, 0.2194173, 0.2103813, 
    0.2870398, 0.2376373, 0.1469893, 0.1600164, 0.1819649, 0.1533887, 
    0.1305756, 0.2125641, 0.1805788, 0.1451085, 0.1480704,
  0.2752971, 0.3303174, 0.2450447, 0.2457277, 0.2542695, 0.2056887, 
    0.2481308, 0.1997634, 0.2050724, 0.2102001, 0.1232687, 0.087074, 
    0.2175803, 0.1797017, 0.2610365, 0.193821, 0.1469814, 0.2667248, 
    0.2974443, 0.223847, 0.122858, 0.140422, 0.1425084, 0.2549662, 0.1649241, 
    0.116286, 0.1835795, 0.2720111, 0.2278141,
  0.2296336, 0.1786658, 0.3130409, 0.2208409, 0.1609933, 0.1622615, 
    0.1989625, 0.2077672, 0.1182781, 0.1889829, 0.1486821, 0.114209, 
    0.1735313, 0.1541505, 0.1628743, 0.1433018, 0.1137543, 0.1410623, 
    0.08766986, 0.1401394, 0.1802042, 0.1152027, 0.02152076, 0.008755863, 
    0.1698138, 0.0322859, 0.01959095, 0.3158392, 0.2059936,
  0.08253787, 0.1024711, 0.09981383, 0.1171127, 0.109821, 0.1018457, 
    0.1246142, 0.2167795, 0.1926207, 0.2069631, 0.218957, 0.1595543, 
    0.1475981, 0.2086979, 0.2250981, 0.2644818, 0.3211262, 0.3013433, 
    0.1904368, 0.1070864, 0.09643853, 0.08822347, 0.03643783, -0.0001726851, 
    0.1113164, 0.02528814, 0.0461239, 0.09258667, 0.1358154,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0003183224, -0.0003183224, 
    -0.0003183224, -0.0003183224, -0.0003183224, -0.0003183224, 
    -0.0003183224, 0, 0, 0, 0, 0, 0, 0, 0,
  0.0223729, 0.004021255, -9.234048e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0004235262, 0.195961, 0.2337268, 0.2331291, 0.2447111, 0.2953301, 
    0.2434568, 0.1265682, 0.05332172, 0.01420843, 0.09094834, 0.3075281, 
    0.3670296, 0.4438245, 0.5106391, 0.397843, 0.1100109,
  0.1355631, 0.2030481, 0.3143632, 0.3567931, 0.05727657, 0.03763818, 
    0.2105583, 0.1019966, 0.08038334, 0.1681672, 0.2382542, 0.1342635, 
    0.1781356, 0.3221549, 0.2274861, 0.2390141, 0.3245586, 0.2878636, 
    0.2278797, 0.199212, 0.2340465, 0.2902838, 0.2691027, 0.4290781, 
    0.4808933, 0.3281486, 0.317549, 0.3417115, 0.2173274,
  0.2099235, 0.2014179, 0.2310977, 0.2924302, 0.3077396, 0.2673489, 
    0.2383783, 0.2760408, 0.2630474, 0.2958228, 0.2660162, 0.3336478, 
    0.301095, 0.2523125, 0.2234526, 0.1944506, 0.1469833, 0.1692137, 
    0.3102622, 0.2969151, 0.2571487, 0.2777052, 0.2762694, 0.2443218, 
    0.3004933, 0.3042526, 0.1965509, 0.1993708, 0.2034755,
  0.1592934, 0.1974308, 0.1935723, 0.1884443, 0.1821868, 0.1736959, 0.154114, 
    0.1260942, 0.1439312, 0.1773264, 0.1836925, 0.1851023, 0.1786509, 
    0.1121866, 0.1104167, 0.04347706, 0.09068439, 0.1629711, 0.1708305, 
    0.1577211, 0.1274554, 0.1335882, 0.1911788, 0.1475396, 0.07590216, 
    0.1368762, 0.1911445, 0.1290227, 0.1184973,
  0.09142992, 0.08047426, 0.03545841, 0.05856743, 0.07283885, 0.03863621, 
    0.08267062, 0.0403729, 0.03111156, 0.03727909, 0.0945966, 0.03508098, 
    0.1044672, 0.1440795, 0.04385303, 0.0259144, 0.1055466, 0.06885595, 
    0.07645205, 0.05212538, 0.08836897, 0.1094561, 0.07197756, 0.02713181, 
    0.04804122, 0.05919876, 0.0229472, 0.08984859, 0.1083734,
  0.0165056, 4.056113e-06, 0.01925872, 0.01347332, 0.03119264, 0.1137158, 
    0.03887765, 0.05820767, 0.05204415, 0.02417153, 0.100921, 0.1406194, 
    0.05224738, 0.147808, 0.01768821, 0.001168236, 0.06748842, 0.128807, 
    0.1250781, 0.07670137, 0.0668745, 0.02691705, 0.0115983, 1.073211e-05, 
    0.03574273, 0.01104587, 0.1063924, 0.05333506, 0.0439419,
  1.470552e-05, 0.07553728, 0.002550911, 0.004175331, 0.1534035, 0.006382106, 
    0.03859049, 0.0631012, 0.0472801, 0.004151623, 0.06939614, 0.008588379, 
    0.004753818, 0.07205456, 0.04159452, 0.1604171, 0.06281462, 0.08864287, 
    0.08369874, 0.01821253, 0.002170665, 3.390255e-05, 8.318979e-05, 
    0.0008382619, 0.05418974, 0.09204867, 0.09843983, 0.006873481, 
    2.128441e-06,
  0.008372654, 0.1280396, 0.2654451, 0.1343599, 0.04785331, 0.07270981, 
    0.06831802, 0.07667214, 0.1188325, 0.008929625, 0.08868945, 0.07315432, 
    0.02503651, 0.02839663, 0.05668715, 0.0467011, 0.09087825, 0.06824618, 
    0.02355246, 0.001020186, -6.505466e-05, -0.0006830087, 0.001672753, 
    0.2246524, 0.2421742, 0.1187708, 0.02003107, 0.001081169, 0.0003115072,
  0.09716203, 0.07443456, 0.1122665, 0.02253587, 0.002246629, 0.005664043, 
    0.004772039, 0.01408469, 0.09738977, 0.1761482, 0.02544923, 0.04961377, 
    0.07090974, 0.04469983, 0.01255343, 0.03729477, 0.02443382, 0.002362191, 
    0.002662348, 0.003852751, 0.01659219, 0.02779627, 0.1099045, 0.07641708, 
    0.1450069, 0.05433118, 0.01036029, 0.008959525, 0.07579795,
  0.0001994762, 3.551908e-05, 0.01910132, 0.01817129, 3.936339e-06, 
    0.0002527803, 0.00366347, 0.06530643, 0.02745364, 0.03671524, 0.0688146, 
    0.04109204, 0.02667895, 0.03203657, 0.01191039, 0.07328826, 0.06348903, 
    0.05407812, 0.1130997, 0.1033897, 0.02500381, 0.01441091, 0.001487629, 
    0.0004133343, 0.004876952, 2.796075e-06, 4.535648e-07, 1.795215e-06, 
    0.007077802,
  6.707508e-07, 0.007573467, 8.08924e-08, 0.0001561698, -5.182407e-05, 
    5.488738e-08, 0.005425287, 7.367642e-05, 0.0004325961, 0.04323949, 
    0.007454359, 0.0323744, 0.0003932297, 0.01094724, 8.675509e-05, 
    0.001031812, 0.02288833, 0.0004882424, 0.05051471, 0.01856189, 
    0.02484953, 0.005406358, 0.01086932, 0.004169572, 0.0009163005, 
    0.01615813, 0.003239148, 3.011965e-07, 0.0009775945,
  0.001454536, 0.000358223, 0.01420902, 0.01037702, 0.1025294, 0.02032518, 
    0.05025692, 0.04537028, 0.219836, 0.1799962, 0.1564623, 0.1029767, 
    0.1037489, 0.0874323, 0.05026889, 0.02803015, 0.03910638, 0.0150209, 
    0.01780668, 0.02254989, 0.01635394, 0.05482724, 0.09259532, 0.04234428, 
    0.06225556, 0.05471672, 0.05938872, 0.04009826, 0.009184026,
  0.01668141, 0.05197199, 0.09188907, 0.124883, 0.1200749, 0.09113405, 
    0.2002736, 0.06728303, 0.0754347, 0.06399086, 0.1208818, 0.07572905, 
    0.1361758, 0.1551377, 0.1790992, 0.1381979, 0.1687179, 0.1380238, 
    0.1448491, 0.1708306, 0.1717435, 0.1567864, 0.148592, 0.1980638, 
    0.1833666, 0.2562635, 0.07031604, 0.08079094, 0.0499227,
  0.1042924, 0.2192964, 0.2148252, 0.1471849, 0.1381663, 0.1450236, 
    0.1875029, 0.1323826, 0.1159675, 0.07560983, 0.105685, 0.1188259, 
    0.1198516, 0.1462634, 0.1926643, 0.2044152, 0.2235767, 0.2148719, 
    0.2841966, 0.2421703, 0.1350099, 0.1322235, 0.1767015, 0.1738959, 
    0.1224675, 0.2089757, 0.1765761, 0.1368159, 0.1234404,
  0.2783501, 0.3366188, 0.2307526, 0.2246293, 0.2692713, 0.2068748, 
    0.2492057, 0.1974122, 0.2292894, 0.2761365, 0.130888, 0.1641922, 
    0.2483117, 0.1846556, 0.2683449, 0.1798025, 0.1499699, 0.2885006, 
    0.3187718, 0.2007497, 0.117813, 0.1205334, 0.138991, 0.2772048, 
    0.1667593, 0.1206896, 0.1720028, 0.2760243, 0.2570423,
  0.233388, 0.1703261, 0.2966493, 0.212184, 0.1742186, 0.172075, 0.2268268, 
    0.2815036, 0.1351609, 0.1828192, 0.1481601, 0.1318015, 0.1745465, 
    0.1301731, 0.1585456, 0.1477048, 0.1318103, 0.130134, 0.09528475, 
    0.1318024, 0.1731141, 0.1149358, 0.04976366, 0.03482736, 0.2307482, 
    0.05636434, 0.05316038, 0.3509523, 0.1821144,
  0.08507047, 0.1337658, 0.1189375, 0.126388, 0.1363049, 0.1226807, 
    0.1691506, 0.2572884, 0.2941155, 0.2892463, 0.2771411, 0.1693668, 
    0.1331227, 0.1860307, 0.22767, 0.2575317, 0.3103052, 0.2703893, 
    0.1681232, 0.1069391, 0.0948588, 0.1046752, 0.1061049, 0.03765782, 
    0.1651058, 0.05215966, 0.0978247, 0.1377541, 0.1337465,
  0, 0, 0, 0, 0, 0, 0, -0.000539644, -0.0003567138, -0.0001737837, 
    9.146507e-06, 0.0001920767, 0.0003750068, 0.000557937, -0.001319912, 
    -0.001253392, -0.001186872, -0.001120352, -0.001053832, -0.0009873121, 
    -0.0009207919, 0.0004748928, 0.0002254426, -2.400757e-05, -0.0002734578, 
    -0.000522908, -0.0007723582, -0.001021808, 0,
  0.06323196, 0.03809451, 0.002313688, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.004333755, 0.2665286, 0.2553008, 0.2417393, 0.287313, 0.3127555, 
    0.2970343, 0.2050428, 0.09680932, 0.05595027, 0.184464, 0.3437552, 
    0.3980395, 0.4653608, 0.5455257, 0.4271663, 0.218286,
  0.1486648, 0.2226713, 0.2993512, 0.3249733, 0.1142175, 0.04955529, 
    0.2211774, 0.2055662, 0.1434824, 0.2210556, 0.2848759, 0.1691916, 
    0.1770188, 0.3469745, 0.2526777, 0.2689724, 0.3495904, 0.2945414, 
    0.2523839, 0.2126391, 0.2322811, 0.2687959, 0.2551906, 0.3928166, 
    0.5112602, 0.3332934, 0.3103738, 0.3291882, 0.2321463,
  0.2191784, 0.2079056, 0.2382154, 0.3168787, 0.2586567, 0.2636827, 
    0.2551398, 0.323117, 0.2858456, 0.3258493, 0.2212133, 0.3199757, 
    0.2819467, 0.2422391, 0.2118672, 0.1595972, 0.1669527, 0.1926748, 
    0.3222209, 0.2679384, 0.2119022, 0.2231837, 0.2991073, 0.2503071, 
    0.3010439, 0.296979, 0.2563044, 0.2223161, 0.1978287,
  0.1574063, 0.2116186, 0.1957146, 0.1878101, 0.1779244, 0.1536521, 
    0.1563307, 0.1440427, 0.1420348, 0.2011034, 0.2169074, 0.1751406, 
    0.1694117, 0.1170819, 0.1142482, 0.04840959, 0.09266987, 0.173945, 
    0.1547161, 0.1858542, 0.1331365, 0.1205848, 0.191415, 0.1435691, 
    0.07683499, 0.1223331, 0.1978844, 0.1115597, 0.1299391,
  0.09268308, 0.08008192, 0.0392985, 0.06537959, 0.0651084, 0.03535692, 
    0.08092579, 0.04215613, 0.04118849, 0.0434841, 0.07577351, 0.03913728, 
    0.1115965, 0.1547239, 0.04216112, 0.0218011, 0.1194123, 0.07408977, 
    0.08148632, 0.06125888, 0.08407652, 0.09956513, 0.06935829, 0.02261375, 
    0.04320577, 0.05882252, 0.02278006, 0.08456995, 0.1161676,
  0.01511902, 1.828328e-05, 0.0176173, 0.01115211, 0.04005424, 0.119449, 
    0.04214288, 0.07891385, 0.0400931, 0.02349538, 0.08601066, 0.1266557, 
    0.05316188, 0.1457933, 0.01683321, 0.008582532, 0.07239397, 0.1256119, 
    0.1213137, 0.07591692, 0.06796606, 0.04855486, 0.01416871, 0.0003242962, 
    0.03180226, 0.01182089, 0.1080041, 0.04815547, 0.04572508,
  0.0002024658, 0.08332622, 0.003258783, 0.008242226, 0.1782728, 0.005684626, 
    0.0490502, 0.07289799, 0.04612545, 0.005059131, 0.07170428, 0.008779677, 
    0.005051534, 0.08419292, 0.05013008, 0.1624083, 0.07640809, 0.09682051, 
    0.0988927, 0.03357038, 0.005484475, 3.976578e-05, 0.0001070912, 
    0.000651294, 0.05667202, 0.09364963, 0.1189689, 0.003880517, 3.10108e-06,
  0.006553216, 0.1297338, 0.2978507, 0.1637826, 0.05400215, 0.07329217, 
    0.07076624, 0.08604789, 0.1311213, 0.009971489, 0.09644704, 0.1054511, 
    0.04637097, 0.03280596, 0.0611912, 0.06257652, 0.1056539, 0.06913764, 
    0.02323517, 0.001869412, -3.258414e-05, -0.001054763, 0.001975852, 
    0.267326, 0.2819277, 0.171867, 0.0411082, 0.001258163, 0.000200844,
  0.1149627, 0.1023967, 0.1467914, 0.04203818, 0.001995605, 0.006831606, 
    0.009672975, 0.01208169, 0.1147883, 0.2129535, 0.03276109, 0.05286251, 
    0.07848372, 0.05904846, 0.01460333, 0.03994181, 0.02859931, 0.002523259, 
    0.004487617, 0.001404991, 0.01173623, 0.03176725, 0.117802, 0.1219973, 
    0.1621424, 0.06908298, 0.008339748, 0.00752859, 0.02554844,
  0.003002298, 1.389272e-06, 0.01527633, 0.08151007, 9.612912e-06, 
    0.0001680086, 0.004483776, 0.08310913, 0.0337873, 0.03931102, 0.08079883, 
    0.05068455, 0.04231668, 0.03700895, 0.01823965, 0.06965169, 0.06648535, 
    0.04048572, 0.1063424, 0.1018763, 0.0329006, 0.01990627, 0.002500849, 
    0.001163824, 0.002693825, 2.139999e-05, 3.562982e-07, -5.208576e-06, 
    0.02754146,
  3.602167e-06, -4.897095e-05, 2.592804e-07, -2.828038e-06, -1.808511e-05, 
    5.68783e-08, 0.01478936, 0.0004989372, 0.001175066, 0.0541116, 
    0.004655775, 0.04859203, 0.0001588184, 0.01281464, -8.807688e-05, 
    0.001680649, 0.03053429, 0.004630825, 0.04451624, 0.01974432, 0.01983665, 
    0.006315109, 0.01093493, 0.009615042, 0.001812804, 0.03549657, 
    0.005443034, 1.228219e-07, 1.638827e-06,
  3.52635e-05, 5.551376e-05, 0.01965639, 0.01340214, 0.1131423, 0.01703112, 
    0.03072698, 0.05085017, 0.2205543, 0.1832001, 0.1653203, 0.1004629, 
    0.1091727, 0.09228551, 0.05023436, 0.03065891, 0.04631979, 0.01377037, 
    0.022594, 0.01521865, 0.01207638, 0.06001399, 0.08844405, 0.04002887, 
    0.06137966, 0.06422935, 0.04407687, 0.03106838, 0.005880383,
  0.01077273, 0.05981962, 0.08108356, 0.138847, 0.1131172, 0.07898393, 
    0.2070401, 0.0429181, 0.0747555, 0.07835775, 0.1298279, 0.0818138, 
    0.1266152, 0.1468323, 0.1736174, 0.1367642, 0.1594265, 0.1360242, 
    0.1512619, 0.1667129, 0.1618866, 0.1666828, 0.1387454, 0.1852427, 
    0.1773722, 0.2575822, 0.07961067, 0.06957109, 0.04938933,
  0.09114947, 0.2209689, 0.1971501, 0.1485005, 0.1487504, 0.1523498, 
    0.1750522, 0.1163264, 0.1060163, 0.1119685, 0.1016009, 0.1156934, 
    0.1136186, 0.1473945, 0.1944094, 0.2116079, 0.2289969, 0.2194196, 
    0.2712342, 0.2341695, 0.132736, 0.1168862, 0.1588888, 0.174911, 
    0.1343476, 0.2094774, 0.1740478, 0.1272621, 0.1058005,
  0.2621518, 0.3401049, 0.2065668, 0.2120771, 0.2842006, 0.2144496, 
    0.2305473, 0.1987943, 0.2326103, 0.3228, 0.1595398, 0.1839181, 0.2411748, 
    0.1965929, 0.2584118, 0.1583162, 0.1451756, 0.3089501, 0.3356674, 
    0.1771462, 0.1076928, 0.1225077, 0.1387427, 0.2997063, 0.1590474, 
    0.09988545, 0.1413899, 0.27571, 0.2278345,
  0.2195918, 0.1678805, 0.2916196, 0.2163525, 0.2014423, 0.1757151, 0.241161, 
    0.3197435, 0.1805026, 0.1887438, 0.1453629, 0.1539271, 0.1699272, 
    0.1224627, 0.1427969, 0.1518686, 0.1378483, 0.1362869, 0.1024474, 
    0.1334704, 0.1912415, 0.1201275, 0.08009775, 0.1079242, 0.2831309, 
    0.0935426, 0.08202314, 0.3516219, 0.1809585,
  0.0802814, 0.133475, 0.1277924, 0.1334852, 0.1374887, 0.1288909, 0.1702246, 
    0.2884523, 0.2923454, 0.2919994, 0.27659, 0.1691469, 0.1234747, 0.15279, 
    0.2381376, 0.2394722, 0.2873537, 0.2281276, 0.1508352, 0.1028281, 
    0.0903988, 0.1139173, 0.1249875, 0.08722693, 0.1947335, 0.1214478, 
    0.1434617, 0.1300842, 0.1110777,
  0.002499975, 0.001813969, 0.001127962, 0.0004419556, -0.000244051, 
    -0.0009300576, -0.001616064, -0.001412549, -0.0007473484, -8.214777e-05, 
    0.0005830528, 0.001248253, 0.001913454, 0.002578655, -0.002462793, 
    -0.0004517538, 0.001559286, 0.003570325, 0.005581365, 0.007592404, 
    0.009603444, 0.01535166, 0.01336143, 0.0113712, 0.009380965, 0.007390731, 
    0.005400497, 0.003410264, 0.003048781,
  0.1488183, 0.03445232, 0.02368113, -0.0002060283, 0, -0.0008181843, 
    -0.0005882164, -0.0001171175, 0, 0, 0, 0.001646066, 0.06478896, 
    0.2783527, 0.2221462, 0.245205, 0.2551973, 0.309858, 0.305832, 0.2255095, 
    0.1920248, 0.2279655, 0.2476252, 0.3274505, 0.4000269, 0.492679, 
    0.6026374, 0.4618652, 0.3587185,
  0.1905726, 0.2271934, 0.2973143, 0.2895028, 0.1314627, 0.04273991, 
    0.2639786, 0.261964, 0.1715019, 0.259299, 0.3157426, 0.1944834, 
    0.1912661, 0.3705319, 0.261265, 0.2962096, 0.3854905, 0.2818673, 
    0.1968462, 0.185555, 0.2014172, 0.2638227, 0.2465081, 0.4005333, 
    0.5108014, 0.3361913, 0.3620947, 0.352595, 0.2461157,
  0.2144539, 0.2112754, 0.2403618, 0.3303895, 0.2926598, 0.3013358, 
    0.2856552, 0.360765, 0.3189623, 0.3321224, 0.2353977, 0.312543, 
    0.3331208, 0.219685, 0.228333, 0.1689124, 0.1824768, 0.205747, 0.2972746, 
    0.2393442, 0.2015929, 0.2469179, 0.3080308, 0.2349565, 0.2813515, 
    0.2985396, 0.2651169, 0.2305105, 0.2115603,
  0.180528, 0.216031, 0.1902915, 0.1777387, 0.1969745, 0.1645637, 0.157449, 
    0.1534303, 0.1524296, 0.1741549, 0.2061726, 0.1813649, 0.1835993, 
    0.1374964, 0.1065364, 0.07619992, 0.09904119, 0.1835491, 0.1881088, 
    0.1985777, 0.1395901, 0.1343353, 0.1866065, 0.1362138, 0.07614236, 
    0.1216823, 0.1923927, 0.1088908, 0.1347719,
  0.1002558, 0.08556587, 0.04062376, 0.0669013, 0.07028749, 0.04256463, 
    0.09183202, 0.05169352, 0.05402379, 0.04121968, 0.06290273, 0.05763372, 
    0.1219895, 0.1631684, 0.05378275, 0.02317717, 0.1395131, 0.09610886, 
    0.08342204, 0.06177599, 0.08809423, 0.09277372, 0.07715465, 0.026112, 
    0.04548196, 0.06117875, 0.03557883, 0.08705234, 0.1196717,
  0.01197992, 0.0006574758, 0.02505287, 0.008982311, 0.04713753, 0.1109758, 
    0.05516435, 0.06702964, 0.02301785, 0.02276088, 0.07320176, 0.1104893, 
    0.05161672, 0.1519983, 0.02844358, 0.01235651, 0.09380145, 0.1236352, 
    0.1223963, 0.08209449, 0.0750581, 0.06356176, 0.0181662, 0.001334298, 
    0.04065532, 0.01150802, 0.1055869, 0.05615887, 0.04176027,
  0.0002223004, 0.1007709, 0.00691205, 0.018503, 0.1703898, 0.005927569, 
    0.05467525, 0.04783644, 0.02160081, 0.004311403, 0.063461, 0.009119765, 
    0.01155079, 0.07312189, 0.05429409, 0.1542955, 0.07056928, 0.07078534, 
    0.0959998, 0.03902448, 0.016045, 0.0004276677, 3.67956e-05, 0.0003066408, 
    0.05315547, 0.1271506, 0.1179247, 0.02040298, 1.008954e-06,
  0.004049649, 0.1163649, 0.3456879, 0.1667459, 0.04392513, 0.06497609, 
    0.05503825, 0.06426585, 0.1039826, 0.009184158, 0.08916209, 0.07035975, 
    0.04862786, 0.02823616, 0.06655166, 0.06487998, 0.08910215, 0.06539488, 
    0.02169742, 0.002294602, 9.211284e-05, -0.001170539, 0.001207125, 
    0.2789519, 0.2775256, 0.2000962, 0.02907502, 0.001239399, 0.0002781875,
  0.03783212, 0.1077985, 0.1441043, 0.04372862, 0.001811326, 0.006147815, 
    0.006189893, 0.007060484, 0.1348306, 0.2305304, 0.04073662, 0.03759908, 
    0.0650891, 0.04641694, 0.01354263, 0.04246062, 0.02808727, 0.003107355, 
    0.003030604, 0.001050523, 0.008154552, 0.00946282, 0.1028054, 0.1532983, 
    0.157175, 0.07793514, 0.009464173, 0.00753731, 0.005698413,
  0.0007240196, 0.0001928347, 0.0005040613, 0.1498922, 1.926946e-06, 
    0.0004982375, 0.005337563, 0.0843087, 0.02704949, 0.03826612, 0.07965829, 
    0.04800304, 0.04218429, 0.03538289, 0.01268234, 0.06755296, 0.0610168, 
    0.02084214, 0.08393855, 0.09608898, 0.02965005, 0.01856113, 0.002218283, 
    0.00170619, 0.001600865, 7.189046e-06, 4.470676e-07, -7.96623e-06, 
    0.04338774,
  1.316569e-06, -8.684507e-07, 1.820301e-07, 1.549893e-07, -8.832534e-07, 
    4.180666e-08, 0.02591226, 0.0004303578, 0.01601046, 0.04886432, 
    0.002429025, 0.05756808, 0.0002513322, 0.01299568, 4.415048e-05, 
    0.002428802, 0.03284384, 0.002119476, 0.03348767, 0.03442241, 
    0.004358933, 0.01392391, 0.02192266, 0.0267741, 0.003160083, 0.0397335, 
    3.083736e-05, 7.806524e-08, 7.783368e-07,
  9.741974e-06, 0.0001139014, 0.01555827, 0.01398409, 0.111246, 0.01229973, 
    0.005029697, 0.06415526, 0.2121159, 0.200083, 0.1617496, 0.1047707, 
    0.108481, 0.08923171, 0.05377612, 0.03672613, 0.05214033, 0.01603756, 
    0.01888691, 0.008976148, 0.01354781, 0.05407327, 0.07105587, 0.04193844, 
    0.06321976, 0.0703885, 0.04117775, 0.01920057, 0.001683228,
  0.007639192, 0.05202879, 0.07504409, 0.1563732, 0.1037572, 0.0674184, 
    0.2047157, 0.02916498, 0.06827274, 0.08477682, 0.1297769, 0.09449349, 
    0.1225813, 0.1583005, 0.1735806, 0.1419658, 0.147695, 0.1434141, 
    0.1471427, 0.162329, 0.1577459, 0.1647591, 0.1329022, 0.180897, 0.170485, 
    0.2404104, 0.07402108, 0.06411855, 0.04293473,
  0.08717148, 0.2201457, 0.2097092, 0.1508219, 0.140671, 0.1528121, 
    0.1620476, 0.1067427, 0.09246851, 0.1213647, 0.1016425, 0.1132528, 
    0.1134997, 0.1467519, 0.1869332, 0.2327649, 0.2456401, 0.2418813, 
    0.2498397, 0.2151512, 0.1402283, 0.1137801, 0.1701607, 0.1769775, 
    0.1269232, 0.2112659, 0.1687924, 0.1220338, 0.1012597,
  0.2653148, 0.329183, 0.2121962, 0.2219509, 0.2679305, 0.2008639, 0.2398061, 
    0.1798392, 0.2189658, 0.3244612, 0.1909485, 0.1872253, 0.2419212, 
    0.2222485, 0.2719543, 0.1845489, 0.1581551, 0.3223328, 0.3325889, 
    0.1902934, 0.1161333, 0.1342733, 0.1611326, 0.3671817, 0.1684908, 
    0.1117404, 0.1493636, 0.2956513, 0.2344291,
  0.2508745, 0.1634544, 0.2887157, 0.2340089, 0.2400271, 0.1732149, 
    0.2597302, 0.3374809, 0.1937723, 0.1827961, 0.1815313, 0.1997786, 
    0.1861678, 0.1400438, 0.1228131, 0.1496406, 0.1347938, 0.1359479, 
    0.0990229, 0.1342023, 0.2206778, 0.1317754, 0.1122453, 0.1149737, 
    0.2897493, 0.1700575, 0.1178082, 0.355678, 0.2093373,
  0.0743095, 0.1161754, 0.123092, 0.1387593, 0.1260159, 0.1400744, 0.1878397, 
    0.3093488, 0.2931236, 0.2719445, 0.2499265, 0.1795422, 0.1198104, 
    0.1301954, 0.2309062, 0.2294357, 0.2691389, 0.1872647, 0.1363987, 
    0.0988621, 0.09374914, 0.1337821, 0.129768, 0.1062201, 0.2045488, 
    0.1321918, 0.1488128, 0.1130164, 0.0876282,
  0.03642909, 0.03419077, 0.03195245, 0.02971412, 0.0274758, 0.02523748, 
    0.02299915, 0.04027967, 0.04441135, 0.04854302, 0.05267469, 0.05680636, 
    0.06093803, 0.06506971, 0.06182339, 0.06245338, 0.06308337, 0.06371335, 
    0.06434333, 0.06497332, 0.06560331, 0.0627626, 0.06023926, 0.05771592, 
    0.05519259, 0.05266925, 0.05014592, 0.04762258, 0.03821975,
  0.3008322, 0.05210298, 0.02892633, 0.001891331, -0.000219788, 0.003802068, 
    0.006376036, 0.00335084, 0.006660798, -4.75819e-05, -0.0007815904, 
    0.02032733, 0.1490217, 0.3121953, 0.236053, 0.2843893, 0.3081797, 
    0.3357571, 0.2915398, 0.2180521, 0.2189282, 0.30538, 0.2906042, 
    0.3487171, 0.5008333, 0.5274289, 0.6002336, 0.5376021, 0.3829695,
  0.2249184, 0.2734199, 0.2965854, 0.3024439, 0.131214, 0.04121823, 
    0.3473857, 0.2799918, 0.1719442, 0.3099567, 0.3649928, 0.2167724, 
    0.2012118, 0.4066606, 0.2803608, 0.2746646, 0.373384, 0.2831233, 
    0.2407536, 0.2065617, 0.231385, 0.2633964, 0.2749569, 0.3893376, 
    0.4805931, 0.3597403, 0.3872732, 0.3926852, 0.2458005,
  0.2042781, 0.2317182, 0.2595004, 0.3482832, 0.259238, 0.3012213, 0.2641378, 
    0.3343917, 0.2718069, 0.3508219, 0.2270616, 0.2876575, 0.3312742, 
    0.2390051, 0.2366844, 0.1688468, 0.181386, 0.238242, 0.3001942, 
    0.2706432, 0.227384, 0.2296015, 0.3122777, 0.2653193, 0.2875412, 
    0.3392027, 0.2522797, 0.2277781, 0.2195739,
  0.1893319, 0.2108539, 0.2090596, 0.2111878, 0.2095805, 0.1899788, 
    0.1740419, 0.1631571, 0.1604344, 0.1751917, 0.2406257, 0.176408, 
    0.1745585, 0.1417196, 0.113461, 0.09227411, 0.1188517, 0.1905303, 
    0.1844641, 0.2228357, 0.1544404, 0.1379669, 0.2181904, 0.1357639, 
    0.08225352, 0.1441351, 0.1802384, 0.1233037, 0.1511038,
  0.1088662, 0.09186976, 0.04485271, 0.06918623, 0.08221938, 0.05720551, 
    0.1083379, 0.06772301, 0.0689333, 0.04519027, 0.06880001, 0.03780187, 
    0.1371348, 0.1723984, 0.06673394, 0.03027853, 0.1507348, 0.1124533, 
    0.09212629, 0.07975706, 0.08833158, 0.1005982, 0.08312561, 0.03085576, 
    0.05935844, 0.0663274, 0.04252651, 0.08539589, 0.1346897,
  0.01234056, 9.59004e-05, 0.04160434, 0.004264665, 0.05185921, 0.1033415, 
    0.08754092, 0.05504341, 0.004494789, 0.01779056, 0.07616346, 0.08344208, 
    0.05719037, 0.1747927, 0.03831556, 0.02563833, 0.1157772, 0.1093458, 
    0.1289278, 0.09470592, 0.07025447, 0.07612757, 0.02453887, 0.001655511, 
    0.04698174, 0.0139595, 0.0973409, 0.06034353, 0.038571,
  0.0004858335, 0.1113251, 0.008238916, 0.02759745, 0.159301, 0.008267228, 
    0.05938843, 0.03652638, 0.01452641, 0.001558067, 0.06239655, 0.0157839, 
    0.02122278, 0.06733061, 0.05419433, 0.1410623, 0.06409883, 0.05432813, 
    0.1027521, 0.05056815, 0.03928516, 0.001495835, 8.278847e-06, 
    4.410917e-05, 0.04802726, 0.1367583, 0.09434924, 0.02861518, 0.0001647863,
  0.000996907, 0.08991126, 0.3726707, 0.123542, 0.03021832, 0.05423895, 
    0.04212366, 0.04802231, 0.0872195, 0.008778089, 0.09186283, 0.05044501, 
    0.04773904, 0.02214669, 0.0649285, 0.0579634, 0.08445704, 0.06854326, 
    0.02442555, 0.004446459, -2.099308e-05, -0.001247486, 0.0007292153, 
    0.2325597, 0.2207751, 0.1489436, 0.01558392, 0.001269679, 0.0005420916,
  0.007713831, 0.0657898, 0.08086955, 0.03866927, 0.001564749, 0.006597598, 
    0.005004273, 0.006441731, 0.1184038, 0.1884434, 0.04078766, 0.03037922, 
    0.0496651, 0.04046548, 0.01365461, 0.04000297, 0.0285287, 0.005069339, 
    0.002422153, 0.001903931, 0.01022645, 0.008051319, 0.09453147, 0.1487579, 
    0.1462687, 0.08786888, 0.01348504, 0.01165535, 0.003411542,
  -0.0001752943, 5.475983e-06, 1.448114e-05, 0.2308651, -8.547382e-06, 
    0.001190725, 0.006829679, 0.08279137, 0.02338836, 0.03941308, 0.09076244, 
    0.04705937, 0.04026431, 0.03244787, 0.0109315, 0.0674121, 0.05260302, 
    0.007680308, 0.06708408, 0.0756387, 0.02897178, 0.01220334, 0.00249225, 
    0.00246809, 0.0008141018, 1.338075e-06, 3.016521e-07, 7.546381e-07, 
    0.01462972,
  7.138083e-07, 2.626815e-07, 2.826235e-08, 2.59667e-07, -2.884834e-06, 
    2.63589e-08, 0.02096158, 2.71973e-05, 0.03758111, 0.04490583, 
    0.004084934, 0.03935731, 0.003713394, 0.01335268, 0.0009499589, 
    0.004930735, 0.03027381, 0.0001486777, 0.03939759, 0.01874178, 
    0.001459166, 0.01661649, 0.02383484, 0.035165, 0.002970145, 0.04451109, 
    -0.0001032853, 5.346643e-08, 1.50755e-07,
  1.97334e-06, 3.449387e-05, 0.02338546, 0.01851614, 0.1028081, 0.006711984, 
    -0.001059736, 0.07174911, 0.1952847, 0.2153376, 0.1646965, 0.1117768, 
    0.1250259, 0.1023189, 0.06509502, 0.05282161, 0.06770222, 0.02513796, 
    0.02278093, 0.009782053, 0.01688998, 0.05106457, 0.06260497, 0.04911625, 
    0.0713526, 0.07791173, 0.038134, 0.008425387, 0.0002051871,
  0.005131231, 0.05367554, 0.08309975, 0.1647809, 0.09390001, 0.05600551, 
    0.2071364, 0.02549141, 0.04485862, 0.07786807, 0.1267677, 0.09011076, 
    0.1184054, 0.1721074, 0.1688757, 0.1435123, 0.1373642, 0.1462041, 
    0.1495649, 0.1785835, 0.1438424, 0.1569369, 0.1457025, 0.1877739, 
    0.173387, 0.2457574, 0.06673165, 0.05983782, 0.03821742,
  0.08811311, 0.2551629, 0.2149582, 0.1784252, 0.1707478, 0.1629041, 
    0.1476578, 0.1031942, 0.08761519, 0.1227605, 0.09433486, 0.113905, 
    0.1150889, 0.1525846, 0.2174127, 0.2410314, 0.2394613, 0.2337778, 
    0.2356566, 0.2193123, 0.1568525, 0.1134864, 0.1968002, 0.2203666, 
    0.1482431, 0.200943, 0.1731715, 0.1175598, 0.1149334,
  0.2838813, 0.3183765, 0.245871, 0.2487324, 0.3229329, 0.2113496, 0.2513642, 
    0.1699385, 0.2318905, 0.336266, 0.2156317, 0.185777, 0.2380266, 
    0.2309869, 0.3002274, 0.1582337, 0.1605702, 0.3349986, 0.3342567, 
    0.2492763, 0.09100831, 0.1635173, 0.2079917, 0.3896036, 0.191756, 
    0.1231857, 0.1410119, 0.3112452, 0.2420776,
  0.2508239, 0.1862139, 0.2767281, 0.2549512, 0.2399443, 0.174986, 0.2423515, 
    0.3401867, 0.205565, 0.2134908, 0.2102804, 0.2026412, 0.2119714, 
    0.1455871, 0.1062875, 0.1749904, 0.1564008, 0.1514445, 0.08459424, 
    0.1269379, 0.2435773, 0.1247729, 0.1490903, 0.1102326, 0.3008498, 
    0.2344916, 0.1601072, 0.3809493, 0.2049415,
  0.06236723, 0.119234, 0.1164165, 0.1395572, 0.1164233, 0.144623, 0.1811693, 
    0.3267398, 0.3050555, 0.2607428, 0.2307454, 0.181863, 0.138382, 
    0.1200261, 0.20276, 0.2418687, 0.2539001, 0.1672674, 0.1190192, 
    0.08060414, 0.081585, 0.1383778, 0.1301751, 0.1116604, 0.1993468, 
    0.1713579, 0.1703813, 0.09035853, 0.08074943,
  0.07355022, 0.06964004, 0.06572986, 0.06181968, 0.0579095, 0.05399933, 
    0.05008915, 0.06886929, 0.07231622, 0.07576317, 0.07921011, 0.08265705, 
    0.08610399, 0.08955093, 0.07810053, 0.08435509, 0.09060964, 0.0968642, 
    0.1031188, 0.1093733, 0.1156279, 0.1263573, 0.120566, 0.1147747, 
    0.1089833, 0.103192, 0.0974007, 0.09160937, 0.07667837,
  0.3423942, 0.1291718, 0.03176899, 0.01247251, -0.0002380924, 0.01198573, 
    0.0162224, 0.01774679, 0.01439813, -7.068585e-05, 0.008461281, 
    0.09298785, 0.2092523, 0.3324412, 0.3268489, 0.3056848, 0.3235977, 
    0.3567365, 0.311722, 0.2277775, 0.2418059, 0.3405001, 0.2880791, 
    0.3127567, 0.4120748, 0.5230333, 0.5931301, 0.6041402, 0.3929296,
  0.2078594, 0.2521833, 0.3338584, 0.2897385, 0.1223985, 0.05372635, 
    0.3236777, 0.2718672, 0.1878478, 0.3329723, 0.3783868, 0.2174935, 
    0.1952864, 0.4377426, 0.3248493, 0.3281495, 0.370717, 0.2747398, 
    0.2200684, 0.2244846, 0.2575346, 0.274147, 0.3437589, 0.4537162, 
    0.525814, 0.3995032, 0.344084, 0.4110695, 0.2571935,
  0.2101319, 0.2530899, 0.2833941, 0.342204, 0.2999476, 0.3639749, 0.3321227, 
    0.370999, 0.3681442, 0.3645887, 0.2660261, 0.3017726, 0.3794185, 
    0.2568158, 0.2414579, 0.2136308, 0.2012874, 0.2551182, 0.318217, 
    0.2990199, 0.2285435, 0.2443839, 0.3063996, 0.2860176, 0.275335, 
    0.3121473, 0.2474853, 0.2289727, 0.2914921,
  0.1874429, 0.2646689, 0.2312218, 0.2267286, 0.2113182, 0.1724197, 
    0.1869468, 0.190779, 0.1700603, 0.17643, 0.2453002, 0.1806342, 0.1850564, 
    0.1651829, 0.1188661, 0.1043884, 0.1424904, 0.2036433, 0.2121629, 
    0.2460494, 0.1684629, 0.1441175, 0.221457, 0.1359215, 0.08190747, 
    0.1589925, 0.2049089, 0.1396839, 0.1513264,
  0.109594, 0.102481, 0.04593313, 0.07199667, 0.09633683, 0.06099695, 
    0.1349234, 0.08118404, 0.0617232, 0.07754112, 0.07819316, 0.04496598, 
    0.1508169, 0.1901382, 0.07841834, 0.04704066, 0.1848459, 0.1346085, 
    0.09172028, 0.09015983, 0.09164073, 0.1118178, 0.0870982, 0.03684314, 
    0.06246573, 0.06782027, 0.0251058, 0.08375058, 0.1473408,
  0.01759881, 0.000483405, 0.02808782, 0.004744797, 0.05384217, 0.08152486, 
    0.09060966, 0.04388753, 0.00543743, 0.01606019, 0.04562408, 0.05484587, 
    0.08746593, 0.1485454, 0.0387659, 0.04012619, 0.1083578, 0.0833106, 
    0.1239967, 0.103292, 0.06969367, 0.1002708, 0.04297844, 0.0006092669, 
    0.04248882, 0.02317394, 0.07474995, 0.04724254, 0.04207538,
  0.002674964, 0.0868633, 0.01444595, 0.03309463, 0.1536412, 0.01084249, 
    0.07188095, 0.03965094, 0.01445062, 0.001352732, 0.07920641, 0.02724846, 
    0.03412287, 0.06996234, 0.05778546, 0.1439177, 0.06522492, 0.05200387, 
    0.107389, 0.05765127, 0.05848117, 0.002478044, 3.5773e-06, 1.210305e-05, 
    0.04993738, 0.1015705, 0.08299822, 0.03154174, 0.004392738,
  0.0004824374, 0.08245116, 0.3001597, 0.1004567, 0.02522947, 0.04853133, 
    0.03853971, 0.04124687, 0.07369617, 0.009603029, 0.09176864, 0.04501674, 
    0.04763722, 0.02162606, 0.05838989, 0.05119655, 0.08207891, 0.07326907, 
    0.03238903, 0.01003011, -4.489515e-05, -0.001503861, 7.500218e-05, 
    0.2212679, 0.2138301, 0.1269202, 0.008379439, 0.001043767, 0.0007261022,
  0.002207764, 0.02406608, 0.02668593, 0.03273353, 0.001681401, 0.007224648, 
    0.005884977, 0.007693825, 0.09765205, 0.1753794, 0.04206607, 0.02623428, 
    0.04096742, 0.02948211, 0.01789489, 0.0430487, 0.03392448, 0.008127257, 
    0.002919404, 0.009577862, 0.01420401, 0.01472826, 0.09223668, 0.1387852, 
    0.1548654, 0.08819779, 0.02001816, 0.01162987, 0.003842822,
  1.317e-05, 1.811937e-06, 4.568465e-06, 0.2144525, -3.705518e-05, 
    0.002240236, 0.005548866, 0.08253411, 0.02110789, 0.04211262, 0.1069882, 
    0.05696942, 0.04176366, 0.03191724, 0.0135514, 0.05282326, 0.03686417, 
    0.006636954, 0.06375919, 0.0673822, 0.03636548, 0.011268, 0.007988122, 
    0.009353533, 0.003526931, 2.128016e-06, 1.626027e-07, 5.892817e-07, 
    0.003638681,
  2.528359e-07, 3.02774e-07, -2.523266e-05, 9.152147e-07, 1.050129e-09, 
    1.334053e-08, 0.004083785, -6.929772e-05, 0.05210654, 0.03480518, 
    0.002592049, 0.03573044, 0.01173387, 0.01445684, 0.006163503, 0.01018327, 
    0.03978132, 0.0001120422, 0.04399926, 0.0150758, 0.0001173829, 
    0.04506892, 0.02419492, 0.04766014, 0.004249396, 0.03967016, 
    -6.600495e-05, 4.213261e-08, 1.195824e-07,
  1.085981e-06, -2.425116e-05, 0.02952664, 0.03826321, 0.0929801, 0.00249705, 
    -0.002540639, 0.06492653, 0.1703056, 0.205498, 0.1666997, 0.1268378, 
    0.1228143, 0.1029531, 0.07223739, 0.07033017, 0.07399683, 0.05216927, 
    0.02306023, 0.01488325, 0.01644455, 0.05104976, 0.06796504, 0.05113736, 
    0.07715973, 0.0787012, 0.03297237, 0.006361934, 5.774825e-05,
  0.004385617, 0.05107866, 0.1025362, 0.1725485, 0.07889269, 0.04034154, 
    0.2207696, 0.02305694, 0.01733787, 0.06087161, 0.1193434, 0.07698963, 
    0.1256081, 0.1901268, 0.165373, 0.1402461, 0.1288223, 0.1509441, 
    0.1526784, 0.1649139, 0.1324837, 0.1563171, 0.1834089, 0.2034272, 
    0.1764666, 0.2680466, 0.0727346, 0.05890858, 0.03606296,
  0.1005353, 0.2590158, 0.2251578, 0.2173513, 0.2379109, 0.1968617, 
    0.1485353, 0.1104977, 0.08762926, 0.1038738, 0.07548476, 0.1135416, 
    0.1269813, 0.1704021, 0.2524699, 0.2793228, 0.2472707, 0.2552597, 
    0.2207513, 0.2074009, 0.1664956, 0.1124123, 0.2164301, 0.2380266, 
    0.136575, 0.2046407, 0.1804156, 0.1132454, 0.1399437,
  0.2915456, 0.2986934, 0.2170867, 0.2613184, 0.3993919, 0.2257819, 
    0.2444739, 0.1838584, 0.2598253, 0.3525877, 0.2463699, 0.1784954, 
    0.2786216, 0.2472005, 0.3021714, 0.2053857, 0.1509995, 0.3449193, 
    0.3568527, 0.2304422, 0.09699801, 0.1588153, 0.2467491, 0.3969945, 
    0.1761135, 0.124633, 0.1539025, 0.3311011, 0.2447597,
  0.2409285, 0.1942904, 0.3368599, 0.3577519, 0.3129297, 0.2224808, 
    0.2852018, 0.3499767, 0.2194089, 0.2404003, 0.2339017, 0.1932035, 
    0.1996382, 0.1226373, 0.08990043, 0.1969867, 0.1145042, 0.1369302, 
    0.07443878, 0.1202875, 0.1847384, 0.1083949, 0.1565255, 0.1083182, 
    0.2945553, 0.3549512, 0.2155006, 0.3866732, 0.2286317,
  0.06790544, 0.1410542, 0.1260017, 0.1559623, 0.1348682, 0.1515696, 
    0.1956508, 0.3344482, 0.3323868, 0.2537666, 0.1902219, 0.1688015, 
    0.1566546, 0.1031032, 0.1763227, 0.214802, 0.2395395, 0.1466742, 
    0.102553, 0.06503814, 0.08041032, 0.1458911, 0.1185496, 0.09803472, 
    0.1810096, 0.1855157, 0.1752972, 0.06812251, 0.07076327,
  0.1716236, 0.1668534, 0.1620831, 0.1573128, 0.1525425, 0.1477723, 0.143002, 
    0.1805175, 0.1864962, 0.1924749, 0.1984536, 0.2044323, 0.210411, 
    0.2163897, 0.2013099, 0.2087491, 0.2161883, 0.2236274, 0.2310666, 
    0.2385058, 0.2459449, 0.2157071, 0.2070595, 0.1984119, 0.1897643, 
    0.1811167, 0.1724692, 0.1638216, 0.1754399,
  0.3654023, 0.2743756, 0.03027598, 0.02915926, 0.01169514, 0.01804756, 
    0.02132039, 0.02064863, 0.01474268, 8.608571e-05, 0.02311922, 0.1017639, 
    0.2824987, 0.3543196, 0.3283395, 0.2282524, 0.2611841, 0.344253, 
    0.3346078, 0.2148331, 0.2344726, 0.3464718, 0.2767603, 0.2732132, 
    0.3269026, 0.3867058, 0.4976779, 0.5791278, 0.4073985,
  0.2160498, 0.2047776, 0.33067, 0.2740968, 0.1070133, 0.06299648, 0.2859092, 
    0.2519247, 0.2176337, 0.3350116, 0.3770907, 0.213871, 0.1854514, 
    0.4293626, 0.3673777, 0.3336765, 0.3312412, 0.2938466, 0.2038547, 
    0.2490003, 0.2530189, 0.2423093, 0.2601551, 0.3692887, 0.4760927, 
    0.3562187, 0.3153664, 0.4482391, 0.2545782,
  0.2225719, 0.2791109, 0.3065229, 0.3334863, 0.2808646, 0.3317071, 
    0.3659959, 0.3667449, 0.3708818, 0.331746, 0.2886713, 0.3606909, 
    0.3656091, 0.2404506, 0.2666641, 0.2323349, 0.2337804, 0.2604734, 
    0.3493524, 0.3373525, 0.2389903, 0.2503752, 0.310257, 0.283997, 
    0.2773418, 0.3211859, 0.2661716, 0.2543821, 0.2832943,
  0.2129921, 0.2625791, 0.2463419, 0.232958, 0.2364886, 0.1907316, 0.1839957, 
    0.2190587, 0.178292, 0.2037052, 0.2626095, 0.2026441, 0.2225985, 
    0.188244, 0.1253371, 0.1180767, 0.1462361, 0.2671563, 0.266786, 0.26172, 
    0.2028787, 0.1539979, 0.2455971, 0.152129, 0.07866377, 0.1743234, 
    0.2211225, 0.1587646, 0.1739648,
  0.1268626, 0.118289, 0.04664176, 0.0790024, 0.1054405, 0.06466082, 
    0.1294428, 0.09206687, 0.06590017, 0.1005416, 0.08992516, 0.05023473, 
    0.1381629, 0.2124906, 0.1016468, 0.06208232, 0.1978598, 0.1432752, 
    0.08552683, 0.1132926, 0.08808031, 0.1158162, 0.09388781, 0.03955109, 
    0.06200012, 0.06549332, 0.02795394, 0.08491915, 0.1651652,
  0.01348691, 0.002253021, 0.01674615, 0.01345481, 0.05409918, 0.07822037, 
    0.09498418, 0.04693845, 0.007179865, 0.01527588, 0.0247942, 0.02360552, 
    0.09368303, 0.1072963, 0.03613862, 0.04552992, 0.1021878, 0.09458143, 
    0.1266955, 0.1141872, 0.06902659, 0.1302271, 0.05628889, 0.0002823484, 
    0.01507364, 0.03927293, 0.07190213, 0.04052798, 0.05364473,
  0.005244348, 0.07111364, 0.02223649, 0.03029091, 0.1551062, 0.017501, 
    0.08369891, 0.05080077, 0.01937897, 0.001938267, 0.05066665, 0.01562139, 
    0.02719724, 0.06710777, 0.05315069, 0.1454009, 0.06798471, 0.04992256, 
    0.1141258, 0.05481265, 0.09552544, 0.008401642, -1.657827e-06, 
    0.0001834329, 0.0551807, 0.1004093, 0.07210823, 0.03695612, 0.008004633,
  0.001418924, 0.06968707, 0.2659564, 0.09469973, 0.02576401, 0.04367805, 
    0.03792516, 0.04064802, 0.06746446, 0.01031901, 0.08879641, 0.04367388, 
    0.0578086, 0.02062277, 0.05212207, 0.04425069, 0.08000324, 0.07747642, 
    0.03668941, 0.013103, 0.0004975105, -0.001218327, 0.000201349, 0.2104865, 
    0.1944203, 0.1130278, 0.01117198, 0.001871688, 0.001374294,
  0.001714181, 0.01050529, 0.01043979, 0.03507696, 0.002527281, 0.009242062, 
    0.007481053, 0.008857416, 0.09820591, 0.164262, 0.04203395, 0.02534649, 
    0.03071147, 0.02405949, 0.01916733, 0.04307269, 0.03096554, 0.01240076, 
    0.005649502, 0.01741024, 0.02508063, 0.02722214, 0.09291092, 0.1189375, 
    0.1474449, 0.09014007, 0.02633298, 0.01309744, 0.00365058,
  -1.833077e-05, 5.294469e-07, 8.373266e-07, 0.1027219, 0.0005206715, 
    0.00213719, 0.009551597, 0.07508374, 0.019107, 0.04895074, 0.1322627, 
    0.06447, 0.04399038, 0.03890429, 0.02257279, 0.04794281, 0.02890539, 
    0.008584286, 0.07672095, 0.06704895, 0.04722119, 0.01316335, 0.01668445, 
    0.01044937, 0.01736408, 9.756978e-06, 7.186411e-08, 1.219452e-07, 
    0.0006099474,
  1.564637e-07, 3.256783e-07, -6.707627e-06, -6.882973e-07, 1.758961e-08, 
    4.306233e-07, 0.0004917846, 0.0001602479, 0.02674257, 0.02500053, 
    0.001899628, 0.02606919, 0.01886257, 0.01957623, 0.01164049, 0.01661871, 
    0.0366766, 0.004305927, 0.03816051, 0.0226157, 5.765441e-06, 0.05907869, 
    0.02361178, 0.05293238, 0.007729825, 0.03156391, -1.627636e-05, 
    2.011453e-08, 5.912379e-08,
  4.478578e-07, 0.002171825, 0.03973309, 0.0213531, 0.06540838, 0.0002512866, 
    -0.002007635, 0.05985484, 0.1254172, 0.1806606, 0.1621573, 0.1344899, 
    0.1307193, 0.1062469, 0.07503141, 0.08635432, 0.07202013, 0.08172631, 
    0.03016913, 0.02375825, 0.01748326, 0.06032388, 0.09833858, 0.04802943, 
    0.09262123, 0.08078393, 0.03248208, 0.005656552, 3.698144e-05,
  0.004159347, 0.05792434, 0.1138742, 0.1694875, 0.06725465, 0.03803497, 
    0.2222625, 0.02201062, 0.003766448, 0.04206897, 0.1049848, 0.07197475, 
    0.1458749, 0.1998756, 0.1686047, 0.146348, 0.1272701, 0.1639184, 
    0.1830896, 0.1751674, 0.1141863, 0.1671393, 0.204174, 0.2031143, 
    0.2100944, 0.3095207, 0.08731788, 0.06248135, 0.02429041,
  0.1219833, 0.2648331, 0.2418415, 0.170767, 0.2380466, 0.1689098, 0.1574114, 
    0.1163138, 0.09112758, 0.07500909, 0.05516811, 0.1131618, 0.1217589, 
    0.2094468, 0.3186275, 0.2780744, 0.2522678, 0.2758509, 0.2132151, 
    0.1942565, 0.1480422, 0.10033, 0.1653064, 0.2419634, 0.137187, 0.2378999, 
    0.2003547, 0.1505717, 0.1546195,
  0.2862427, 0.3208343, 0.2183599, 0.3073853, 0.3742292, 0.2312598, 
    0.2544746, 0.2329142, 0.2652323, 0.3861386, 0.2914452, 0.1750595, 
    0.2717368, 0.3112875, 0.3153821, 0.2255282, 0.1898846, 0.3412795, 
    0.3777706, 0.1535531, 0.0845267, 0.205826, 0.1873602, 0.432038, 
    0.1690989, 0.153982, 0.1961605, 0.3577203, 0.2662654,
  0.2393909, 0.1838085, 0.3012541, 0.3092442, 0.3019961, 0.1923954, 
    0.2310804, 0.3559523, 0.241265, 0.2599758, 0.2361535, 0.1938827, 
    0.2243223, 0.1524671, 0.1244538, 0.2145063, 0.07876766, 0.1211843, 
    0.06461412, 0.1137684, 0.1446743, 0.09613591, 0.1688197, 0.1065016, 
    0.2882898, 0.4536432, 0.2931458, 0.3767099, 0.2296382,
  0.0612152, 0.1507619, 0.1770146, 0.2073627, 0.1482997, 0.1853294, 
    0.2564974, 0.3625211, 0.3339002, 0.2655824, 0.1673651, 0.1417584, 
    0.1361898, 0.1091953, 0.1973664, 0.2006343, 0.2091942, 0.1182667, 
    0.1201497, 0.06905368, 0.0872141, 0.1306091, 0.1118719, 0.09519365, 
    0.1568951, 0.1597334, 0.1801952, 0.07146858, 0.07730092,
  0.2285265, 0.2252701, 0.2220137, 0.2187573, 0.215501, 0.2122446, 0.2089882, 
    0.2791836, 0.288071, 0.2969585, 0.3058459, 0.3147334, 0.3236208, 
    0.3325083, 0.3116772, 0.3165931, 0.321509, 0.3264249, 0.3313408, 
    0.3362567, 0.3411726, 0.2978101, 0.2872632, 0.2767162, 0.2661693, 
    0.2556223, 0.2450753, 0.2345283, 0.2311316,
  0.3632489, 0.3423707, 0.11327, 0.03186522, 0.02278268, 0.03008545, 
    0.02573099, 0.01793945, 0.01294091, 0.01164576, 0.0419769, 0.116599, 
    0.2870525, 0.3316834, 0.2698842, 0.1775374, 0.2769314, 0.3302407, 
    0.3171429, 0.236104, 0.2567428, 0.3657499, 0.2943103, 0.276654, 
    0.3678409, 0.3598498, 0.5737269, 0.5480472, 0.3947706,
  0.1461193, 0.1945245, 0.3152439, 0.3269175, 0.1078739, 0.07103604, 
    0.305184, 0.2475339, 0.2777878, 0.3488165, 0.3809364, 0.1785589, 
    0.1751153, 0.4558686, 0.4049732, 0.3221493, 0.3154709, 0.2726108, 
    0.2854969, 0.2607896, 0.2669437, 0.2065145, 0.263526, 0.3630183, 
    0.3870704, 0.347039, 0.3472473, 0.4168386, 0.2382956,
  0.2112089, 0.2701056, 0.2830469, 0.3266552, 0.2590874, 0.2681697, 
    0.3470006, 0.303495, 0.3436737, 0.3332546, 0.2749192, 0.3208638, 
    0.3343256, 0.2415842, 0.2634995, 0.2318656, 0.2560318, 0.2414917, 
    0.3695221, 0.3548534, 0.2517713, 0.2856831, 0.3438894, 0.2892473, 
    0.2788846, 0.2897921, 0.2694079, 0.2780361, 0.300685,
  0.2076654, 0.241126, 0.2505435, 0.2509944, 0.2376071, 0.1956384, 0.2061071, 
    0.2228325, 0.1903873, 0.2156442, 0.2380231, 0.2145166, 0.2306196, 
    0.2216723, 0.1126877, 0.1235337, 0.161829, 0.3222865, 0.3019521, 
    0.2855763, 0.1985484, 0.1752798, 0.2636752, 0.1708188, 0.06891199, 
    0.1647773, 0.2282456, 0.1701254, 0.1837569,
  0.1323885, 0.1344417, 0.05503702, 0.08895471, 0.1137563, 0.06822386, 
    0.1168761, 0.09876645, 0.09608097, 0.09549531, 0.09475399, 0.08557364, 
    0.1260258, 0.1922438, 0.1192775, 0.08216508, 0.2118303, 0.1573111, 
    0.09017023, 0.1193978, 0.07448714, 0.1405723, 0.1243766, 0.04554428, 
    0.04138197, 0.07410429, 0.05446187, 0.0980619, 0.175835,
  0.01263103, 0.007981991, 0.01520768, 0.02403769, 0.07145574, 0.07975665, 
    0.1043007, 0.04651352, 0.01730113, 0.01439018, 0.02253831, 0.001946343, 
    0.1034694, 0.1071688, 0.04691669, 0.04982077, 0.1339922, 0.1088816, 
    0.1135701, 0.1261015, 0.06465562, 0.1497085, 0.05864326, 5.665616e-05, 
    0.01040762, 0.04088192, 0.07551698, 0.04509635, 0.05357832,
  0.009827766, 0.06157843, 0.0233466, 0.02868606, 0.1439102, 0.02126442, 
    0.07748863, 0.0740061, 0.0249175, 0.002789701, 0.03523768, 0.006295725, 
    0.02397615, 0.06614874, 0.04804875, 0.1422163, 0.06672166, 0.04247387, 
    0.1081346, 0.04841008, 0.09160393, 0.03392395, -2.062198e-05, 
    0.0002831588, 0.05966391, 0.09108483, 0.06066383, 0.0593195, 0.02598451,
  0.002312954, 0.04305961, 0.2340235, 0.09192232, 0.02711629, 0.03533743, 
    0.03595039, 0.03750157, 0.05693309, 0.01197943, 0.08491622, 0.041397, 
    0.05626482, 0.02114652, 0.03972501, 0.03487743, 0.07076609, 0.06483786, 
    0.03656641, 0.01882276, 0.008679633, -3.352318e-06, 0.006495391, 
    0.1975667, 0.168559, 0.09818427, 0.02045037, 0.002948134, 0.002839424,
  0.001517455, 0.008252488, 0.008964444, 0.0223768, 0.004297582, 0.01377961, 
    0.00814012, 0.01265435, 0.09651319, 0.1744839, 0.04033963, 0.02420332, 
    0.0281464, 0.02309946, 0.01817532, 0.0359164, 0.03663436, 0.01652321, 
    0.01642034, 0.01718402, 0.02709814, 0.03180153, 0.09096199, 0.09282933, 
    0.146048, 0.08279447, 0.02756469, 0.01520534, 0.003372339,
  -4.141409e-06, 1.657601e-07, 2.42658e-07, 0.03855503, 0.003200784, 
    0.002668367, 0.01264492, 0.05807656, 0.01544719, 0.05409624, 0.1246322, 
    0.07016821, 0.05085541, 0.03525027, 0.02577668, 0.04528099, 0.02804727, 
    0.0165609, 0.09384493, 0.07370003, 0.04385955, 0.01529051, 0.03496355, 
    0.01652297, 0.01876758, 0.0002083593, 3.682869e-07, 9.169403e-09, 
    0.0002669482,
  9.689077e-08, 1.093115e-07, -3.375308e-06, -7.013743e-06, 5.950742e-09, 
    9.027838e-07, 6.985189e-05, 0.0002149686, 0.003003453, 0.02160387, 
    0.004080118, 0.03113598, 0.02186279, 0.02420998, 0.01449666, 0.02405639, 
    0.03510762, 0.02354952, 0.04662354, 0.02137163, 2.891064e-06, 0.07703532, 
    0.01887076, 0.05247347, 0.03047412, 0.03014061, 0.0009312545, 
    -3.044778e-09, 2.921494e-08,
  1.678122e-07, 0.007781891, 0.04313662, 0.01210446, 0.03868058, 
    -2.789443e-05, -0.001695793, 0.05128909, 0.09792479, 0.1566833, 
    0.1520021, 0.1409822, 0.1292462, 0.1051279, 0.08398134, 0.09497492, 
    0.1182117, 0.09083591, 0.04449631, 0.0322411, 0.01435765, 0.07921268, 
    0.08618771, 0.05521583, 0.1117345, 0.09177745, 0.03593231, 0.005322214, 
    1.813018e-05,
  0.004844736, 0.05511192, 0.1092657, 0.1853086, 0.06270263, 0.04985985, 
    0.202355, 0.02447299, 0.001580449, 0.05595762, 0.08675598, 0.08667767, 
    0.1763322, 0.2278327, 0.194087, 0.1569386, 0.1480312, 0.1957919, 
    0.2112005, 0.1724426, 0.1171991, 0.1899544, 0.2112218, 0.1765963, 
    0.2590365, 0.3233932, 0.125827, 0.06958935, 0.02219866,
  0.1330965, 0.2605357, 0.2401664, 0.1441144, 0.1672806, 0.1167498, 
    0.1149249, 0.1325003, 0.09312684, 0.04956611, 0.04463952, 0.1166489, 
    0.1025119, 0.2713037, 0.3351158, 0.258387, 0.248414, 0.2783788, 
    0.2113367, 0.1807015, 0.1308939, 0.093053, 0.1417339, 0.2334857, 
    0.1314052, 0.2634142, 0.2285862, 0.1732092, 0.1785761,
  0.274619, 0.3113652, 0.2572435, 0.2812523, 0.3156739, 0.2072656, 0.2745276, 
    0.310484, 0.2896255, 0.3927393, 0.318442, 0.1905876, 0.2641234, 
    0.2896471, 0.296849, 0.2218506, 0.1559647, 0.3372436, 0.350119, 
    0.1589225, 0.08378334, 0.1561085, 0.1918306, 0.4122635, 0.1852987, 
    0.1699554, 0.2653532, 0.3551658, 0.3132832,
  0.2369605, 0.2040177, 0.2448596, 0.2875177, 0.2574599, 0.2156672, 
    0.2624504, 0.3474934, 0.2306479, 0.2826635, 0.2555875, 0.1810439, 
    0.2043114, 0.08967368, 0.1542881, 0.1533399, 0.08510713, 0.1175256, 
    0.06537346, 0.1113531, 0.1112417, 0.09249183, 0.1864265, 0.1143521, 
    0.2705487, 0.5281039, 0.3649959, 0.3415942, 0.2161508,
  0.06730755, 0.1664041, 0.1853381, 0.2244756, 0.189087, 0.2323415, 
    0.2713007, 0.3806784, 0.3323629, 0.2580196, 0.1747455, 0.1216598, 
    0.1232297, 0.1678446, 0.2186248, 0.1840189, 0.2091729, 0.100524, 
    0.1171836, 0.05419908, 0.08223833, 0.1278491, 0.1167372, 0.10263, 
    0.1364361, 0.1529684, 0.1875337, 0.08504287, 0.1144607,
  0.3042807, 0.3001232, 0.2959658, 0.2918083, 0.2876508, 0.2834933, 
    0.2793358, 0.3396861, 0.349467, 0.359248, 0.369029, 0.3788099, 0.3885909, 
    0.3983718, 0.3858623, 0.3902589, 0.3946556, 0.3990522, 0.4034489, 
    0.4078455, 0.4122422, 0.394963, 0.3849429, 0.3749228, 0.3649026, 
    0.3548825, 0.3448624, 0.3348423, 0.3076067,
  0.342408, 0.3600067, 0.2477805, 0.03915924, 0.03202185, 0.03489638, 
    0.03298906, 0.01553867, 0.01054582, 0.01016696, 0.07281701, 0.129438, 
    0.3119286, 0.2898817, 0.2127975, 0.2028375, 0.3019084, 0.3418905, 
    0.362819, 0.2443832, 0.3057082, 0.3733386, 0.3079605, 0.2825462, 
    0.3983274, 0.432219, 0.5734386, 0.5109123, 0.3873539,
  0.1734843, 0.2028964, 0.3057694, 0.3352035, 0.1073888, 0.08536555, 
    0.3549838, 0.2587341, 0.2912581, 0.3756413, 0.3691526, 0.1658914, 
    0.1891361, 0.4614157, 0.4534077, 0.3859715, 0.3817888, 0.3401602, 
    0.3777525, 0.2924497, 0.2984301, 0.1970374, 0.2806749, 0.4186222, 
    0.3535463, 0.404906, 0.3622786, 0.4011928, 0.3179031,
  0.2528444, 0.2913645, 0.2533208, 0.4002036, 0.2887705, 0.2799053, 
    0.3767803, 0.3836107, 0.3621676, 0.4254127, 0.2797392, 0.336314, 
    0.3928965, 0.2662838, 0.2737574, 0.2627814, 0.2726796, 0.2698391, 
    0.434117, 0.3898204, 0.2744873, 0.3626852, 0.4039457, 0.3593691, 
    0.2890697, 0.3194454, 0.2838984, 0.2888562, 0.2896912,
  0.2345231, 0.2602888, 0.2982891, 0.3070515, 0.2530838, 0.221363, 0.2429237, 
    0.2822629, 0.2064873, 0.241556, 0.2408512, 0.218052, 0.2452613, 
    0.2313519, 0.1038851, 0.1209304, 0.1720542, 0.3739733, 0.3142768, 
    0.3061776, 0.2241311, 0.2059859, 0.2561078, 0.1868526, 0.07291061, 
    0.1669391, 0.2442944, 0.2249984, 0.2108813,
  0.1681208, 0.155564, 0.07754764, 0.1160124, 0.1216808, 0.1036258, 
    0.1679063, 0.1403337, 0.1189909, 0.08562043, 0.1262135, 0.1142933, 
    0.1243934, 0.1722209, 0.1410524, 0.1091338, 0.242126, 0.1974645, 
    0.1083516, 0.1538375, 0.0774993, 0.1678067, 0.1576381, 0.0530717, 
    0.03740557, 0.09919763, 0.09851409, 0.1190422, 0.1753152,
  0.03501154, 0.0124647, 0.01895416, 0.04231596, 0.09516542, 0.09737078, 
    0.1292644, 0.07190786, 0.03728829, 0.01698246, 0.02591796, -3.376617e-05, 
    0.08510137, 0.1106657, 0.04619057, 0.05722526, 0.1367489, 0.1363592, 
    0.1213362, 0.1229388, 0.06480987, 0.1602427, 0.08262753, -2.619768e-05, 
    0.008672114, 0.04438616, 0.0720152, 0.05613391, 0.05134417,
  0.01117229, 0.05166038, 0.03912365, 0.03078496, 0.1409196, 0.02472808, 
    0.07338937, 0.08417284, 0.03155762, 0.003238463, 0.02392235, 0.002790797, 
    0.02540703, 0.06478398, 0.04478469, 0.123036, 0.06160756, 0.0337904, 
    0.1001581, 0.03885211, 0.05740424, 0.0868098, 0.003702051, 0.0004804034, 
    0.06555483, 0.1141072, 0.04187801, 0.04586528, 0.05804554,
  0.005930852, 0.03155124, 0.1924233, 0.09934173, 0.02509848, 0.0288422, 
    0.03422186, 0.02913145, 0.04796463, 0.01541533, 0.08336115, 0.04261633, 
    0.06003884, 0.02393388, 0.03216944, 0.02865241, 0.05914529, 0.03512267, 
    0.0341161, 0.01984944, 0.00986341, 0.0027855, 0.02146106, 0.1785395, 
    0.1497651, 0.08134598, 0.03009092, 0.01055458, 0.00739324,
  0.001711566, 0.01050002, 0.008233317, 0.0242288, 0.007235067, 0.0181528, 
    0.01065872, 0.01852957, 0.1003119, 0.1803542, 0.03234028, 0.02433245, 
    0.02595115, 0.02464065, 0.0165923, 0.03394433, 0.03243756, 0.02213987, 
    0.02623315, 0.01891877, 0.02171725, 0.02619717, 0.07460124, 0.07019226, 
    0.1332482, 0.06460803, 0.02595043, 0.018499, 0.00465057,
  -1.44709e-07, 6.76111e-08, 5.897098e-08, 0.0134818, 0.01804918, 
    0.004137222, 0.01988775, 0.04357887, 0.01431857, 0.05564416, 0.1232405, 
    0.0656975, 0.04511373, 0.03714462, 0.02395821, 0.03562045, 0.02889502, 
    0.02924739, 0.1152307, 0.07969863, 0.03706307, 0.01702156, 0.04131273, 
    0.01611108, 0.01865236, 0.002257059, 1.127602e-06, 2.866721e-09, 
    9.412037e-05,
  6.407415e-08, 9.454948e-09, -1.180761e-06, 2.138716e-05, 1.046005e-09, 
    2.594767e-06, 1.661055e-05, 0.0001404148, 0.0003381304, 0.03236457, 
    0.02228303, 0.05831754, 0.02791976, 0.04113336, 0.04448589, 0.01814582, 
    0.04861363, 0.03689676, 0.07638123, 0.02635093, 1.994708e-06, 0.100437, 
    0.01886506, 0.0417994, 0.04832797, 0.06691086, 0.03910908, -8.130676e-06, 
    1.603417e-08,
  8.043747e-08, 0.0116313, 0.04238556, 0.01128599, 0.02714838, -1.951828e-05, 
    -0.001376933, 0.0376499, 0.08007056, 0.1508845, 0.1548581, 0.1912899, 
    0.1845559, 0.1768996, 0.1147187, 0.1756258, 0.1771357, 0.1231284, 
    0.07368775, 0.03823683, 0.007710967, 0.09441439, 0.07578966, 0.1023907, 
    0.1345295, 0.1012131, 0.03663233, 0.006796539, 1.42914e-05,
  0.002709838, 0.05981643, 0.1096451, 0.1947196, 0.06642394, 0.02732624, 
    0.1821384, 0.02660141, 0.001312257, 0.07418738, 0.07193604, 0.1078826, 
    0.2136644, 0.2889767, 0.2245638, 0.1813951, 0.1821765, 0.2208323, 
    0.2419813, 0.1805875, 0.1320885, 0.2071817, 0.2321338, 0.1765425, 
    0.3251401, 0.3279671, 0.145052, 0.09661397, 0.02069647,
  0.1141301, 0.2974915, 0.2630732, 0.2122952, 0.1541871, 0.1404039, 0.105111, 
    0.1258993, 0.0830333, 0.03049223, 0.05634024, 0.0992147, 0.09606881, 
    0.3445993, 0.3573341, 0.2949705, 0.2815432, 0.2800709, 0.2186411, 
    0.1833175, 0.1630785, 0.1208268, 0.1450349, 0.2450621, 0.1393216, 
    0.2881846, 0.2528001, 0.2079824, 0.1777111,
  0.2712075, 0.3143331, 0.304498, 0.3178258, 0.4061565, 0.2635831, 0.2735672, 
    0.2918029, 0.3254466, 0.4448262, 0.3467796, 0.2119964, 0.2582873, 
    0.3231522, 0.3041316, 0.1772333, 0.1321788, 0.3285231, 0.3247609, 
    0.1756635, 0.1161528, 0.1188963, 0.2182386, 0.3684963, 0.2043137, 
    0.1858566, 0.3470815, 0.3706701, 0.3055926,
  0.2289463, 0.2396892, 0.2807119, 0.3565764, 0.271886, 0.2124741, 0.2650821, 
    0.3628298, 0.2227139, 0.2961608, 0.2688664, 0.1789147, 0.216546, 
    0.05640909, 0.1525369, 0.1154715, 0.1521255, 0.1288701, 0.06627104, 
    0.1110903, 0.09908234, 0.0966757, 0.1928319, 0.1139236, 0.2600963, 
    0.5425909, 0.4236912, 0.3156648, 0.2245861,
  0.05919493, 0.1625886, 0.2161357, 0.2417896, 0.169717, 0.2404811, 
    0.2747934, 0.4088815, 0.3454659, 0.2711162, 0.1755217, 0.1024057, 
    0.09842131, 0.1843464, 0.2151601, 0.2312801, 0.2242752, 0.1460791, 
    0.1339272, 0.09063028, 0.1156896, 0.1447203, 0.1339806, 0.1058802, 
    0.1240564, 0.1467429, 0.1847463, 0.1222111, 0.1421323,
  0.3715583, 0.3692498, 0.3669414, 0.3646329, 0.3623244, 0.360016, 0.3577075, 
    0.3759928, 0.3851427, 0.3942926, 0.4034425, 0.4125924, 0.4217422, 
    0.4308921, 0.4578198, 0.4605326, 0.4632455, 0.4659582, 0.468671, 
    0.4713838, 0.4740966, 0.4510046, 0.4414504, 0.4318962, 0.4223419, 
    0.4127877, 0.4032335, 0.3936793, 0.373405,
  0.3142951, 0.3875316, 0.3401209, 0.09784902, 0.04715704, 0.0770342, 
    0.06706024, 0.05215, 0.01468905, 0.02291628, 0.09337619, 0.1713874, 
    0.3299958, 0.2272995, 0.1854682, 0.2217037, 0.2993436, 0.3195569, 
    0.378184, 0.23244, 0.3431641, 0.3717547, 0.3402673, 0.3559991, 0.4104017, 
    0.4267308, 0.5200174, 0.4429104, 0.3828372,
  0.1736813, 0.1802128, 0.334325, 0.3080199, 0.1130495, 0.1039967, 0.3503858, 
    0.272827, 0.3042659, 0.3517577, 0.3401578, 0.1555707, 0.2075133, 
    0.455752, 0.5095982, 0.4599759, 0.5181532, 0.4918557, 0.3858741, 
    0.3207501, 0.2871678, 0.1911783, 0.2309664, 0.4255791, 0.4026433, 
    0.5188212, 0.3791836, 0.5315297, 0.4015035,
  0.3161049, 0.3865359, 0.3237851, 0.3935033, 0.2846855, 0.3337345, 
    0.4344065, 0.4376084, 0.4573242, 0.3927246, 0.3410205, 0.4188207, 
    0.4566296, 0.2976663, 0.3310412, 0.2978113, 0.2969759, 0.3230419, 
    0.4298145, 0.4102097, 0.3250735, 0.382738, 0.3879383, 0.3666697, 
    0.3478253, 0.4132507, 0.3746952, 0.3417268, 0.3038937,
  0.2942943, 0.2975219, 0.3134381, 0.299511, 0.2823311, 0.2499255, 0.2539801, 
    0.2987216, 0.2136805, 0.268224, 0.3134095, 0.2723135, 0.2940045, 
    0.2492793, 0.11984, 0.1815754, 0.2500786, 0.3957029, 0.3074004, 
    0.3245521, 0.2571498, 0.2280874, 0.3002838, 0.1758095, 0.06350729, 
    0.1691867, 0.2607474, 0.2650615, 0.2753926,
  0.1889684, 0.1638102, 0.09972253, 0.1461449, 0.1643879, 0.1365725, 
    0.1840475, 0.1539846, 0.1518879, 0.09890833, 0.1933837, 0.137232, 
    0.1244158, 0.1976953, 0.1878335, 0.1333278, 0.2796023, 0.2268016, 
    0.1299049, 0.1639514, 0.1711686, 0.2074661, 0.1682958, 0.06020983, 
    0.03911371, 0.1343479, 0.1272471, 0.1601634, 0.2479407,
  0.06007139, 0.01284412, 0.0130268, 0.08969954, 0.1148878, 0.1206971, 
    0.1693305, 0.1007075, 0.08662723, 0.04113651, 0.02522421, -3.453451e-05, 
    0.07594881, 0.1254206, 0.08397812, 0.06134603, 0.1393322, 0.1664121, 
    0.1469302, 0.1220633, 0.07178444, 0.1879, 0.1481061, -6.054482e-06, 
    0.0106337, 0.06669129, 0.09349991, 0.076298, 0.05260678,
  0.01227603, 0.0432923, 0.01899312, 0.05305757, 0.1291483, 0.02799172, 
    0.0705725, 0.08627867, 0.05365236, 0.004110879, 0.01537491, 0.001248744, 
    0.03329288, 0.0629241, 0.04207689, 0.09955028, 0.05970171, 0.0300692, 
    0.09103734, 0.04213304, 0.0475999, 0.1301144, 0.0739364, 0.000733444, 
    0.07931749, 0.1685994, 0.05043799, 0.04255452, 0.05701261,
  0.01718337, 0.03660427, 0.1479053, 0.1178963, 0.02564466, 0.02893741, 
    0.03579468, 0.02688205, 0.04218838, 0.02334365, 0.08100116, 0.03780315, 
    0.06791162, 0.02998347, 0.02887042, 0.02768871, 0.04959104, 0.03313841, 
    0.03422912, 0.02336897, 0.0132602, 0.01744322, 0.04295417, 0.1749921, 
    0.1284033, 0.06837796, 0.04587927, 0.03952636, 0.03271633,
  0.002770984, 0.01360774, 0.006356446, 0.02082377, 0.01220112, 0.02533947, 
    0.01716507, 0.02442634, 0.09958386, 0.1600775, 0.03170376, 0.02551179, 
    0.02763975, 0.02714597, 0.01781914, 0.03087293, 0.02949027, 0.02447786, 
    0.01947572, 0.01784083, 0.02048337, 0.02649591, 0.05546454, 0.05635899, 
    0.1325449, 0.05080607, 0.02529922, 0.01985506, 0.008872871,
  -4.859208e-07, 3.70159e-08, 2.069342e-08, 0.002323153, 0.01479164, 
    0.01198066, 0.02379199, 0.03577702, 0.01209965, 0.05519856, 0.1248029, 
    0.05740713, 0.03716481, 0.03381021, 0.02276037, 0.03164655, 0.0284941, 
    0.0371486, 0.1237766, 0.08736145, 0.03524883, 0.02111504, 0.04064813, 
    0.02405341, 0.02526844, 0.02130785, 0.0001619083, 8.773732e-10, 
    4.091813e-05,
  3.581582e-08, 8.815018e-09, -5.035535e-08, 0.0005767414, 3.031273e-10, 
    4.24462e-05, -4.913274e-07, -7.720162e-06, 1.137275e-05, 0.05839211, 
    0.04878357, 0.1060782, 0.07033061, 0.06616864, 0.06715133, 0.03222161, 
    0.07075972, 0.06366219, 0.09318179, 0.1126389, 9.446339e-07, 0.1205903, 
    0.0561635, 0.06127153, 0.09816302, 0.09062259, 0.0807106, 9.169098e-05, 
    1.072045e-08,
  3.962101e-08, 0.007241115, 0.05789099, 0.00894432, 0.01741922, 
    8.905682e-07, -0.001116302, 0.02652603, 0.0746107, 0.1491913, 0.1844492, 
    0.1740863, 0.153059, 0.1557272, 0.2267583, 0.2090417, 0.1542884, 
    0.2069919, 0.1301982, 0.06700431, 0.006053585, 0.1253877, 0.07326027, 
    0.1902129, 0.1456283, 0.1125936, 0.03579824, 0.01596662, 1.339364e-05,
  0.0005950892, 0.03699462, 0.1144874, 0.2359297, 0.09580491, 0.02189968, 
    0.1449503, 0.01795754, 0.00145311, 0.04627926, 0.05742907, 0.1001215, 
    0.2218808, 0.2600103, 0.1880332, 0.1917005, 0.2070395, 0.2190177, 
    0.2701432, 0.1825767, 0.1148168, 0.2318615, 0.2529817, 0.1970328, 
    0.3660555, 0.3512735, 0.1467172, 0.1455838, 0.02318064,
  0.1058385, 0.3154019, 0.2246609, 0.2279036, 0.1521778, 0.1821035, 
    0.1132414, 0.1298041, 0.06911856, 0.02488083, 0.01495655, 0.09353209, 
    0.07705193, 0.394668, 0.3544656, 0.3209071, 0.2929156, 0.2731044, 
    0.2297507, 0.2059434, 0.1790009, 0.113654, 0.1272717, 0.3061879, 
    0.1560561, 0.3625482, 0.316667, 0.2624269, 0.1979329,
  0.2836032, 0.3078116, 0.2892626, 0.3001604, 0.4371047, 0.27657, 0.3105812, 
    0.2619587, 0.3500385, 0.4569038, 0.3634157, 0.2219327, 0.2375877, 
    0.3501429, 0.4183507, 0.2375556, 0.1461364, 0.3246128, 0.3070222, 
    0.1598705, 0.1155799, 0.1802529, 0.2133967, 0.3598655, 0.3516768, 
    0.2320883, 0.3677546, 0.3635059, 0.2780455,
  0.2448129, 0.3035243, 0.3430406, 0.448823, 0.2769125, 0.222459, 0.2699878, 
    0.371686, 0.2671231, 0.3084987, 0.274395, 0.1706464, 0.2196655, 
    0.09527298, 0.1428852, 0.08246402, 0.1215688, 0.168952, 0.06830925, 
    0.129209, 0.1023082, 0.1521886, 0.2128873, 0.1282062, 0.2324481, 0.52255, 
    0.4618984, 0.3096351, 0.2260329,
  0.09820673, 0.234408, 0.2791788, 0.2577484, 0.2184541, 0.2703308, 
    0.3128983, 0.4145845, 0.367582, 0.3008989, 0.1975657, 0.1167196, 
    0.1074439, 0.1779913, 0.2606298, 0.2336224, 0.2088773, 0.1578324, 
    0.1139658, 0.1117604, 0.1199003, 0.1608137, 0.1418249, 0.09764045, 
    0.1060754, 0.1267656, 0.1878, 0.1316877, 0.1618471,
  0.4237208, 0.4234163, 0.4231118, 0.4228072, 0.4225027, 0.4221982, 
    0.4218937, 0.4195724, 0.4269175, 0.4342626, 0.4416077, 0.4489529, 
    0.456298, 0.4636431, 0.4922089, 0.4923983, 0.4925876, 0.492777, 
    0.4929664, 0.4931557, 0.4933451, 0.459016, 0.451786, 0.4445561, 
    0.4373261, 0.4300961, 0.4228661, 0.4156361, 0.4239644,
  0.2903997, 0.4068105, 0.3840458, 0.1499677, 0.08281808, 0.1022293, 
    0.1344891, 0.09407662, 0.01406528, 0.03163778, 0.1119608, 0.2062263, 
    0.3147834, 0.1856736, 0.2032945, 0.2029082, 0.2777569, 0.2717761, 
    0.274819, 0.2912374, 0.361618, 0.4055172, 0.3543775, 0.361636, 0.4616736, 
    0.4442229, 0.4485595, 0.3565775, 0.3501268,
  0.1906446, 0.1836646, 0.3208746, 0.2508774, 0.1283452, 0.1443024, 
    0.2914408, 0.3088028, 0.3263368, 0.3484078, 0.329392, 0.1508867, 
    0.2346123, 0.432321, 0.4672534, 0.4052018, 0.5029774, 0.4178985, 
    0.4375431, 0.3633725, 0.3378136, 0.2604159, 0.2268022, 0.4305277, 
    0.4463938, 0.536433, 0.6221992, 0.6139204, 0.4767886,
  0.4158467, 0.377064, 0.3467583, 0.3847836, 0.317657, 0.4206303, 0.4626195, 
    0.5113959, 0.5270188, 0.3881422, 0.3731728, 0.4463298, 0.4673776, 
    0.4041184, 0.3650184, 0.3234181, 0.3576112, 0.3890706, 0.4974616, 
    0.3872593, 0.3630864, 0.3468086, 0.3827207, 0.4177828, 0.4376218, 
    0.5019681, 0.4973694, 0.5185786, 0.4246536,
  0.3385297, 0.3333271, 0.3283885, 0.2876715, 0.3011793, 0.2718794, 0.262361, 
    0.3040786, 0.2535607, 0.2876196, 0.3393129, 0.266727, 0.2632722, 
    0.2668025, 0.1392645, 0.1976938, 0.3947848, 0.4097972, 0.3796933, 
    0.3602499, 0.3370257, 0.2977151, 0.3126137, 0.1766988, 0.04616076, 
    0.1853414, 0.2750303, 0.2750303, 0.3599854,
  0.2018782, 0.2307318, 0.1878893, 0.2077743, 0.1868702, 0.1605648, 0.224081, 
    0.2886024, 0.2336668, 0.2114464, 0.2706776, 0.1403696, 0.110552, 
    0.2308052, 0.1573887, 0.1644027, 0.2940387, 0.2596289, 0.1779583, 
    0.1659909, 0.2327947, 0.2148914, 0.1415231, 0.07692017, 0.05250265, 
    0.1715216, 0.1292808, 0.1690184, 0.2410787,
  0.1047718, 0.01873258, 0.005487948, 0.1229337, 0.1421003, 0.1301744, 
    0.1750002, 0.1477994, 0.2111855, 0.06197075, 0.03193117, -6.739717e-05, 
    0.06354748, 0.1426814, 0.07732162, 0.04917018, 0.160831, 0.2024122, 
    0.1888337, 0.1715784, 0.0795826, 0.1983317, 0.1270862, 9.239512e-05, 
    0.006192877, 0.05843002, 0.1013376, 0.08189144, 0.06865884,
  0.08020548, 0.03155131, 0.01328292, 0.06473647, 0.1165619, 0.03622739, 
    0.07575534, 0.08536937, 0.09638823, 0.01603322, 0.009639976, 
    0.0004117994, 0.06036199, 0.07971632, 0.06049201, 0.1177846, 0.06164814, 
    0.03466554, 0.1138374, 0.05620273, 0.05361185, 0.1027604, 0.3178749, 
    0.001047683, 0.08021532, 0.1639505, 0.05625755, 0.04941426, 0.05842371,
  0.05529225, 0.03953844, 0.1089452, 0.1172387, 0.03408624, 0.03347452, 
    0.04503787, 0.0302221, 0.04210619, 0.03051687, 0.07706811, 0.03501683, 
    0.07197178, 0.04286385, 0.02584769, 0.04368058, 0.04227375, 0.05661593, 
    0.04230262, 0.04153401, 0.02648778, 0.03852414, 0.08527008, 0.1575284, 
    0.09875426, 0.05491184, 0.06863638, 0.1260228, 0.1072518,
  0.007133407, 0.01133203, 0.004193009, 0.01576746, 0.0282792, 0.03670033, 
    0.06438962, 0.04560751, 0.09786128, 0.1359623, 0.03252841, 0.0279845, 
    0.03238959, 0.03074254, 0.04895978, 0.03160648, 0.02603656, 0.02451318, 
    0.01873895, 0.01872303, 0.02512406, 0.02618929, 0.03313299, 0.03487018, 
    0.1119248, 0.04646863, 0.02990905, 0.02567083, 0.01534473,
  -7.296007e-07, 2.526466e-08, 8.514738e-09, 3.396436e-05, 0.03997933, 
    0.06609368, 0.02255551, 0.05967884, 0.01331057, 0.07699484, 0.1252076, 
    0.05083014, 0.03480427, 0.04230536, 0.02594615, 0.03820448, 0.03341488, 
    0.04256108, 0.1205122, 0.08964872, 0.06143537, 0.04140127, 0.03685063, 
    0.03678776, 0.06104923, 0.1166308, 0.004135809, -2.718737e-10, 
    2.179895e-05,
  1.91757e-08, 5.526343e-10, -1.004068e-08, 0.0003705977, 2.607212e-10, 
    9.140749e-06, -3.86752e-07, -8.859846e-05, -1.711491e-05, 0.06953258, 
    0.08393537, 0.124825, 0.1108162, 0.09949955, 0.05651169, 0.05351484, 
    0.1279239, 0.07837801, 0.1876792, 0.1663764, -5.11333e-07, 0.129581, 
    0.05543499, 0.05292505, 0.08592676, 0.08594517, 0.1045478, 0.001415358, 
    8.4771e-09,
  1.841415e-08, 0.003849237, 0.04646854, 0.01569936, 0.01134538, 
    1.649916e-06, -0.0008872077, 0.01665978, 0.0705665, 0.1598239, 0.1641145, 
    0.1462186, 0.1420455, 0.1756184, 0.2058157, 0.2588245, 0.2039948, 
    0.2251211, 0.1578686, 0.05302882, 0.009128997, 0.1612618, 0.07851467, 
    0.176352, 0.1410073, 0.1232436, 0.06217845, 0.0212394, 8.76251e-06,
  -0.0007075482, 0.02869071, 0.1011519, 0.2177279, 0.07139535, 0.02291409, 
    0.1185898, 0.008370088, 0.002458444, 0.01781473, 0.05080401, 0.08035185, 
    0.1989874, 0.1979155, 0.1590889, 0.2221947, 0.2033329, 0.256251, 
    0.2777669, 0.1871482, 0.0930325, 0.2258705, 0.2374979, 0.216566, 
    0.3488853, 0.3374423, 0.1760475, 0.1785079, 0.06955296,
  0.1207696, 0.3502082, 0.2310257, 0.2665855, 0.2008253, 0.1723818, 
    0.1529699, 0.1446768, 0.04840602, 0.01729147, 0.006192173, 0.09080978, 
    0.09767738, 0.3720693, 0.2298522, 0.2952151, 0.2381474, 0.2729886, 
    0.2191285, 0.2241476, 0.1537893, 0.09901735, 0.1235038, 0.3077756, 
    0.1403014, 0.427897, 0.3581916, 0.2577551, 0.2007853,
  0.2698211, 0.2900952, 0.2847669, 0.2943976, 0.5120142, 0.3390354, 
    0.2970269, 0.2393116, 0.3076272, 0.4220208, 0.3188453, 0.208515, 
    0.2297425, 0.3310924, 0.5702435, 0.2537559, 0.1639242, 0.3132434, 
    0.2901211, 0.1363705, 0.120119, 0.1815927, 0.2505633, 0.3724059, 
    0.5801396, 0.1339211, 0.2361936, 0.3185913, 0.2377754,
  0.2695712, 0.2239646, 0.3431697, 0.4390846, 0.2606928, 0.215281, 0.2629552, 
    0.386382, 0.3065575, 0.3278029, 0.3133186, 0.1581315, 0.2219036, 
    0.1342686, 0.2157484, 0.09787165, 0.1269733, 0.1802133, 0.08428989, 
    0.1614556, 0.1508819, 0.1791127, 0.2375083, 0.1301798, 0.2335498, 
    0.5104893, 0.4773434, 0.2945381, 0.314577,
  0.1012726, 0.2991294, 0.2772453, 0.2449627, 0.2375076, 0.3070575, 
    0.3288562, 0.4295792, 0.3818498, 0.3408858, 0.2600454, 0.1513483, 
    0.1649531, 0.2169217, 0.2692397, 0.2047084, 0.2302974, 0.1948787, 
    0.1475339, 0.1333761, 0.1358505, 0.1810401, 0.1438251, 0.09048068, 
    0.09838233, 0.115243, 0.1957151, 0.1495482, 0.1858426,
  0.4688378, 0.469766, 0.4706942, 0.4716223, 0.4725505, 0.4734787, 0.4744069, 
    0.452673, 0.4596007, 0.4665285, 0.4734562, 0.4803839, 0.4873116, 
    0.4942393, 0.5007465, 0.4969566, 0.4931667, 0.4893768, 0.4855869, 
    0.481797, 0.478007, 0.4523965, 0.4483305, 0.4442645, 0.4401986, 
    0.4361326, 0.4320666, 0.4280006, 0.4680952,
  0.3047067, 0.4441353, 0.4229309, 0.1741353, 0.1080248, 0.1377142, 
    0.1797576, 0.1340829, 0.01974818, 0.04502572, 0.1520784, 0.2327211, 
    0.3297672, 0.1386382, 0.24769, 0.1985885, 0.262925, 0.2571861, 0.2107564, 
    0.3356282, 0.3960576, 0.4129839, 0.4004021, 0.3344049, 0.4646302, 
    0.5125348, 0.4558474, 0.2973675, 0.365232,
  0.2052137, 0.1599326, 0.3162629, 0.1568876, 0.1500304, 0.1648245, 
    0.2437598, 0.2928615, 0.3738895, 0.3455234, 0.3367869, 0.1445453, 
    0.2386152, 0.3619315, 0.3545487, 0.4036499, 0.4136778, 0.394916, 
    0.429398, 0.4023266, 0.3666577, 0.2831895, 0.2273596, 0.4285897, 
    0.4804598, 0.4102161, 0.4744672, 0.5733131, 0.3746251,
  0.3372297, 0.2894879, 0.2929543, 0.3490636, 0.3226367, 0.4199911, 
    0.4849884, 0.5088764, 0.5084633, 0.3923453, 0.3324551, 0.4081473, 
    0.5326618, 0.4520885, 0.3942017, 0.3729749, 0.3907089, 0.4488012, 
    0.5358442, 0.411753, 0.4053111, 0.3671178, 0.4125089, 0.4107207, 
    0.4235251, 0.5416858, 0.5146547, 0.5447888, 0.4283074,
  0.3640115, 0.3485361, 0.3514259, 0.3360555, 0.3070337, 0.3573158, 0.299352, 
    0.311602, 0.2764459, 0.3318485, 0.3614519, 0.2788194, 0.2615051, 
    0.339502, 0.1609276, 0.2349591, 0.4026367, 0.4701967, 0.3648687, 
    0.3638837, 0.293937, 0.2839174, 0.2804239, 0.1879321, 0.04703326, 
    0.2104444, 0.3000257, 0.3710048, 0.4211514,
  0.2391436, 0.2879357, 0.1710171, 0.2051292, 0.2568767, 0.2139314, 
    0.2373019, 0.3202475, 0.2515623, 0.2786658, 0.218307, 0.132725, 
    0.07521765, 0.1984088, 0.1686772, 0.1096047, 0.2472892, 0.2359473, 
    0.1692171, 0.1667213, 0.1753094, 0.1556818, 0.1567485, 0.09549321, 
    0.02364627, 0.1751046, 0.1895007, 0.2592471, 0.2606691,
  0.1552885, 0.07745973, 0.002645311, 0.1118023, 0.1476855, 0.1728353, 
    0.1501231, 0.1122642, 0.1673393, 0.07048532, 0.02753977, -2.717097e-05, 
    0.04840321, 0.09234551, 0.07243846, 0.0314908, 0.1455259, 0.2237607, 
    0.1617672, 0.1452378, 0.1734884, 0.1637156, 0.2093139, 0.0003288474, 
    0.01196196, 0.06427488, 0.1072678, 0.1172924, 0.09585027,
  0.2322633, 0.03048917, 0.005770909, 0.09004479, 0.09450276, 0.06781265, 
    0.08210761, 0.07393093, 0.1003614, 0.03684976, 0.00495824, 7.331586e-05, 
    0.09986189, 0.1725006, 0.04238229, 0.09021363, 0.1311751, 0.0577031, 
    0.1117512, 0.08826678, 0.07141061, 0.08417766, 0.2596352, 0.00346412, 
    0.0653576, 0.1399078, 0.05408464, 0.1750386, 0.1173959,
  0.2566093, 0.0816345, 0.06985474, 0.0784637, 0.04796395, 0.08442161, 
    0.04684659, 0.05168286, 0.05796588, 0.1019171, 0.08938795, 0.07545418, 
    0.1213897, 0.1057531, 0.1065293, 0.1315848, 0.1480474, 0.1155029, 
    0.09320559, 0.1197771, 0.1337739, 0.1547594, 0.1828163, 0.121145, 
    0.07326102, 0.03546299, 0.0978562, 0.1457956, 0.2254114,
  0.05989001, 0.004579332, 0.001919668, 0.01267612, 0.1857372, 0.2254144, 
    0.266494, 0.1326884, 0.06808979, 0.1011912, 0.03830904, 0.08478994, 
    0.05676884, 0.08389207, 0.1025989, 0.0745895, 0.03446738, 0.03245658, 
    0.02660893, 0.02571163, 0.03032826, 0.03257387, 0.02207263, 0.01525719, 
    0.08253101, 0.05333786, 0.04787724, 0.03650177, 0.03243588,
  -4.864526e-07, 2.079518e-08, 3.699834e-09, -0.0003876644, 0.05885946, 
    0.2350326, 0.0585101, 0.1813256, 0.03256349, 0.104514, 0.1328935, 
    0.06299561, 0.04030737, 0.03501652, 0.06694492, 0.0282087, 0.04265174, 
    0.07237214, 0.1059182, 0.09452004, 0.08453036, 0.06043966, 0.1042462, 
    0.05465979, 0.0537817, 0.1592296, 0.1319421, -5.106244e-09, 9.6428e-06,
  9.026786e-09, 1.578331e-09, -3.734673e-09, 0.0003067566, 3.028404e-10, 
    5.020096e-05, -1.508681e-08, 0.0001056584, -5.129039e-06, 0.0970237, 
    0.0797829, 0.1362562, 0.1133724, 0.09470256, 0.0798315, 0.05007557, 
    0.0484181, 0.03178799, 0.1366066, 0.2477382, -0.0001050624, 0.1178549, 
    0.04748222, 0.0279968, 0.05835889, 0.05700947, 0.1380516, 0.01336184, 
    7.65047e-09,
  9.448254e-09, 0.01239527, 0.03999365, 0.01497991, 0.008147152, 
    2.324521e-06, -0.0006491417, 0.01052101, 0.05958607, 0.1544362, 
    0.1763972, 0.1198043, 0.1389372, 0.1632613, 0.1578154, 0.2173948, 
    0.1656818, 0.2591341, 0.2354628, 0.08479849, 0.006857702, 0.1647955, 
    0.07984285, 0.139837, 0.07671754, 0.09340727, 0.2513438, 0.09656062, 
    -4.014483e-05,
  -0.0009548064, 0.03527345, 0.08784228, 0.2338442, 0.05328834, 0.01337076, 
    0.1029772, 0.006030774, 0.001242822, 0.006498527, 0.04629862, 0.06064931, 
    0.1707846, 0.1606851, 0.1534782, 0.1989443, 0.2162048, 0.2048991, 
    0.313174, 0.2020594, 0.08397423, 0.2210112, 0.2241668, 0.1908899, 
    0.2681107, 0.3186797, 0.2282961, 0.2741344, 0.1128357,
  0.2078419, 0.3466441, 0.2363775, 0.2846872, 0.1768067, 0.1651412, 
    0.2072429, 0.1588662, 0.03295429, 0.01811414, 0.003728065, 0.08542981, 
    0.09212581, 0.263394, 0.1632434, 0.2336751, 0.19752, 0.270705, 0.217883, 
    0.2691978, 0.1275149, 0.1023637, 0.1126575, 0.2739826, 0.1094264, 
    0.3587124, 0.3198276, 0.2437449, 0.2515981,
  0.2824051, 0.2861844, 0.2958153, 0.3438185, 0.4696376, 0.2377354, 0.256411, 
    0.2197207, 0.2574989, 0.3412777, 0.2684399, 0.2050296, 0.2343775, 
    0.3011159, 0.6318049, 0.2539604, 0.2235014, 0.283295, 0.3295556, 0.12806, 
    0.1562251, 0.1821756, 0.2762645, 0.3678696, 0.5792692, 0.07926592, 
    0.1606914, 0.2907088, 0.2251252,
  0.1755148, 0.1552034, 0.3078457, 0.3209494, 0.2809316, 0.2369204, 
    0.2803146, 0.4250145, 0.3092918, 0.3433946, 0.3686197, 0.158562, 
    0.2287872, 0.198555, 0.2807941, 0.1281927, 0.1576712, 0.2041211, 
    0.09618928, 0.2332587, 0.1883446, 0.2525012, 0.2710766, 0.1373737, 
    0.2270781, 0.5025458, 0.4878418, 0.2434244, 0.3800316,
  0.1238046, 0.2750675, 0.2950811, 0.2178441, 0.2418126, 0.3227863, 
    0.3477938, 0.4488879, 0.4201984, 0.3880768, 0.3310349, 0.2200053, 
    0.2314216, 0.2978489, 0.2725433, 0.2435998, 0.295682, 0.2721554, 
    0.2396128, 0.1422192, 0.1503315, 0.1922836, 0.1450178, 0.07903948, 
    0.091253, 0.1052285, 0.1913082, 0.1723809, 0.2196898,
  0.4858305, 0.4872543, 0.4886782, 0.490102, 0.4915259, 0.4929497, 0.4943736, 
    0.4887264, 0.4940849, 0.4994433, 0.5048018, 0.5101602, 0.5155187, 
    0.5208771, 0.5269574, 0.5229, 0.5188427, 0.5147853, 0.510728, 0.5066707, 
    0.5026133, 0.4702916, 0.4675666, 0.4648417, 0.4621167, 0.4593918, 
    0.4566668, 0.4539419, 0.4846914,
  0.322566, 0.5097123, 0.4512324, 0.1942824, 0.1266537, 0.1571934, 0.1967883, 
    0.1668871, 0.01885242, 0.07758469, 0.2229841, 0.282537, 0.3222406, 
    0.09758325, 0.2233383, 0.2242044, 0.2607066, 0.2417157, 0.1917982, 
    0.3197546, 0.4820155, 0.4326514, 0.4187864, 0.3239885, 0.399734, 
    0.5026711, 0.3978817, 0.216934, 0.3835669,
  0.1926368, 0.1226104, 0.2728332, 0.100928, 0.1421538, 0.1666638, 0.1687902, 
    0.2754966, 0.394047, 0.3306688, 0.3362791, 0.1350045, 0.2158206, 
    0.2716516, 0.2803495, 0.3776824, 0.389423, 0.3323785, 0.3531193, 
    0.4025574, 0.3866687, 0.3277997, 0.268575, 0.4205985, 0.4637792, 
    0.4062859, 0.4158351, 0.5228019, 0.2575391,
  0.2905194, 0.242593, 0.2470794, 0.3146628, 0.2964609, 0.404317, 0.4457991, 
    0.4371099, 0.4650033, 0.3432729, 0.3017156, 0.3773159, 0.5782961, 
    0.4666923, 0.3972519, 0.4233411, 0.4304108, 0.4804425, 0.5066193, 
    0.4675321, 0.4166486, 0.4087708, 0.455853, 0.3612768, 0.4165194, 
    0.5378612, 0.51335, 0.4782123, 0.366118,
  0.4204619, 0.424123, 0.4028966, 0.3470823, 0.3336397, 0.3713237, 0.3493918, 
    0.370479, 0.3104193, 0.3546162, 0.3623928, 0.2961898, 0.2876598, 
    0.3571037, 0.140581, 0.3455368, 0.3374192, 0.4562207, 0.3403923, 
    0.3337408, 0.2712027, 0.2529508, 0.284303, 0.2038755, 0.02549358, 
    0.22145, 0.3262298, 0.3698167, 0.4203236,
  0.2973155, 0.2581161, 0.1107233, 0.1783826, 0.1932585, 0.2214464, 0.264973, 
    0.2932143, 0.2691754, 0.2336689, 0.1329873, 0.1137195, 0.09064868, 
    0.1553389, 0.1673395, 0.04544939, 0.2025635, 0.1853908, 0.1478769, 
    0.1839062, 0.1286304, 0.1571791, 0.1343593, 0.1261906, 0.02029947, 
    0.1665702, 0.2121594, 0.3075337, 0.247349,
  0.1793923, 0.1235135, 0.0003336077, 0.05964169, 0.1036958, 0.1917306, 
    0.0988043, 0.05970582, 0.09909831, 0.06595849, 0.02711109, 0.0004890042, 
    0.03853456, 0.07177304, 0.03559133, 0.009516057, 0.0841376, 0.2117772, 
    0.1364648, 0.1095662, 0.09361897, 0.09983478, 0.1574429, 0.007796326, 
    0.02360305, 0.02486294, 0.05944696, 0.07284004, 0.09414496,
  0.240034, 0.03384136, 0.001606553, 0.01710637, 0.07575689, 0.04861035, 
    0.05635144, 0.06875139, 0.05904446, 0.02784651, 0.001779541, 
    3.379325e-05, 0.04395651, 0.07550211, 0.03024789, 0.06799824, 0.07809289, 
    0.04413654, 0.08431993, 0.0218815, 0.0229183, 0.03341177, 0.07696028, 
    0.1048842, 0.05364463, 0.1337048, 0.02189813, 0.06292251, 0.09087224,
  0.3163759, 0.121704, 0.04469324, 0.05476739, 0.04604272, 0.02783286, 
    0.03095497, 0.0241269, 0.04326601, 0.1505173, 0.07432714, 0.04144037, 
    0.06336115, 0.0708096, 0.0259518, 0.03679012, 0.04715225, 0.034495, 
    0.02744534, 0.04062752, 0.05252379, 0.07047995, 0.1067496, 0.09738464, 
    0.05555264, 0.01720593, 0.03781159, 0.04083641, 0.08140279,
  0.1222289, 0.002202037, 0.0009835728, 0.01392706, 0.12474, 0.07429026, 
    0.0409111, 0.01501639, 0.04604741, 0.06836476, 0.1114391, 0.1914136, 
    0.04861448, 0.02557686, 0.02803268, 0.07053151, 0.05569333, 0.04467923, 
    0.0473694, 0.05219971, 0.08982404, 0.123902, 0.02436847, 0.004798629, 
    0.04934645, 0.04269435, 0.03283236, 0.05487385, 0.1855128,
  -1.473859e-07, 1.89564e-08, 2.216311e-09, -0.0007084086, 0.05478244, 
    0.04755265, 0.05044533, 0.04591303, 0.03497881, 0.08266873, 0.1197992, 
    0.04373721, 0.02265122, 0.01663224, 0.01706598, 0.01504574, 0.0215322, 
    0.02850071, 0.1019555, 0.06284035, 0.03204577, 0.01490397, 0.2624033, 
    0.08462989, 0.009799768, 0.05090263, 0.1006135, 1.076664e-06, 
    -5.911385e-06,
  4.919981e-09, 1.280614e-09, -1.915425e-09, 0.0003759616, 3.209523e-10, 
    0.001537257, -1.213836e-08, 0.0001151094, -3.65239e-06, 0.1689067, 
    0.09771248, 0.1241723, 0.06551022, 0.06524658, 0.07723709, 0.01008958, 
    0.02081411, 0.01648111, 0.04760285, 0.08347436, 9.215656e-05, 0.1029502, 
    0.02320283, 0.01548033, 0.02594248, 0.04417648, 0.08141826, 0.004762546, 
    7.21401e-09,
  5.789425e-09, 0.01380765, 0.03359989, 0.01028976, 0.007129269, 
    1.403591e-06, -0.0004853112, 0.0071317, 0.04290809, 0.1403393, 0.1820772, 
    0.1088944, 0.1788218, 0.1474094, 0.1424109, 0.203683, 0.1678457, 
    0.1278422, 0.1130414, 0.06331025, 0.005372422, 0.158936, 0.05526317, 
    0.09723105, 0.05826156, 0.06578752, 0.162643, 0.1047, 7.066964e-05,
  6.98647e-05, 0.04428492, 0.05861552, 0.2311088, 0.04996343, 0.009899129, 
    0.0815385, 0.00160268, 0.0005365647, 0.004350144, 0.05206183, 0.05135908, 
    0.1440508, 0.132752, 0.1151741, 0.1558415, 0.2017372, 0.1931855, 
    0.2451373, 0.2147218, 0.06996629, 0.2215736, 0.2078018, 0.1608072, 
    0.2018988, 0.3297583, 0.1905074, 0.2965104, 0.08761342,
  0.2232237, 0.2974094, 0.1762815, 0.202874, 0.1200627, 0.2534439, 0.175779, 
    0.1443757, 0.02006827, 0.01644578, 0.001417922, 0.07692868, 0.119588, 
    0.1892146, 0.1222482, 0.2163022, 0.1693726, 0.2459288, 0.2198282, 
    0.3024689, 0.1175257, 0.09167764, 0.09895783, 0.2295365, 0.09324403, 
    0.2759052, 0.2772578, 0.2965049, 0.276709,
  0.2567648, 0.3013316, 0.3208214, 0.4082962, 0.463175, 0.1795248, 0.2192525, 
    0.199267, 0.2042195, 0.266827, 0.2284639, 0.2311522, 0.2226501, 
    0.2513619, 0.549138, 0.2728468, 0.1885315, 0.2570243, 0.3216813, 
    0.1082598, 0.1457251, 0.1623803, 0.2749664, 0.3584425, 0.4529437, 
    0.04903724, 0.1220815, 0.2613033, 0.2065519,
  0.1258509, 0.109034, 0.2844982, 0.2472072, 0.3324308, 0.2437118, 0.3111013, 
    0.4227859, 0.3012873, 0.3709461, 0.4669992, 0.2134823, 0.2661089, 
    0.2300646, 0.31589, 0.2102272, 0.2056351, 0.2251851, 0.1526949, 
    0.2595136, 0.2499798, 0.305618, 0.2809764, 0.1469509, 0.2103538, 
    0.4585813, 0.4932315, 0.2005793, 0.3999166,
  0.1407248, 0.2160133, 0.3540541, 0.2611252, 0.2766372, 0.369518, 0.3692627, 
    0.4617825, 0.4425671, 0.4284266, 0.4028097, 0.2844851, 0.2804645, 
    0.3605209, 0.3105707, 0.3050103, 0.3257641, 0.3070972, 0.269801, 0.15683, 
    0.1536473, 0.1944638, 0.1499025, 0.07782288, 0.0996564, 0.09993344, 
    0.1537121, 0.1860458, 0.2389702,
  0.4968948, 0.4935788, 0.4902628, 0.4869469, 0.4836309, 0.4803149, 
    0.4769989, 0.4798309, 0.4869626, 0.4940942, 0.5012258, 0.5083574, 
    0.515489, 0.5226207, 0.5417923, 0.5413013, 0.5408103, 0.5403194, 
    0.5398284, 0.5393374, 0.5388464, 0.5155427, 0.512218, 0.5088934, 
    0.5055687, 0.502244, 0.4989194, 0.4955947, 0.4995475,
  0.3785984, 0.5892029, 0.4712025, 0.2176029, 0.1502258, 0.1663073, 
    0.2032041, 0.1901794, 0.03406533, 0.07560285, 0.2592758, 0.2919599, 
    0.3651069, 0.06709781, 0.2121049, 0.2888246, 0.3002139, 0.2175342, 
    0.1967803, 0.2730948, 0.5172323, 0.4493547, 0.4019045, 0.2740054, 
    0.4322627, 0.507843, 0.273255, 0.1281559, 0.3825802,
  0.1577945, 0.08987202, 0.2523509, 0.06963033, 0.1028533, 0.1476896, 
    0.1101742, 0.2438809, 0.3540009, 0.3173204, 0.3174205, 0.1260133, 
    0.1910309, 0.1863839, 0.2475974, 0.3270054, 0.3645464, 0.283765, 
    0.3162092, 0.3656494, 0.3570391, 0.3132622, 0.2617296, 0.4074659, 
    0.4524807, 0.4491981, 0.4029454, 0.4568329, 0.1785177,
  0.2662641, 0.212771, 0.2015279, 0.2973896, 0.2482429, 0.3684551, 0.3959097, 
    0.3689914, 0.418639, 0.3212774, 0.250562, 0.3711924, 0.5618739, 
    0.4461763, 0.396331, 0.3962249, 0.4362538, 0.4926074, 0.4883666, 
    0.4544213, 0.3950923, 0.4175832, 0.4436282, 0.3286896, 0.4328067, 
    0.5316672, 0.5041586, 0.4648088, 0.3273208,
  0.4397013, 0.4534365, 0.3662912, 0.3381978, 0.3480852, 0.3663568, 
    0.3826489, 0.3930022, 0.335898, 0.3617536, 0.3073453, 0.2477897, 
    0.2325702, 0.3837041, 0.1613714, 0.3009135, 0.2865781, 0.3941421, 
    0.3300323, 0.3180084, 0.2789284, 0.2305663, 0.2567095, 0.1959014, 
    0.02831883, 0.2224687, 0.3347688, 0.3663326, 0.4055457,
  0.2611337, 0.2193396, 0.06283575, 0.1235001, 0.1666707, 0.2001363, 
    0.2383654, 0.2075453, 0.2208928, 0.1350324, 0.08324175, 0.07363427, 
    0.04263924, 0.1687182, 0.1628498, 0.02635162, 0.1791607, 0.136043, 
    0.1464732, 0.1490913, 0.09529687, 0.1362522, 0.1085785, 0.1383757, 
    0.02894551, 0.111108, 0.1904355, 0.1832254, 0.2656685,
  0.1480311, 0.06828389, -0.0005469943, 0.01206027, 0.0896304, 0.2211791, 
    0.06880985, 0.0267379, 0.02899583, 0.03889971, 0.02516019, 0.0008840084, 
    0.03519128, 0.05352167, 0.03256182, 0.00235393, 0.04384822, 0.1921639, 
    0.1089008, 0.05820448, 0.04875619, 0.07309262, 0.06792542, 0.05075066, 
    0.02124041, 0.01113914, 0.01734111, 0.01792633, 0.040345,
  0.1365001, 0.04074243, 0.0001049899, 0.003075973, 0.04411408, 0.01943593, 
    0.02597281, 0.03919151, 0.02894983, 0.004029533, 0.0007134598, 
    1.88327e-05, 0.0106262, 0.02710712, 0.01073659, 0.03805933, 0.03577369, 
    0.01382892, 0.03220134, 0.008539748, 0.01188097, 0.006442317, 0.01850687, 
    0.1223557, 0.0439706, 0.1279186, 0.003822126, 0.01911948, 0.03537561,
  0.09260576, 0.08829913, 0.03524779, 0.04000564, 0.006858937, 0.006530944, 
    0.0147342, 0.004723529, 0.02175775, 0.02230082, 0.03444498, 0.01870696, 
    0.0151497, 0.01197308, 0.006058617, 0.01600952, 0.02329567, 0.01121145, 
    0.006577742, 0.007543413, 0.009948358, 0.01386871, 0.01801755, 
    0.08513746, 0.04877242, 0.01248731, 0.001719328, 0.01246382, 0.02792405,
  0.01360375, 0.002431628, 0.0006329332, 0.01840129, 0.02482093, 0.01792005, 
    0.01014286, 0.002770307, 0.04866123, 0.04882835, 0.01950578, 0.03197301, 
    0.01614394, 0.007884596, 0.005303665, 0.02566638, 0.03413941, 0.02496824, 
    0.02542408, 0.09165987, 0.09212168, 0.1567028, 0.07959682, 0.002074082, 
    0.02946314, 0.0115329, 0.00388056, 0.004770223, 0.02401781,
  -3.796297e-08, 1.809886e-08, 1.756432e-09, -0.0007053768, 0.03046337, 
    0.01365454, 0.009358878, 0.01596933, 0.005060419, 0.01790447, 0.08161293, 
    0.01322349, 0.006727084, 0.003078166, 0.00324233, 0.006286175, 
    0.008042244, 0.008095412, 0.05201313, 0.03384233, 0.01037577, 
    0.002201948, 0.2663624, 0.09637383, 0.001106977, 0.01647326, 0.04760318, 
    -1.212664e-05, -1.424818e-05,
  3.548643e-09, 1.096563e-09, -1.023256e-09, 7.591923e-05, 2.701961e-10, 
    0.0001289648, 6.386904e-09, -1.15797e-05, -1.937777e-05, 0.3289783, 
    0.05631511, 0.04687496, 0.01818123, 0.02591481, 0.01626747, 0.001028812, 
    0.009886246, 0.02261577, 0.02403898, 0.07009763, -4.271633e-06, 
    0.08453725, 0.004947219, 0.007515463, 0.01012737, 0.02695453, 0.03389375, 
    0.001017526, 6.902011e-09,
  4.656832e-09, 0.008496506, 0.02189127, 0.01463378, 0.007997207, 
    1.025032e-06, -0.0003711959, 0.005169764, 0.02780992, 0.1198794, 
    0.1807733, 0.110419, 0.1744135, 0.1311534, 0.1546729, 0.1483225, 
    0.1343896, 0.08835942, 0.04461646, 0.04449276, 0.005264616, 0.1527172, 
    0.04071368, 0.08577141, 0.04188688, 0.03782196, 0.1336634, 0.04511934, 
    0.0001439474,
  0.0006615483, 0.01593428, 0.03841417, 0.2369039, 0.02749071, 0.005440573, 
    0.06810801, 0.000588286, 0.0001500748, 0.002716178, 0.05845543, 
    0.04222498, 0.1170058, 0.1133763, 0.09778979, 0.1147936, 0.1679783, 
    0.1733977, 0.1860759, 0.2053519, 0.060194, 0.2208116, 0.1932262, 
    0.1362948, 0.1483004, 0.3137715, 0.1916224, 0.2204828, 0.08319064,
  0.1610051, 0.2292566, 0.132321, 0.1453141, 0.2533475, 0.3205113, 0.1366982, 
    0.1307314, 0.01351949, 0.007876215, 0.0004770039, 0.06982008, 0.1215931, 
    0.1487432, 0.1000505, 0.1805532, 0.1494017, 0.2285318, 0.1755223, 
    0.3238958, 0.099833, 0.08292176, 0.08816025, 0.2104991, 0.06733163, 
    0.2501977, 0.2539441, 0.2694685, 0.2346337,
  0.1954804, 0.2988316, 0.3419903, 0.4830808, 0.4771444, 0.14062, 0.184409, 
    0.1516802, 0.1589909, 0.2137898, 0.1729016, 0.2236941, 0.2061673, 
    0.1860202, 0.4326534, 0.2704567, 0.1639459, 0.2289523, 0.260306, 
    0.1115967, 0.1412049, 0.1279827, 0.2887869, 0.2748719, 0.3707325, 
    0.03345368, 0.1012467, 0.2184081, 0.1757901,
  0.1036882, 0.08568161, 0.2325072, 0.1848172, 0.3800176, 0.2538747, 
    0.3217725, 0.4031657, 0.3224291, 0.3905566, 0.5641294, 0.2801595, 
    0.3366121, 0.2467792, 0.3406065, 0.2911109, 0.2809676, 0.2240402, 
    0.1871466, 0.3152657, 0.2780751, 0.3528307, 0.3099047, 0.1628138, 
    0.1933263, 0.4103829, 0.5042, 0.1716374, 0.3045594,
  0.1192909, 0.2191327, 0.419813, 0.3633708, 0.3548541, 0.454122, 0.4153258, 
    0.4984137, 0.441805, 0.4319436, 0.4497145, 0.3644043, 0.3761816, 
    0.4191172, 0.4201594, 0.3630354, 0.3661747, 0.3321677, 0.2828858, 
    0.1820868, 0.1713279, 0.1977475, 0.167468, 0.07981639, 0.1121245, 
    0.1149158, 0.1396997, 0.1994478, 0.2580298,
  0.3602235, 0.3580395, 0.3558554, 0.3536714, 0.3514873, 0.3493033, 
    0.3471192, 0.3860084, 0.395802, 0.4055955, 0.415389, 0.4251826, 
    0.4349761, 0.4447696, 0.4355595, 0.4369621, 0.4383648, 0.4397675, 
    0.4411701, 0.4425728, 0.4439754, 0.4888912, 0.4798791, 0.470867, 
    0.4618548, 0.4528427, 0.4438306, 0.4348184, 0.3619708,
  0.4308827, 0.5595596, 0.4760357, 0.2272805, 0.1453083, 0.1167936, 0.141626, 
    0.174095, 0.02795917, 0.04337525, 0.1910334, 0.3119688, 0.4079672, 
    0.04143358, 0.2573038, 0.345846, 0.3779869, 0.2167339, 0.1544049, 
    0.2374199, 0.4844382, 0.4769331, 0.3705147, 0.2106982, 0.4315033, 
    0.5382953, 0.1753055, 0.05522206, 0.3569557,
  0.1164833, 0.05706066, 0.1823202, 0.04070281, 0.06875546, 0.1244096, 
    0.06799381, 0.1765078, 0.3129284, 0.2910112, 0.2686969, 0.1262304, 
    0.1722195, 0.13041, 0.2214503, 0.275222, 0.3296518, 0.2344558, 0.2738117, 
    0.3236484, 0.306108, 0.3014674, 0.2635361, 0.4218553, 0.4143698, 
    0.5057677, 0.3792304, 0.3778545, 0.1524006,
  0.2293346, 0.1926045, 0.1713317, 0.2470397, 0.1959349, 0.2884699, 0.342512, 
    0.3141534, 0.3518686, 0.2927506, 0.2050685, 0.3392324, 0.5226296, 
    0.3991969, 0.3463455, 0.3553631, 0.4102345, 0.4735963, 0.4421228, 
    0.3875039, 0.3584488, 0.3875943, 0.370177, 0.3082627, 0.4338036, 
    0.5695361, 0.5098688, 0.4392465, 0.2964841,
  0.4015081, 0.4257274, 0.3321433, 0.3068234, 0.3348759, 0.3293803, 
    0.3900673, 0.3702442, 0.3059862, 0.3238314, 0.234618, 0.1783156, 
    0.2308799, 0.3425691, 0.1862695, 0.244395, 0.217129, 0.3344221, 
    0.3142841, 0.3094232, 0.2652959, 0.2028183, 0.2149981, 0.1648618, 
    0.03086403, 0.2147413, 0.3548853, 0.3539831, 0.3930161,
  0.1896013, 0.1514841, 0.03049617, 0.07978913, 0.146074, 0.1827256, 
    0.1945712, 0.1252949, 0.1507681, 0.07981692, 0.05932355, 0.0368668, 
    0.02208815, 0.1841513, 0.1638297, 0.02173897, 0.1550909, 0.127024, 
    0.1136643, 0.1152805, 0.08261128, 0.102009, 0.08471552, 0.1423371, 
    0.02564487, 0.06742171, 0.111459, 0.1224017, 0.2122373,
  0.03771968, 0.02318056, -4.964974e-06, 0.003563634, 0.06709352, 0.1824735, 
    0.04502215, 0.01353131, 0.01166787, 0.01543075, 0.01785111, 0.0009173363, 
    0.02972856, 0.04610698, 0.03511039, 0.0005288573, 0.02221829, 0.1591815, 
    0.06436955, 0.02671921, 0.01866137, 0.03703627, 0.02763517, 0.04773249, 
    0.01301628, 0.007075432, 0.007645999, 0.004913582, 0.006780635,
  0.0489955, 0.06200501, -4.955644e-05, 0.0009634635, 0.02041693, 
    0.002164317, 0.01028252, 0.01610462, 0.01202223, 0.001225034, 
    0.0001706742, 1.394466e-05, 0.002751756, 0.009479471, 0.002852844, 
    0.0197542, 0.01186825, 0.001826128, 0.014177, 0.003072399, 0.00450794, 
    0.002308054, 0.006862403, 0.04049185, 0.03602385, 0.1084571, 0.001788243, 
    0.008509467, 0.01302468,
  0.034657, 0.03222366, 0.02956055, 0.0260748, 0.0005685549, 0.001111735, 
    0.00836921, 0.000555362, 0.01013877, 0.006261729, 0.02178058, 0.00652418, 
    0.002483143, 0.002538095, 0.001199908, 0.008401793, 0.01152398, 
    0.00288708, 0.001355015, 0.002761777, 0.003476713, 0.003489101, 
    0.005732429, 0.08080806, 0.04404895, 0.00994577, -0.0007384836, 
    0.004700098, 0.008841435,
  0.003542926, 0.001462647, 0.0004436042, 0.009968208, 0.008164799, 
    0.006135287, 0.003563812, 0.001018703, 0.05663242, 0.03919529, 
    0.007809547, 0.007991095, 0.005419658, 0.001102618, 0.001106699, 
    0.006317772, 0.008530623, 0.002621438, 0.004604596, 0.01567376, 
    0.0173671, 0.04487403, 0.08472712, 0.001514583, 0.02251543, 0.001593194, 
    0.0002163238, 0.0003265697, 0.004785759,
  -3.16755e-08, 1.775507e-08, 1.594324e-09, -0.0004605264, 0.01365082, 
    0.006364554, 0.001563098, 0.007526319, 0.000944318, 0.007411702, 
    0.03928459, 0.001432779, 0.002590992, 0.0005314809, 0.0009448823, 
    0.0002905327, 0.002217368, 0.001428429, 0.02210435, 0.01456293, 
    0.002395042, 0.0008210311, 0.1864499, 0.08871163, 0.0004596045, 
    0.006365378, 0.01971478, 4.043608e-06, -1.751567e-05,
  3.035436e-09, 9.211968e-10, -5.190524e-10, -1.088678e-06, 2.714455e-10, 
    8.645612e-06, 1.107767e-08, -1.32072e-06, -6.489724e-05, 0.2329402, 
    0.01621044, 0.01545617, 0.006112494, 0.01238619, 0.004152223, 
    0.0004280257, 0.01132701, 0.007784734, 0.01140042, 0.0496633, 
    -1.754275e-06, 0.0646602, 0.001219361, 0.001805085, 0.002934039, 
    0.0103589, 0.01566977, 0.0004092651, 6.518068e-09,
  4.216758e-09, 0.002250496, 0.01300766, 0.01105102, 0.00704838, 
    8.852091e-07, -0.0003142696, 0.005557576, 0.01986115, 0.1017196, 
    0.1824162, 0.1044372, 0.1385765, 0.08980469, 0.1282276, 0.09260669, 
    0.1023633, 0.0644491, 0.02351915, 0.05365189, 0.003601787, 0.1286029, 
    0.03367005, 0.07787807, 0.0281635, 0.01945404, 0.05112128, 0.01873188, 
    -5.847615e-05,
  0.0005990643, 0.004701353, 0.02421004, 0.2281072, 0.01347336, 0.00291309, 
    0.05635066, 0.0003684178, 1.718222e-05, 0.00176578, 0.06380732, 
    0.0325483, 0.09619827, 0.09613337, 0.07712303, 0.08928458, 0.1305378, 
    0.1434566, 0.1430911, 0.183179, 0.05275558, 0.18401, 0.1703115, 
    0.1225166, 0.1072759, 0.2462432, 0.1552481, 0.1441559, 0.05028263,
  0.08996295, 0.1660151, 0.1064614, 0.123658, 0.2419185, 0.2679743, 
    0.1004449, 0.1123012, 0.007860827, 0.003249662, 0.0001303751, 0.06162428, 
    0.1875098, 0.1205929, 0.08283173, 0.1476394, 0.1369547, 0.1930342, 
    0.1444968, 0.288729, 0.08495961, 0.06822922, 0.07886999, 0.1990191, 
    0.05304281, 0.2260952, 0.2434001, 0.1947298, 0.1902718,
  0.1503646, 0.3174372, 0.346392, 0.5017528, 0.4443526, 0.09675944, 
    0.1425347, 0.1149069, 0.1228477, 0.1748239, 0.1331344, 0.2158051, 
    0.2004337, 0.1287034, 0.363856, 0.2999186, 0.1418654, 0.2014043, 
    0.1944973, 0.121718, 0.1287087, 0.1032193, 0.3450823, 0.2230726, 
    0.3215654, 0.02177369, 0.08832166, 0.1715392, 0.1453348,
  0.09002253, 0.07089563, 0.1737057, 0.1414464, 0.4396209, 0.2711978, 
    0.3558272, 0.3569472, 0.3792504, 0.3699341, 0.5687133, 0.2855509, 
    0.3919441, 0.2877815, 0.3741274, 0.3476872, 0.339038, 0.2231814, 
    0.2236762, 0.3434295, 0.3081091, 0.4089237, 0.3585092, 0.194562, 
    0.1775211, 0.3352115, 0.5001333, 0.1498602, 0.2257764,
  0.2042124, 0.253839, 0.485517, 0.382045, 0.4086333, 0.5745741, 0.4898987, 
    0.4966834, 0.4805946, 0.4680854, 0.4820672, 0.4112906, 0.4033192, 
    0.4516797, 0.4741575, 0.4291503, 0.3938181, 0.3487567, 0.3051309, 
    0.2480851, 0.2141644, 0.2093173, 0.1863264, 0.1202111, 0.1250146, 
    0.1128235, 0.1352044, 0.2205955, 0.3121615,
  0.2271547, 0.227679, 0.2282032, 0.2287275, 0.2292517, 0.229776, 0.2303003, 
    0.2631919, 0.2782507, 0.2933095, 0.3083682, 0.323427, 0.3384857, 
    0.3535445, 0.3920082, 0.3888677, 0.3857271, 0.3825866, 0.379446, 
    0.3763055, 0.373165, 0.3517806, 0.3393381, 0.3268956, 0.3144532, 
    0.3020107, 0.2895682, 0.2771257, 0.2267353,
  0.4199008, 0.4808587, 0.3178482, 0.1573866, 0.153267, 0.07681764, 
    0.09912172, 0.1533397, 0.01427033, 0.004599411, 0.08611097, 0.2347335, 
    0.4020317, 0.0145449, 0.3657908, 0.3970742, 0.5132601, 0.278322, 
    0.1349567, 0.2196104, 0.4378113, 0.4940748, 0.3203818, 0.1627652, 
    0.430629, 0.5721841, 0.1140873, 0.01754793, 0.2858803,
  0.08820839, 0.03843893, 0.1175191, 0.02571342, 0.05136772, 0.09966121, 
    0.04834467, 0.1151648, 0.2701845, 0.2379223, 0.2164339, 0.1200271, 
    0.1509627, 0.09675509, 0.1891676, 0.2106541, 0.2579129, 0.1722553, 
    0.2213697, 0.2532034, 0.2471485, 0.2798174, 0.2577228, 0.3990098, 
    0.3710728, 0.4768938, 0.325744, 0.2728528, 0.1173835,
  0.1853171, 0.1722277, 0.1391565, 0.1836742, 0.1421375, 0.2235651, 
    0.2773743, 0.2432832, 0.2752926, 0.2466922, 0.1755682, 0.2944469, 
    0.4560544, 0.3139549, 0.2684519, 0.2905765, 0.3467265, 0.425292, 
    0.3931549, 0.3311816, 0.298138, 0.3245087, 0.2900028, 0.2332411, 
    0.393907, 0.5556238, 0.4643958, 0.4125792, 0.2672304,
  0.3368302, 0.3486791, 0.2880734, 0.2579486, 0.290872, 0.2789261, 0.3572217, 
    0.3094581, 0.24891, 0.2485015, 0.1639876, 0.1216948, 0.1918611, 0.284046, 
    0.2160879, 0.1765911, 0.1561804, 0.2522893, 0.2782031, 0.2811385, 
    0.2314996, 0.1557657, 0.182777, 0.1317269, 0.03228928, 0.2215241, 
    0.3439187, 0.3112703, 0.3617565,
  0.1520375, 0.1123402, 0.01927287, 0.05074598, 0.1188976, 0.1468907, 
    0.181124, 0.09336183, 0.1006201, 0.04635352, 0.04027503, 0.0178376, 
    0.01381122, 0.1456272, 0.1558775, 0.02046839, 0.1279911, 0.1198095, 
    0.08108894, 0.08817806, 0.06932403, 0.07878911, 0.06094776, 0.1355642, 
    0.01190991, 0.04927025, 0.05665844, 0.08489871, 0.1557387,
  0.01660017, 0.01036356, 0.0005418501, 0.001862179, 0.02170685, 0.1170665, 
    0.0135086, 0.005398788, 0.006406195, 0.00712625, 0.006942603, 
    0.0003719561, 0.0206767, 0.02693156, 0.033845, 0.0002662693, 0.01267207, 
    0.1253218, 0.02909558, 0.01126229, 0.009760071, 0.01439132, 0.01234056, 
    0.02606193, 0.009103729, 0.003857568, 0.002930448, 0.002257087, 
    0.001829349,
  0.02329807, 0.06682921, -2.114807e-05, 0.0005253759, 0.006678691, 
    0.000571931, 0.001980651, 0.00344312, 0.008838241, 0.0006661465, 
    7.410323e-05, 6.932889e-06, 0.001262976, 0.003849221, 0.001005401, 
    0.008837054, 0.003769462, 0.0003545678, 0.005719405, 0.001088022, 
    0.001381391, 0.001116539, 0.003589761, 0.02013889, 0.02852344, 
    0.08542372, 0.0007454344, 0.00364568, 0.005635082,
  0.01794437, 0.01468849, 0.02719043, 0.01942798, 0.0001130873, 0.0004560383, 
    0.00459008, 0.0001305639, 0.004454678, 0.003543752, 0.01450286, 
    0.002653638, 0.0002489503, 0.001206372, 0.0004901395, 0.005091696, 
    0.00472606, 0.001104579, 0.000567262, 0.001516167, 0.001778681, 
    0.001637721, 0.00294641, 0.08312272, 0.04408122, 0.006595016, 
    -0.0001276946, 0.002400051, 0.004573082,
  0.001709548, 0.001175136, 0.000287298, 0.006266539, 0.003980852, 
    0.003364848, 0.001937605, 0.0005460602, 0.04735901, 0.04531003, 
    0.002653931, 0.003441894, 0.003408724, 0.0004283899, 0.0005191888, 
    0.001757668, 0.002041045, 0.0004149036, 0.0007506717, 0.003763888, 
    0.00348158, 0.0142666, 0.02384296, 0.001968439, 0.01976455, 0.0004260234, 
    6.221253e-05, 0.0001022743, 0.002290769,
  2.2106e-10, 1.746776e-08, 1.528463e-09, -9.634224e-05, 0.008539767, 
    0.003791018, 0.0003932253, 0.003895455, 0.0003042689, 0.002543018, 
    0.0172022, -4.973786e-06, 0.0003992909, 0.0001149517, 0.0004418081, 
    -4.903702e-05, 0.0006500212, 0.0004910947, 0.01045242, 0.007928331, 
    0.000898206, 0.0004894703, 0.1110322, 0.07734389, 0.0002683657, 
    0.0035187, 0.009818912, -1.372294e-07, -8.126012e-05,
  2.802079e-09, 8.289e-10, -2.062437e-10, -5.056356e-08, 2.516286e-10, 
    3.81086e-06, 9.315828e-09, 7.997817e-08, -9.357117e-05, 0.1053039, 
    0.006501078, 0.005886425, 0.003461609, 0.005505184, 0.001980401, 
    0.0002499886, 0.005728292, 0.00281348, 0.005113395, 0.03032177, 
    -1.000266e-06, 0.05172715, 0.0006423062, 4.53282e-05, 0.001497164, 
    0.004852027, 0.009066, 0.0002206427, 6.441953e-09,
  4.090994e-09, 0.0008511515, 0.008036712, 0.006101916, 0.007185395, 
    8.144161e-07, -0.0002877254, 0.01073758, 0.014615, 0.07365908, 0.1640814, 
    0.08047163, 0.08896552, 0.05721082, 0.081235, 0.07456642, 0.07988714, 
    0.04625107, 0.01533894, 0.04251811, 0.002835108, 0.09755519, 0.02600673, 
    0.05970311, 0.01802579, 0.008344318, 0.02528634, 0.01060392, -0.0001056518,
  0.0003081242, 0.001969856, 0.01550326, 0.2078971, 0.008325529, 0.001841827, 
    0.04417046, 0.0001588205, -5.417021e-06, 0.0009003917, 0.07570328, 
    0.02130334, 0.07991965, 0.07238927, 0.05808597, 0.06950166, 0.09156669, 
    0.1040862, 0.1003394, 0.1613783, 0.04304593, 0.1395703, 0.1427962, 
    0.1089451, 0.07731818, 0.1754653, 0.0950585, 0.08670736, 0.02321116,
  0.05165685, 0.118047, 0.07378325, 0.1076099, 0.1780788, 0.1837313, 
    0.07381994, 0.09156317, 0.009443833, 0.001748152, 6.8151e-05, 0.05600367, 
    0.2246427, 0.09011176, 0.06906842, 0.1244215, 0.1165709, 0.1514748, 
    0.1044371, 0.2440405, 0.06883941, 0.05821486, 0.07141331, 0.187474, 
    0.04742928, 0.2043669, 0.1998342, 0.1490801, 0.1511494,
  0.122108, 0.3120869, 0.3309102, 0.4476887, 0.3764382, 0.07116516, 
    0.0972708, 0.08865118, 0.09096057, 0.1371408, 0.1041014, 0.2099171, 
    0.2240172, 0.1103262, 0.2967623, 0.2284583, 0.1511204, 0.1718759, 
    0.1395155, 0.1213698, 0.1159477, 0.0750527, 0.3104174, 0.2201287, 
    0.2901166, 0.01487301, 0.07351439, 0.1235861, 0.110471,
  0.07933525, 0.05485157, 0.1471033, 0.1091275, 0.3646197, 0.3034872, 
    0.3582936, 0.3171279, 0.3660229, 0.3352702, 0.5820109, 0.28006, 
    0.4051146, 0.2876933, 0.3437314, 0.365398, 0.36421, 0.2064736, 0.2788165, 
    0.3313366, 0.3397938, 0.4219412, 0.3842219, 0.2286917, 0.1964295, 
    0.2700113, 0.5065317, 0.1360085, 0.1826513,
  0.3930906, 0.2676068, 0.5300423, 0.4534225, 0.5133716, 0.6840414, 
    0.5115978, 0.458934, 0.5375394, 0.515882, 0.5083129, 0.4827177, 
    0.4246172, 0.4452451, 0.5125213, 0.5211061, 0.4159778, 0.3718632, 
    0.348235, 0.2871725, 0.2760945, 0.2081463, 0.2253323, 0.1624712, 
    0.1119327, 0.09656396, 0.1319999, 0.1966037, 0.4167355,
  0.07568359, 0.07368695, 0.07169032, 0.06969368, 0.06769705, 0.06570041, 
    0.06370378, 0.09061539, 0.1115911, 0.1325669, 0.1535426, 0.1745184, 
    0.1954941, 0.2164699, 0.3041536, 0.3023537, 0.3005538, 0.2987539, 
    0.296954, 0.2951542, 0.2933543, 0.2399513, 0.2227721, 0.2055928, 
    0.1884136, 0.1712344, 0.1540551, 0.1368759, 0.07728089,
  0.395285, 0.4188643, 0.1423357, 0.01724516, 0.09788232, 0.05513539, 
    0.06849866, 0.03001795, -0.0001458917, 0.000375685, 0.05955901, 
    0.1408713, 0.316228, 0.004852881, 0.4352686, 0.4449829, 0.5488642, 
    0.2782513, 0.1222829, 0.2309694, 0.4069593, 0.5378768, 0.2552741, 
    0.1177617, 0.4322754, 0.5842563, 0.1065663, 0.005044947, 0.2022827,
  0.07162957, 0.02889536, 0.07662498, 0.01821407, 0.03793856, 0.06950173, 
    0.03465097, 0.08069751, 0.2251195, 0.1749759, 0.1573669, 0.1113787, 
    0.1235477, 0.07638258, 0.146035, 0.1554859, 0.1853765, 0.1239295, 
    0.169734, 0.1933719, 0.1834577, 0.2536971, 0.2379247, 0.3601816, 
    0.3202071, 0.3737021, 0.2395188, 0.1731629, 0.08989272,
  0.1291378, 0.1332786, 0.1008385, 0.1276983, 0.1012692, 0.1747275, 0.215778, 
    0.1839428, 0.2113243, 0.1985738, 0.1464256, 0.23647, 0.3682982, 
    0.2386557, 0.1875116, 0.2121807, 0.2708896, 0.3616428, 0.3412673, 
    0.2836818, 0.229162, 0.2444233, 0.2052118, 0.1509838, 0.3252492, 
    0.4786659, 0.3858626, 0.3362758, 0.2055332,
  0.2613674, 0.2778386, 0.2280525, 0.1997022, 0.2408045, 0.2309953, 0.30124, 
    0.2447632, 0.1931437, 0.1806845, 0.1038426, 0.07522962, 0.1494511, 
    0.224052, 0.1963948, 0.1237735, 0.1067571, 0.175562, 0.2206655, 0.224095, 
    0.1743832, 0.1010812, 0.1218817, 0.105844, 0.03247142, 0.1940464, 
    0.2866207, 0.258235, 0.3021771,
  0.123475, 0.07411835, 0.01362245, 0.03165828, 0.08411052, 0.1141238, 
    0.1327555, 0.0560981, 0.06665795, 0.02747788, 0.02487301, 0.009444105, 
    0.008443883, 0.09371491, 0.1373529, 0.01405543, 0.08218405, 0.07875012, 
    0.0525754, 0.05773934, 0.04317363, 0.05986688, 0.03983756, 0.1204439, 
    0.005166294, 0.03301035, 0.03227401, 0.05561621, 0.1161816,
  0.01037624, 0.006424628, 0.0003973856, 0.001207202, 0.00668593, 0.05898185, 
    0.004364241, 0.002229551, 0.004149017, 0.004040774, 0.002953338, 
    0.0001437467, 0.01700151, 0.00975339, 0.02601988, 0.0001759423, 
    0.007721104, 0.0914858, 0.01272268, 0.005249171, 0.004760034, 
    0.005280626, 0.007015863, 0.01653999, 0.006576327, 0.001676171, 
    0.001701517, 0.001280116, 0.0009766145,
  0.01453347, 0.05458402, 5.812748e-06, 0.0003473885, -0.0008419774, 
    0.0003707972, 0.000787566, 0.001369957, 0.002916856, 0.0004364517, 
    4.810788e-05, 2.435195e-06, 0.0007699652, 0.001928601, 0.0002661606, 
    0.003253781, 0.001413825, 0.0001739171, 0.001578711, 0.0003683985, 
    0.0004664761, 0.0006924809, 0.002242892, 0.0128497, 0.02001411, 
    0.06904181, 0.0003352613, 0.002092664, 0.003251656,
  0.01150553, 0.007635194, 0.02658834, 0.02566436, 6.681785e-05, 
    0.0003039486, 0.001951034, 6.476489e-05, 0.001814238, 0.002374341, 
    0.007173833, 0.0009811177, -5.437305e-05, 0.0007811278, 0.0002899998, 
    0.002565237, 0.001747995, 0.0005613926, 0.0003659198, 0.0009863677, 
    0.001106857, 0.001103068, 0.00189401, 0.07048456, 0.03946964, 
    0.004826806, 0.0001126268, 0.001552574, 0.002937117,
  0.001041244, 0.0007863431, 0.0001422862, 0.004901229, 0.002531653, 
    0.002208013, 0.00130469, 0.000346946, 0.03594508, 0.05700268, 
    0.001083786, 0.001992873, 0.001335816, 0.0002618802, 0.0003245734, 
    0.0006779497, 0.0009418977, 0.0002092904, 0.0003911721, 0.002000944, 
    0.001623736, 0.006590165, 0.005618322, 0.002443433, 0.01503574, 
    0.0001584734, 3.217063e-05, 5.610742e-05, 0.00142218,
  2.26729e-09, 1.733416e-08, 1.520891e-09, -7.679781e-05, 0.007255327, 
    0.002601417, 0.0001476711, 0.001935228, 0.0001412296, 0.001395409, 
    0.007538347, 2.224045e-05, 0.0001261477, 5.22197e-05, 0.0002831533, 
    -2.448917e-05, 0.000242278, 0.0002709381, 0.004911928, 0.003918596, 
    0.0003837442, 0.0003383283, 0.07742725, 0.06326693, 0.0001780574, 
    0.002303836, 0.006043922, -5.431914e-08, -0.0002021135,
  2.716458e-09, 7.916447e-10, -1.309861e-10, -1.412296e-06, 2.335549e-10, 
    1.622869e-05, 7.789585e-09, 1.199885e-07, -7.041177e-05, 0.04601797, 
    0.003761878, 0.002983916, 0.002821094, 0.002749431, 0.001283896, 
    0.00017069, 0.001619129, 0.001358849, 0.002584319, 0.01314232, 
    -6.698497e-07, 0.04171776, 0.0004128717, -0.0004824103, 0.0009354295, 
    0.002416951, 0.006147052, 0.0001418353, 6.115159e-09,
  4.092497e-09, 0.0002639517, 0.004890536, 0.00403141, 0.006276883, 
    7.613705e-07, -0.0002559636, 0.02353331, 0.01243501, 0.05357153, 
    0.1390598, 0.05319072, 0.04943588, 0.03360073, 0.05213533, 0.04353992, 
    0.05738686, 0.03342176, 0.01018425, 0.02985169, 0.001342573, 0.069779, 
    0.01665549, 0.0383834, 0.01000039, 0.003535299, 0.01574312, 0.006872726, 
    -9.337905e-05,
  3.933597e-05, 0.00118537, 0.01067298, 0.189539, 0.004894524, 0.001374001, 
    0.03531343, 8.835673e-05, -1.436786e-05, 0.0005375909, 0.07214658, 
    0.01354715, 0.06216512, 0.05382014, 0.04121808, 0.04984963, 0.06106136, 
    0.06907662, 0.06162287, 0.1398189, 0.03589878, 0.104917, 0.1147692, 
    0.09513786, 0.05640165, 0.1080525, 0.05263149, 0.04559978, 0.01481755,
  0.03028712, 0.08425099, 0.04854242, 0.08933239, 0.1353458, 0.1544753, 
    0.05396265, 0.07977595, 0.01706823, 0.001107711, 3.475379e-05, 
    0.05005365, 0.2180368, 0.07457379, 0.056157, 0.1007737, 0.09403972, 
    0.1163647, 0.0633646, 0.2162038, 0.053573, 0.05295511, 0.062994, 
    0.1654905, 0.04068721, 0.1856865, 0.1409103, 0.1090581, 0.1122099,
  0.08402808, 0.2921593, 0.2993528, 0.3920393, 0.3004535, 0.04907025, 
    0.07434185, 0.07254213, 0.06736083, 0.1083857, 0.08146577, 0.2197592, 
    0.243195, 0.0992528, 0.2463264, 0.1658291, 0.1708966, 0.146119, 
    0.1196565, 0.1076409, 0.1044946, 0.06373701, 0.242754, 0.1975987, 
    0.2698991, 0.01165545, 0.05418332, 0.08722249, 0.07470779,
  0.06397562, 0.03832239, 0.1367819, 0.07883705, 0.3329783, 0.264734, 
    0.356336, 0.3105565, 0.3414042, 0.3412359, 0.5550362, 0.2845303, 
    0.4243541, 0.296256, 0.2991718, 0.3391848, 0.3748927, 0.1950064, 
    0.3184583, 0.2926152, 0.3125523, 0.4158083, 0.4137203, 0.2652044, 
    0.2150821, 0.2167096, 0.5089168, 0.131814, 0.1500029,
  0.4264787, 0.3020801, 0.5421416, 0.5067453, 0.5471228, 0.6308046, 
    0.5125386, 0.4258057, 0.5079234, 0.4789225, 0.5052299, 0.4597379, 
    0.4380805, 0.4302081, 0.4784352, 0.4798865, 0.3603257, 0.3147005, 
    0.3365154, 0.3039327, 0.2633034, 0.2000139, 0.2411495, 0.2368819, 
    0.09642004, 0.08137226, 0.124938, 0.1835074, 0.3865738,
  0.04348774, 0.04363547, 0.04378319, 0.04393091, 0.04407863, 0.04422636, 
    0.04437408, 0.07167407, 0.08739101, 0.103108, 0.1188249, 0.1345418, 
    0.1502588, 0.1659757, 0.2379444, 0.2365483, 0.2351522, 0.2337562, 
    0.2323601, 0.230964, 0.2295679, 0.1568652, 0.1423967, 0.1279281, 
    0.1134595, 0.09899093, 0.08452235, 0.07005378, 0.04336957,
  0.4133147, 0.325191, 0.08230443, 0.001305809, 0.06698117, 0.05498514, 
    0.03837438, -0.0006227142, 0.0002654412, 7.224286e-05, 0.03841329, 
    0.0863466, 0.2186341, 0.002572999, 0.4273753, 0.4758146, 0.5006552, 
    0.2513014, 0.1020688, 0.2915971, 0.3730793, 0.5479596, 0.1983098, 
    0.0991025, 0.3873709, 0.5807356, 0.08194833, 0.003848597, 0.146693,
  0.0618856, 0.0240012, 0.05780829, 0.01485513, 0.02778129, 0.04654972, 
    0.02863699, 0.06415056, 0.1943218, 0.1426418, 0.1399607, 0.1004046, 
    0.1053123, 0.06065125, 0.1121664, 0.1198873, 0.1395081, 0.09423752, 
    0.1412475, 0.1571319, 0.1462048, 0.2274425, 0.215169, 0.3163348, 
    0.2634415, 0.2917196, 0.1781346, 0.128474, 0.07184406,
  0.09894324, 0.1025794, 0.07781374, 0.09498431, 0.07961793, 0.1446013, 
    0.1704558, 0.1463055, 0.1698212, 0.1720611, 0.1266319, 0.1927101, 
    0.2953509, 0.1907458, 0.140991, 0.1601808, 0.2148927, 0.3077796, 
    0.2963097, 0.2320605, 0.174532, 0.1849003, 0.141397, 0.1036002, 
    0.2613819, 0.3912155, 0.3120486, 0.2727582, 0.1582541,
  0.20593, 0.2223591, 0.1834653, 0.1616367, 0.2000486, 0.1982282, 0.2644175, 
    0.2005699, 0.1524605, 0.1353106, 0.07185958, 0.05014383, 0.1099771, 
    0.1709456, 0.1594839, 0.08913622, 0.07662877, 0.1243265, 0.171098, 
    0.1741978, 0.1337827, 0.0699291, 0.08275931, 0.09291854, 0.02969344, 
    0.1554229, 0.2323121, 0.2133206, 0.2477085,
  0.09203821, 0.04803421, 0.009932174, 0.0186523, 0.05280472, 0.08461659, 
    0.09289549, 0.03387461, 0.04167755, 0.01959454, 0.01383371, 0.006149759, 
    0.006126932, 0.05649783, 0.1156943, 0.01063181, 0.04411924, 0.04479593, 
    0.03278536, 0.03773336, 0.0237189, 0.04308244, 0.02472555, 0.1064936, 
    0.002694165, 0.02059787, 0.02164129, 0.03749225, 0.08686713,
  0.007572849, 0.004658255, 0.001390628, 0.0008949295, 0.003404983, 
    0.03046015, 0.002099397, 0.001224918, 0.003079477, 0.002862472, 
    0.00176613, 9.366134e-05, 0.01204738, 0.003086845, 0.01994975, 
    0.0001319668, 0.005261361, 0.05707183, 0.006431784, 0.002998421, 
    0.002257691, 0.002589996, 0.004977894, 0.01289256, 0.005051082, 
    0.0006916866, 0.001188634, 0.0009159974, 0.0006679016,
  0.01065284, 0.0408573, 1.00102e-05, 0.0002591662, -0.001618481, 
    0.0002728276, 0.0004844653, 0.0008575374, 0.001738922, 0.0003258037, 
    5.125751e-05, -8.298588e-06, 0.0005517351, 0.001258282, 0.000146819, 
    0.001588533, 0.000780933, 0.0001162416, 0.000593143, 0.000206927, 
    0.0002426012, 0.0004907206, 0.001626124, 0.009434399, 0.01304052, 
    0.0601685, 0.0002014923, 0.001420431, 0.002219657,
  0.008437648, 0.004268357, 0.02217556, 0.03175374, 5.375467e-05, 0.00023208, 
    0.0008309299, 4.312418e-05, 0.0009019073, 0.001761929, 0.003984258, 
    0.0005120527, -7.185803e-05, 0.0005743435, 0.0002053755, 0.001382634, 
    0.0008073565, 0.0003767823, 0.0002580652, 0.0007271505, 0.0007934914, 
    0.0008987372, 0.001375772, 0.05392887, 0.02794856, 0.006612704, 
    -6.679767e-05, 0.001148286, 0.002155953,
  0.0007352078, 0.003139923, 6.954789e-05, 0.004254583, 0.0018385, 
    0.001637928, 0.0009798985, 0.0002502821, 0.02847171, 0.06721622, 
    0.0005913202, 0.00135408, 0.000640257, 0.0001933691, 0.000245351, 
    0.0004337642, 0.0005834733, 0.0001616049, 0.0002615099, 0.001355881, 
    0.001032293, 0.00432856, 0.002855167, 0.003880392, 0.01051377, 
    7.686163e-05, 2.143173e-05, 3.915013e-05, 0.001023755,
  2.596678e-09, 1.727426e-08, 1.523308e-09, -1.69851e-05, 0.00573863, 
    0.001989982, -0.0001544007, 0.001255827, 3.384947e-05, 0.0009503767, 
    0.003653856, 3.72075e-05, 5.901072e-05, 3.64915e-05, 0.0002077085, 
    -3.384776e-06, 0.0001107952, 0.0001895397, 0.002318994, 0.001946503, 
    0.0001945924, 0.0002511392, 0.04594811, 0.04748867, 0.000129375, 
    0.001709757, 0.004315392, -2.827888e-08, -0.0004836009,
  2.694175e-09, 7.715067e-10, -4.88792e-11, -1.90248e-06, 2.098683e-10, 
    1.73968e-06, 5.864934e-09, 1.545722e-07, 2.422665e-05, 0.02530053, 
    0.002677115, 0.001893862, 0.00203709, 0.001403654, 0.0009603873, 
    0.0001291841, 0.0008377975, 0.0008807681, 0.00186444, 0.007538048, 
    -4.960392e-07, 0.03484511, 0.0003111299, -0.0004913812, 0.0006938638, 
    0.001541669, 0.004677261, 0.0001046541, 5.998311e-09,
  4.132928e-09, 0.0002412234, 0.002550488, 0.002696793, 0.005517379, 
    7.307519e-07, -0.000246253, 0.06828551, 0.01241879, 0.04230023, 
    0.1030599, 0.03202774, 0.02860999, 0.01990631, 0.03172029, 0.02318531, 
    0.03861976, 0.022864, 0.007402564, 0.02196834, 0.0007558727, 0.05358052, 
    0.01115048, 0.02479786, 0.006021521, 0.00180453, 0.01150997, 0.005117676, 
    -7.968475e-05,
  0.0002823849, 0.001024069, 0.007661661, 0.1827163, 0.003076251, 
    0.001102049, 0.03042889, 7.075039e-05, -1.8271e-05, 0.0003949004, 
    0.06671698, 0.009326392, 0.04846224, 0.0402906, 0.03171273, 0.03667191, 
    0.042441, 0.04748292, 0.03767404, 0.1206919, 0.03078987, 0.0866551, 
    0.0947845, 0.08732544, 0.04525334, 0.06680659, 0.03150994, 0.03135877, 
    0.01048507,
  0.02041244, 0.06230332, 0.03601985, 0.08069906, 0.1153942, 0.1447308, 
    0.04247373, 0.08500963, 0.03800293, 0.001498076, 1.336929e-05, 
    0.04608585, 0.1992485, 0.06324338, 0.04725932, 0.08126986, 0.07908157, 
    0.09534425, 0.04027006, 0.1947871, 0.04587419, 0.04688742, 0.05707113, 
    0.1405149, 0.03550469, 0.1616494, 0.1055171, 0.07566525, 0.07754572,
  0.05854687, 0.2815175, 0.2863168, 0.3640921, 0.2562987, 0.04309608, 
    0.06362785, 0.06646569, 0.05617993, 0.09106847, 0.07254911, 0.3136314, 
    0.2792822, 0.08555736, 0.2124591, 0.14046, 0.2013468, 0.129954, 0.138708, 
    0.1014202, 0.0966429, 0.06617076, 0.181707, 0.2159788, 0.256714, 
    0.01093679, 0.04172485, 0.06732629, 0.05405072,
  0.04974356, 0.02874999, 0.1444801, 0.06317429, 0.3090407, 0.229388, 
    0.4071504, 0.3276231, 0.3757256, 0.3778592, 0.5341885, 0.3001058, 
    0.4598899, 0.2709151, 0.2642812, 0.2770269, 0.3912798, 0.1705562, 
    0.3367313, 0.2547725, 0.2824398, 0.3349193, 0.474186, 0.3082254, 
    0.2318172, 0.1666206, 0.4891961, 0.1256439, 0.1268941,
  0.4344789, 0.2968606, 0.4746775, 0.4553683, 0.4810512, 0.466059, 0.3443489, 
    0.2621819, 0.3536503, 0.3585484, 0.328054, 0.3276007, 0.3258732, 
    0.3293113, 0.3543514, 0.3298614, 0.2577752, 0.2407726, 0.2563136, 
    0.2078545, 0.1836556, 0.1749432, 0.2788354, 0.3033762, 0.08970984, 
    0.04855449, 0.1222915, 0.1935341, 0.3160166,
  0.03229425, 0.0320038, 0.03171334, 0.03142289, 0.03113243, 0.03084197, 
    0.03055152, 0.03545837, 0.04704227, 0.05862617, 0.07021007, 0.08179396, 
    0.09337787, 0.1049618, 0.1594172, 0.1602597, 0.1611021, 0.1619446, 
    0.1627871, 0.1636295, 0.164472, 0.1267747, 0.1146388, 0.1025029, 
    0.09036695, 0.07823104, 0.06609514, 0.05395924, 0.03252662,
  0.3281704, 0.2329517, 0.046025, 0.001871053, 0.001972769, 0.004534637, 
    0.01499961, -0.0005301597, 0.0001361353, 2.404147e-05, 0.02667458, 
    0.07816225, 0.2044905, 0.001660654, 0.3962765, 0.4489796, 0.4351288, 
    0.2508553, 0.09391547, 0.2949523, 0.3623635, 0.5789992, 0.176627, 
    0.09308571, 0.3348231, 0.5518349, 0.07624783, 0.01241625, 0.1335184,
  0.07795954, 0.02156413, 0.04940538, 0.01332291, 0.02678315, 0.03200908, 
    0.02520244, 0.05647907, 0.1749372, 0.1331212, 0.1283445, 0.09201308, 
    0.09775133, 0.05317332, 0.09604651, 0.1018824, 0.1145218, 0.07928704, 
    0.1242467, 0.1358861, 0.1261759, 0.2053936, 0.196184, 0.2859839, 
    0.2326685, 0.2526718, 0.1423847, 0.1049645, 0.06596022,
  0.07965281, 0.08395213, 0.06499428, 0.07731055, 0.06795615, 0.1258023, 
    0.1463962, 0.1245673, 0.1420923, 0.1482671, 0.1068464, 0.1647088, 
    0.247661, 0.1594337, 0.1162042, 0.1333695, 0.1824505, 0.2580588, 
    0.2492112, 0.1842135, 0.1426174, 0.1505518, 0.1084529, 0.08105537, 
    0.2117851, 0.3234096, 0.2617633, 0.2259217, 0.1296981,
  0.1686823, 0.183181, 0.1493863, 0.132442, 0.1687342, 0.169839, 0.2256948, 
    0.1701225, 0.1286833, 0.1103172, 0.05572737, 0.03551749, 0.08732368, 
    0.1371146, 0.1293311, 0.07316814, 0.05963921, 0.09664657, 0.1321513, 
    0.1318853, 0.1076517, 0.05631686, 0.06124621, 0.1030948, 0.0245991, 
    0.1181591, 0.1872068, 0.1820485, 0.2103114,
  0.06752915, 0.03378644, 0.006997772, 0.01092324, 0.03528231, 0.05853719, 
    0.06322101, 0.02483052, 0.02678595, 0.01399978, 0.008896898, 0.004917118, 
    0.004038037, 0.03914184, 0.1189923, 0.006496263, 0.02661894, 0.0270486, 
    0.02262409, 0.02666878, 0.01556184, 0.02922155, 0.01724787, 0.1080194, 
    0.001810885, 0.01523393, 0.01697561, 0.02720112, 0.06534321,
  0.006165334, 0.003824886, 0.01076436, 0.0007418139, 0.002475344, 
    0.01834044, 0.001261269, 0.0009197872, 0.002594254, 0.002347527, 
    0.001173342, 7.02066e-05, 0.01357025, 0.001809413, 0.01121272, 
    0.000109782, 0.003231036, 0.03551681, 0.004188027, 0.002175181, 
    0.001480582, 0.00173759, 0.00404302, 0.01026143, 0.007438989, 
    0.0004188887, 0.0009741026, 0.0007443512, 0.0005331378,
  0.008759402, 0.03161912, -1.585728e-05, 0.0002082722, -0.001901391, 
    0.0002106862, 0.0003794701, 0.0006385323, 0.001368273, 0.0002709983, 
    0.0007778846, -0.0001059208, 0.0004514753, 0.001006024, 0.0001104125, 
    0.00103841, 0.0005807042, 8.985862e-05, 0.0004000125, 0.0001582084, 
    0.000172911, 0.0003979575, 0.001339681, 0.00769252, 0.03342442, 
    0.09098052, 0.0001492658, 0.001131765, 0.001763624,
  0.006902877, 0.002584079, 0.03616905, 0.05618731, 4.623304e-05, 
    0.0001919257, 0.0004475883, 3.410263e-05, 0.0006007644, 0.001003901, 
    0.002737484, 0.000353427, -5.320397e-05, 0.0004720132, 0.0001641948, 
    0.0009407211, 0.0005484508, 0.0002980433, 0.0002099885, 0.0006017603, 
    0.0006468912, 0.0007886664, 0.001130688, 0.08547279, 0.03838727, 
    0.04822414, -0.0002039818, 0.0009507548, 0.001773132,
  0.0005861409, 0.03463187, 0.005532926, 0.005375985, 0.001501733, 
    0.001344091, 0.0008144037, 0.0002029071, 0.03466529, 0.1105607, 
    0.0004405789, 0.001051942, 0.0004483715, 0.0001581981, 0.0002035439, 
    0.0003469242, 0.0004460476, 0.0001389301, 0.0002104966, 0.001065991, 
    0.0007800801, 0.003336715, 0.001904285, 0.04846003, 0.04155423, 
    5.663433e-05, 1.720978e-05, 3.162534e-05, 0.0008283567,
  2.967507e-09, 1.733921e-08, 1.527174e-09, -4.454883e-06, 0.005629466, 
    0.001678982, -0.0006047981, 0.0009652911, -0.0003571638, 0.0007360663, 
    0.002254085, 3.828659e-05, 4.223957e-05, 2.97082e-05, 0.000172494, 
    4.7901e-06, 8.1214e-05, 0.0001556206, 0.001491898, 0.001155578, 
    0.0001432489, 0.0002336458, 0.0549517, 0.03993125, 0.0001113653, 
    0.001430664, 0.003507333, -1.858045e-08, -0.002186154,
  2.709843e-09, 7.675159e-10, -2.114319e-11, -1.564252e-06, 2.371867e-10, 
    1.36297e-05, 6.688288e-09, 1.601104e-07, 0.0002683465, 0.01736467, 
    0.002170086, 0.001431782, 0.001485685, 0.0009112895, 0.0007997192, 
    0.0001084285, 0.0006742488, 0.0006854353, 0.001573124, 0.005338055, 
    -4.133447e-07, 0.0311231, 0.0002626514, -0.000572969, 0.0005773574, 
    0.001209804, 0.003937782, 8.819239e-05, 6.149536e-09,
  4.305313e-09, 0.0002232054, 0.001795285, 0.002003204, 0.005756315, 
    7.110495e-07, -0.0002836532, 0.1242346, 0.02007163, 0.04069807, 
    0.07021849, 0.02106679, 0.01922519, 0.01219361, 0.02163183, 0.01570411, 
    0.02611544, 0.01463939, 0.005929075, 0.01671293, 0.0006271036, 
    0.05308848, 0.01737838, 0.01762097, 0.004019851, 0.001259253, 
    0.009382436, 0.004332606, -4.882011e-05,
  0.0009266661, 0.0008931324, 0.006131385, 0.1961845, 0.002137447, 
    0.0009182582, 0.02814889, 5.16642e-05, -2.122762e-05, 0.0004511109, 
    0.07066745, 0.007677317, 0.0431481, 0.03181244, 0.02670309, 0.03011992, 
    0.03269572, 0.03242305, 0.02550168, 0.1143983, 0.02889099, 0.07717258, 
    0.08123746, 0.07392336, 0.04070649, 0.04767433, 0.02161041, 0.02405449, 
    0.008531393,
  0.01589931, 0.05034441, 0.0329856, 0.08152696, 0.1038594, 0.1350366, 
    0.03772332, 0.140045, 0.08316673, 0.003775838, -0.0002586556, 0.05475875, 
    0.20205, 0.05550145, 0.04249299, 0.06930209, 0.07025183, 0.08229738, 
    0.03004869, 0.1896871, 0.04642839, 0.04923396, 0.06030652, 0.1357754, 
    0.03445141, 0.141414, 0.08923105, 0.05752175, 0.06051692,
  0.04537438, 0.3220799, 0.3064312, 0.3733121, 0.2450316, 0.05833793, 
    0.06049322, 0.08249792, 0.07396369, 0.101288, 0.08577055, 0.4547796, 
    0.3447295, 0.08677843, 0.1943074, 0.1308931, 0.267793, 0.1305157, 
    0.189508, 0.1380807, 0.1120851, 0.09940954, 0.15557, 0.2777962, 
    0.2521189, 0.01771439, 0.03620872, 0.05705667, 0.04364968,
  0.04036144, 0.02369281, 0.1665654, 0.05478959, 0.2967778, 0.2166136, 
    0.4340171, 0.3596736, 0.4593855, 0.4323905, 0.5538243, 0.4246683, 
    0.4874755, 0.2588643, 0.253877, 0.2393709, 0.4421951, 0.2062147, 
    0.3528028, 0.231912, 0.2640193, 0.3041078, 0.4570622, 0.3410618, 
    0.2145783, 0.1529312, 0.4799653, 0.126918, 0.1154268,
  0.5592085, 0.3057052, 0.4377601, 0.3584729, 0.3686694, 0.340239, 0.2481723, 
    0.1782012, 0.3041644, 0.2572384, 0.2495443, 0.2524601, 0.2589349, 
    0.243151, 0.2787147, 0.266274, 0.2055364, 0.2064146, 0.2209338, 0.199676, 
    0.1540809, 0.1746758, 0.292011, 0.3689937, 0.09320294, 0.03754474, 
    0.1524016, 0.2159808, 0.2548968,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.485034e-09, 0, 0, 0, 0, 0, 
    0, 0, 0, -3.246492e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, -1.076182e-05, 2.556325e-05, 0, 0, 0, 0, 
    -8.566196e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -5.138656e-06, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0.0007285672, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 4.999588e-05, 0, 0, 0, 0, 9.641914e-05, 0.0003097472, 0, 0, 0, 
    -7.821295e-05, 0, 0, -3.615231e-05, 0, 0, 0, 0, 0, 0, 0, 0, 
    -4.551592e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, -2.877696e-05, 3.37807e-05, 0, 0, 0, 0, 
    -1.728509e-05, 0, 0, 0, 0, 0, 0, 0, 0, -7.008615e-06, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001040094, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0.003993544, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0.002093571, 0, 0.001163178, -3.838061e-05, -2.56595e-05, 
    0.001052489, 0.001346419, 0, 0.001532482, 0, -0.0002566254, 9.704621e-05, 
    0, -0.0001122286, -4.56766e-06, -5.347972e-06, 0, 0, 0, 0, 0, 0, 
    3.616396e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, -3.521988e-05, 0.0004264705, 0, 0, -2.170417e-06, 
    0.002654377, -2.893667e-05, 0, 0, 0, 0, 0, 0, 0, 0, -7.542227e-05, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -9.17946e-07, -3.975271e-05, 0, 
    0, 0, 0, 0.003274198, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.36831e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, -7.29915e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0.00637093, 0.0001717262, -3.155813e-05, 0, 0, 0, 0, 0, 0, 
    -2.740708e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0.001279755, 0.002154857, -4.35362e-05, 0.002786013, -0.0001347314, 
    -0.0001054202, 0.001235568, 0.003327506, 0, 0.002280885, 0, 0.003294659, 
    0.0001123254, 0, -0.0001863304, -2.308231e-05, -4.269972e-05, 0, 0, 0, 
    -2.129343e-05, 0, -3.379866e-06, 0.0003355876, 0, 0, 0, 0,
  0, -5.455547e-05, 0, 0, 0, 0, 0, 0, -3.604605e-06, 0.001708657, 
    1.448798e-05, 0, -2.580857e-06, 0.005773464, -3.0536e-05, 0, 0, 0, 0, 0, 
    0, 3.176773e-05, 0, -0.0001335704, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -1.667397e-10, 0, 0, 0, 0, 0, -9.989815e-06, 
    -3.767212e-05, -2.591731e-05, -0.0001062378, 0, 0, 0, 0, 0.005416149, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0003033894, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001656693, 0, 0, 0, 0, 
    0, 0, 0, -3.091141e-06, 0, -8.828522e-06, 0, 0,
  0, 0, 0, 0, 0, 0.0004260326, 0.0007301047, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, -8.268952e-09, 0, 0,
  0, 0, 0, 0, 0, 0.01096768, 0.003246588, -7.12322e-05, -1.704513e-05, 0, 0, 
    0, 0, 0, 6.263088e-05, -1.399929e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0.00776963, 0.003814534, -0.0001496131, 0.004586061, -0.0001680775, 
    -0.000299389, 0.001586499, 0.009992118, 0, 0.006923725, -1.399906e-05, 
    0.009011298, 0.001016641, 0, -0.000272429, -4.862208e-05, 8.302368e-05, 
    0, 0, 0, -2.839124e-05, 0, -8.619977e-05, 0.004114926, 0, 0.0002103924, 
    0, 0,
  0, 0.000448022, 0, 0, 0, 0, 0, 0, 6.8523e-05, 0.003716439, 3.877386e-05, 0, 
    0.0004203898, 0.01432426, 0.005855761, 0, -1.04358e-05, 0, 0, 0, 0, 
    8.850409e-05, 0.0001209641, 0.0003313131, -9.741887e-06, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -3.001605e-05, 0, 0, 0, 0, -2.412765e-05, -2.880889e-05, 
    -0.0002096914, 0.001141134, 0.00131145, 0, 0, 0, -2.44379e-05, 
    0.008137124, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0009244148, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -1.756689e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.336521e-08, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0.0001153057, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001730457, 
    0.0003814468, 0, 0, 0.0001249836, 0, 0, 0, 9.542184e-05, 0.000334461, 
    9.414736e-05, -2.647029e-05, 0,
  0, 0, 0, 0, 0, 0.00385098, 0.003961901, 0, 0, -1.04457e-06, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.002229405, 0, 0, 0, 0, 0, 0, 8.091964e-05, 0.0005501967, 0, 0,
  0, 0, 0, 0, 0, 0.02523786, 0.007155993, -0.000131711, -8.283863e-05, 0, 0, 
    0, 0, -4.239952e-05, 0.0003399289, 0.0003911396, -1.718575e-05, 
    -1.573613e-05, 0, -2.29288e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0.0112377, 0.003851037, -0.000255449, 0.005807656, -0.0001378546, 
    0.001566646, 0.00184782, 0.01691089, -4.252608e-05, 0.00933635, 
    0.001180973, 0.01564445, 0.002164277, -5.138073e-06, 0.001956732, 
    -0.0001117519, 0.0001073418, 0, 0, 0, -5.678249e-05, 0, -0.0001767042, 
    0.008250466, 0, 0.002813668, 0, 0,
  0, 0.001890984, 0.0004995788, 0, 0, 0, 0, 0, 0.0004209651, 0.00883113, 
    6.264244e-05, -2.081162e-05, 0.004798957, 0.01996881, 0.009076185, 0, 
    -2.250185e-05, -3.08142e-05, 0, 0, 0, 0.0004383225, 0.003089899, 
    0.002778736, 0.0006333336, 6.984469e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -0.0001129104, -1.261339e-05, 0, 0, 0, -0.0002623762, 
    -0.0001332493, -0.0001930383, 0.004045258, 0.006105739, -3.069651e-05, 0, 
    0, -2.956709e-05, 0.01829189, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.00126321, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001381229, 0.001446261, 0.0006319294, 
    2.165418e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0008126286, -5.805005e-05, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.055983e-05, 0.0004214199, 0, 0, 
    -1.851177e-06, 0, 0, 0, 0, 0, 0, 0, -1.589439e-07, -2.168994e-06, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9.059507e-07, 0, 
    -4.484294e-06, 0, 0, 0, 0, 0, 0, 0, -4.957259e-06, 0,
  -1.014845e-05, 0, 0, 0.00154455, 0, 0.0002705977, 0, 0, 0, 0, 
    -2.410607e-05, 0, 0, 0, 0, -5.410947e-05, 0.004172671, 0.002022727, 
    -0.0001310918, 0, 0.001881923, 0, 0, 0, 0.001108291, 0.0026533, 
    0.005638597, 0.00152375, 0,
  0, 0, -1.968753e-06, 0, 0, 0.01017006, 0.006865554, 0, 0, -1.516374e-05, 0, 
    0, -2.018912e-06, -2.926515e-06, 0.002489924, 0, 0, 0.0002667526, 
    0.007971463, 0, 0, 0, 0, 0, -2.949862e-05, 0.001405403, 0.001715544, 0, 0,
  0, 0, 0, 0, 0, 0.03688605, 0.009665408, 0.0001396066, 4.912672e-05, 0, 0, 
    0, 0, 0.0007141344, 0.005207636, 0.0008190995, -4.713318e-05, 
    -8.845769e-05, 0, -4.784665e-05, 0, 0, 0, 0, -1.927172e-06, 0, 0, 0, 0,
  0, 0.01860293, 0.009674885, -0.0001659337, 0.008237144, -6.330404e-05, 
    0.005342942, 0.002154211, 0.03431381, -6.378913e-05, 0.01425433, 
    0.002021871, 0.02914177, 0.006171478, 6.160678e-05, 0.007178829, 
    -0.0003044504, 0.0004261953, 0, 0, 0, -0.0001905889, 0, 0.001099283, 
    0.01193366, 0, 0.004038182, -4.914607e-06, 0,
  0, 0.004374609, 0.0005782791, 0, 0, 0, 0, -9.371624e-06, 0.0004289882, 
    0.01600778, 0.0004510845, 3.967363e-05, 0.009873265, 0.03198227, 
    0.01663854, -1.061691e-06, -4.112582e-05, -0.0001456235, 0, 0, 
    9.339937e-06, 0.005001743, 0.005688816, 0.01017548, 0.001042677, 
    0.0002825668, 0, 0, 0,
  0, 0, 0, -2.013302e-05, 0, 0, -0.0003576754, -2.893934e-05, 0, 0, 
    3.055919e-07, -0.0001005845, 0.00099688, 0.003599873, 0.007594375, 
    0.01590409, -0.0001598852, -2.20169e-05, 0, 0.0001070688, 0.02885377, 0, 
    0, 0, 0, 0, 0, -1.395346e-07, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.00237019, 0, 0, 0, 0, 0, 0, 
    -7.761112e-05, 0, 7.858493e-05, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0.008024498, 0.0074294, 0.002485448, 
    0.001724553, 0, 0, 0, 0, 0, 0, 0, 0, -1.679927e-05, 0.001613971, 
    0.0004053866, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0009348916, 0.00235605, -5.758977e-05, 
    6.578447e-07, 0.001160734, 0, 0, 0, 0, 0, 0, -1.662895e-05, 0.0002646075, 
    0.0002119991, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -8.823789e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0.0001338734, 0, 0, 0, 2.661925e-05, 0, 0, 0, 0, 0, 0, -8.587311e-05, 0, 0, 
    0, 2.302609e-05, -2.130918e-05, 0.000131958, 0, 0.001538688, 0, 0, 
    0.0002893094, 0, 0, -9.071608e-06, -0.0001492811, 0.001311992, 
    1.380779e-05,
  -0.0001552895, -1.539372e-05, 0, 0.004382615, 0.001180924, 0.005239136, 
    -3.503501e-05, 0, 0, 0.0004437559, 0.0003822777, 0, 0, 0, -6.378717e-06, 
    -0.0001926506, 0.01111688, 0.006467111, 0.002210864, -8.939925e-06, 
    0.009737215, 0, -1.071152e-05, 0, 0.002285004, 0.009191545, 0.01037723, 
    0.006101168, -1.431427e-05,
  0, 0, -3.690706e-05, 0.0003796487, 8.875579e-05, 0.01380066, 0.01719707, 0, 
    -2.160474e-06, 0.0009864391, 0, 0, -7.101209e-05, -0.0002159024, 
    0.007282651, 5.620605e-07, -1.727512e-06, 0.004307816, 0.02035487, 0, 
    0.001328339, 0, 0, 0, -8.547419e-05, 0.004346741, 0.003709425, 
    1.578847e-06, 0,
  0, -5.722289e-06, 0, 0, 0.0003284574, 0.05269423, 0.01213475, 0.00131014, 
    0.002714224, 0, 0, 0, 0, 0.004944792, 0.02332216, 0.005770362, 
    -6.693108e-05, 0.0009833493, -2.092486e-05, 2.515456e-05, -2.891281e-05, 
    0, 0, 1.852358e-09, 0.00102901, 0, 0, 0, 0,
  0, 0.03944391, 0.015732, 0.002621645, 0.01471965, 8.665826e-05, 0.01018083, 
    0.004068902, 0.06022494, -0.0001722255, 0.01673658, 0.008088783, 
    0.04567088, 0.01466348, 0.0005243767, 0.01115049, -0.0001835688, 
    0.001567802, 0, 0, 0, -0.000243758, 0, 0.003502421, 0.0215355, 
    -9.501437e-06, 0.005423149, -6.343603e-05, 0,
  0, 0.007301294, 0.0009678343, -9.36318e-06, 0, 0, 7.60074e-07, 
    0.0002380434, 0.003543693, 0.02495847, 0.006771569, 0.002861182, 
    0.01783156, 0.05984172, 0.02711874, -7.819791e-07, -8.89732e-05, 
    -0.0001144203, 0, 0, -5.63548e-05, 0.01237088, 0.008980982, 0.02469967, 
    0.002598349, 0.001235197, 1.622869e-06, 0, 0,
  0, 0, 0, -3.803798e-05, -5.03481e-06, 5.454029e-06, -0.0003004926, 
    -0.0001074623, 1.456831e-05, -8.170949e-06, -6.968987e-06, 0.007353322, 
    0.004108368, 0.01339349, 0.01301967, 0.02593487, 0.002485421, 
    -9.543481e-05, -2.525008e-06, 0.000385728, 0.05504544, -0.0001063283, 
    -1.028343e-07, 0, 0, 0, 0, -5.871854e-05, -7.797236e-06,
  0, 0, 0, 0, 0, 0, 3.99861e-05, 0, 2.894987e-05, 0, 0, 0.007970657, 
    -4.238264e-08, -1.199089e-07, 0, 0, 0, 0, 0.001136296, 0.0001981956, 
    0.0003264449, 0, -6.182905e-06, 0, 0, 0, 0, -1.444342e-05, 0,
  0, 0, 0, 0, 0.0007940144, -1.241152e-05, 0, 0, 0, 0.01505642, 0.02461683, 
    0.0040908, 0.01092637, -3.102589e-05, 0, 0, 0, 0.0001323764, 0, 0, 0, 
    -4.560873e-05, 0.00280418, 0.002729267, 2.541305e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.005647028, 0.008891705, 0.0007339765, 
    0.003051614, 0.003567175, 0, 0, 0, 0, 0, 0, -9.455567e-05, 0.003857597, 
    0.001815103, 6.698367e-05, 3.347422e-05, 3.524648e-05, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -2.814296e-05, 0, -5.342902e-07, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.001052739, 0, 4.932472e-06, 0, 0.0009103072, -5.119084e-05, 0.003586339, 
    0, 9.435146e-06, 0, 0, 0.0001144514, 5.053773e-05, 0, 0, 0.001465079, 
    0.004202397, 0.001076696, -2.685172e-06, 0.005752388, 0.006724585, 
    0.00360618, 0.006836544, 0, 0, -0.0001170628, 0.0003487081, 0.004098913, 
    0.004613041,
  0.0003967503, 0.000738097, -2.474248e-07, 0.008121273, 0.002844567, 
    0.007817262, -5.766032e-05, 0, 0, 0.005517207, 0.006498534, 0, 0, 0, 
    -3.423747e-06, 0.001890402, 0.01678001, 0.01954354, 0.0399155, 
    0.008862378, 0.0204488, 0.003860941, 0.0006333169, -0.0001089404, 
    0.006500505, 0.02774813, 0.01650192, 0.01574222, -0.0001335151,
  0, 0, -8.898524e-05, 0.006057976, 0.001975128, 0.02100982, 0.03047643, 0, 
    0.0001499818, 0.008473373, 0.001258323, 0.000302686, 0.00296116, 
    -0.0001038235, 0.01402071, 0.002555108, 0.00418543, 0.01618293, 
    0.03588159, 0.0004260322, 0.006738356, -3.323648e-05, 0, 0, 3.350196e-05, 
    0.006895218, 0.01167643, 0.005517459, -5.848724e-06,
  0, -1.053196e-05, 0, 0, 0.0004063573, 0.07475523, 0.01896167, 0.003695997, 
    0.0106023, -8.351348e-06, 5.882466e-07, 7.503902e-05, -3.575189e-09, 
    0.007975828, 0.03599837, 0.02334446, 0.003969756, 0.005743453, 
    0.006675391, 0.0002278986, -6.132473e-05, 0, 0, 4.341022e-06, 
    0.003121893, -6.270095e-06, -1.402502e-05, 0, 0,
  0, 0.06370898, 0.02343529, 0.01423565, 0.03018553, 0.02374813, 0.02763873, 
    0.01719783, 0.08689652, 0.003394184, 0.02355967, 0.009689189, 0.07745918, 
    0.04046712, 0.00416156, 0.0264127, 0.00537655, 0.0119378, 0.001512813, 0, 
    -0.0001052769, 0.0003826639, 5.325699e-09, 0.01911197, 0.03432807, 
    0.0002908017, 0.005141504, -0.0001414279, 0,
  0.0005471584, 0.02520316, 0.005028463, -1.634373e-05, -5.588255e-06, 
    -8.747125e-06, -7.596303e-06, 0.003898886, 0.03979839, 0.05168647, 
    0.02497412, 0.0153836, 0.05348317, 0.1083102, 0.04437036, -9.032919e-06, 
    -0.000219499, 0.003153065, 8.92412e-07, 0, 0.002867622, 0.0232737, 
    0.01992912, 0.06022201, 0.006256063, 0.002084892, 9.042954e-05, 0, 
    -3.651564e-06,
  2.385731e-06, 2.532595e-05, -1.236456e-05, 5.957644e-05, -2.472056e-05, 
    0.002220235, 0.01253928, 0.001281067, 0.0004151897, 0.004482392, 
    -8.056981e-05, 0.02207487, 0.03146242, 0.03164008, 0.01980561, 
    0.04803661, 0.01091672, 1.690142e-05, 0.0003536752, 0.001501187, 
    0.08293277, -1.641308e-05, -1.818294e-06, 0, 0.000374045, 0, 0, 
    0.0004719211, 0.001580102,
  0, 0, 0, 0, 0.000259642, 0, 1.13257e-06, -1.426653e-07, 4.556547e-05, 
    -8.598949e-12, -1.186891e-06, 0.02351848, 0.00030826, 0.0005669466, 
    0.0005971268, -7.7284e-07, -3.312901e-05, -5.366311e-10, 0.003958281, 
    0.008716203, 0.003680162, 6.561683e-05, -3.041374e-05, 2.351982e-07, 0, 
    0, 0, 0.000127173, -3.096858e-07,
  0, 0, 0, 0, 0.002647772, -7.084305e-05, 0, 0, 0, 0.02893708, 0.0511699, 
    0.006400778, 0.02312928, 0.0001396252, -1.321192e-05, -4.529255e-05, 0, 
    0.00313064, -1.390959e-05, 0, 0, -0.000107518, 0.007339668, 0.004130009, 
    0.00225982, 0.0002904439, 6.651307e-05, 0, 0,
  0, -1.899715e-06, 0, -7.612105e-06, -2.82676e-05, 0, -9.999123e-06, 0, 0, 
    -1.50226e-06, 0.007344054, 0.01680281, 0.002683507, 0.00769715, 
    0.007383033, -2.129366e-05, -8.192425e-07, 0, 0, 0, 0, -0.0002303479, 
    0.006593557, 0.009668436, 0.001671241, 0.004051333, 0.001845667, 0, 0,
  0, 8.992342e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001801685, 0, 0, 0, 
    0, 0, 0, -7.128921e-05, 0, 0, -3.49322e-06, -6.576439e-06, 0, 
    2.158257e-05, 0,
  -3.235816e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.0008906731,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -4.847596e-05, 0, 0.0007735137, 0, 0, 0, 0, 
    0.0003225558, 0.0007441441, 0.0004800179, 6.734907e-05, 0.0008784088, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0.002188033, 4.511376e-06, 0.0005486897, -9.581126e-05, 0.004477536, 
    0.001097633, 0.007435302, 0.003221446, 0.004895935, -1.501576e-05, 
    -5.887101e-07, 0.005290811, 0.0004390421, 0, -1.368023e-05, 0.004898008, 
    0.01092757, 0.003287286, 0.006328184, 0.0134355, 0.01441375, 0.01113153, 
    0.01197654, 0.002619887, 1.37223e-05, 0.002032721, 0.002386837, 
    0.01263779, 0.01016922,
  0.001454952, 0.007164619, -2.579295e-05, 0.01410897, 0.007603526, 
    0.01137768, 2.833212e-05, 1.65873e-05, -3.433528e-06, 0.00782722, 
    0.01295568, 0.000656047, -1.004764e-05, 0.002531938, 0.002710676, 
    0.006842597, 0.0330354, 0.02883323, 0.0859405, 0.03543806, 0.04510303, 
    0.007668802, 0.001564669, 0.0008373857, 0.01665157, 0.05030054, 
    0.02726859, 0.02865578, 0.008191188,
  0, -8.333712e-10, -4.103296e-05, 0.01836651, 0.004828392, 0.02037544, 
    0.04078734, -1.188254e-07, 0.00575721, 0.01734138, 0.005519402, 
    -3.544445e-05, 0.00426054, 0.009154859, 0.02222547, 0.02350326, 
    0.03212266, 0.04863106, 0.08123291, 0.004089771, 0.0226199, 0.001394414, 
    0.003698851, 0.009060415, 0.0002767628, 0.0112734, 0.03134735, 
    0.007868349, -4.077496e-05,
  5.194976e-06, -3.648635e-05, 2.04605e-05, 1.087985e-05, 0.007050085, 
    0.08541027, 0.05273192, 0.009123942, 0.01941327, 0.0002768801, 
    0.001101715, 0.001008342, 3.801525e-05, 0.01276524, 0.08238009, 
    0.08722995, 0.04020527, 0.01978356, 0.02257596, 0.001131354, 0.002276185, 
    -6.45407e-07, -4.697625e-08, 0.01477607, 0.01334189, 0.0001993643, 
    0.00140428, 2.774786e-05, -1.555701e-06,
  -1.298573e-06, 0.1087094, 0.05944592, 0.02684403, 0.04272167, 0.1362699, 
    0.06758991, 0.05812573, 0.2072114, 0.03975962, 0.0496745, 0.01196756, 
    0.1495907, 0.2071189, 0.09931879, 0.07206908, 0.09210348, 0.07306165, 
    0.01592523, 2.474543e-05, 0.0005594956, 0.006634868, 2.759525e-05, 
    0.08025458, 0.0970512, 0.003165679, 0.01078912, 0.0006142832, 3.321718e-08,
  0.01537642, 0.05319509, 0.05341812, -7.161202e-05, 5.235997e-05, 
    4.030169e-05, 0.0005096547, 0.01489816, 0.136129, 0.1125159, 0.1255882, 
    0.1017143, 0.2392196, 0.2025539, 0.1118978, 0.000275532, 0.0001983633, 
    0.004966384, -2.647666e-05, -3.608492e-05, 0.008963615, 0.04147898, 
    0.0406314, 0.1790289, 0.03734039, 0.006556999, 0.002234063, 3.99278e-05, 
    0.004418625,
  0.0005689692, 0.001353286, 0.0002581656, 0.001954945, -0.0002124817, 
    0.009705206, 0.07605492, 0.01934263, 0.03069313, 0.02562873, 0.00789363, 
    0.04419335, 0.180221, 0.1256023, 0.07311858, 0.09165447, 0.04253443, 
    0.009176728, 0.001160009, 0.007980877, 0.1184573, 0.02922113, 
    -0.0002058747, 0.0001382279, 0.009394668, -2.45263e-05, 0.0001461575, 
    0.005133446, 0.02371191,
  0.0001097385, -1.984943e-06, -1.163672e-05, 0.0006289951, 0.0007896781, 
    -1.283657e-07, 8.795138e-05, 0.000866082, 0.001350224, 0.0009044328, 
    0.001429116, 0.0328918, 0.01029726, 0.003868904, 0.007610579, 
    2.683293e-05, 0.001051794, 2.970902e-06, 0.007162238, 0.01565335, 
    0.02094913, 0.004904816, 0.0002436305, -4.145568e-06, -3.032854e-06, 
    -5.118592e-11, -1.431508e-07, 0.00359066, -5.122052e-05,
  0, 0, 0, 7.296079e-07, 0.004141106, 0.002506291, -3.235243e-09, 0, 0, 
    0.05356724, 0.08154403, 0.02633613, 0.03302787, 0.00544685, 0.005702453, 
    0.003050422, 0.001634051, 0.005772716, 0.0002280429, -3.534165e-05, 0, 
    0.001255397, 0.0100038, 0.008780154, 0.008687327, 0.003784995, 
    0.0006870685, 0, 0,
  0, -2.266867e-05, 0, 0.0004452229, 5.020208e-05, -1.106462e-06, 
    0.001856828, 0, -9.120237e-06, -4.404406e-05, 0.01121879, 0.02259219, 
    0.01109246, 0.01902594, 0.01572324, 0.002836202, 0.0009356753, 
    -2.781135e-06, 0, 0, 0, 0.002134692, 0.01302997, 0.03009219, 0.007095271, 
    0.0061696, 0.003552955, 0, 0,
  0, 0.001722189, 0, 0.0005109409, 0, 0, 0, 0, 0, 0, 0, -1.809633e-05, 
    -2.550248e-05, 0, 0.007216093, -4.83073e-06, 2.464031e-05, 0, 0, 0, 0, 
    0.002031569, 0, 0.0006342367, 0.003241668, 0.002617512, 0.001301415, 
    0.003731555, 0,
  0.001125417, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.003988448,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -6.466018e-05, 0, 0, 0, 0, 
    -2.387719e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, -7.338178e-06, -1.512988e-05, 0, -6.976363e-06, 0, 0, 
    0.0004096905, -0.000122308, 0.002804843, 0, 0, 0, -8.357383e-09, 
    0.002360157, 0.005343625, 0.007351507, 0.000217198, 0.003001333, 0, 0, 0, 
    0, 0, 0, -1.015483e-07, 0,
  0.0153071, 0.003190958, 0.005663936, -0.0005136058, 0.02291962, 
    0.007546755, 0.01549668, 0.01046956, 0.0087118, 0.0005850169, 
    0.0001116768, 0.008836514, 0.01381668, 8.426401e-05, 0.001177239, 
    0.01145706, 0.0200104, 0.01127868, 0.05287353, 0.0213645, 0.01974666, 
    0.02188873, 0.01852565, 0.00528559, 0.00316158, 0.003208696, 0.004082414, 
    0.02018315, 0.02132276,
  0.02577194, 0.01207623, 0.0005640595, 0.02586294, 0.0155384, 0.02077522, 
    0.004007919, 0.005693837, -2.455855e-05, 0.01914191, 0.02282103, 
    0.009007861, 0.000531221, 0.0096008, 0.0137438, 0.01882113, 0.0669585, 
    0.04056891, 0.1490406, 0.07902487, 0.09748942, 0.02521665, 0.004365263, 
    0.01052368, 0.027565, 0.07281623, 0.03931133, 0.05783562, 0.03016261,
  0.004281245, 0.001430922, 0.0001948136, 0.02866568, 0.01247577, 0.03698288, 
    0.1006291, 0.02625348, 0.0285272, 0.1147693, 0.02817026, 0.004317607, 
    0.007738268, 0.02141559, 0.05838323, 0.06695248, 0.116915, 0.1014919, 
    0.2341615, 0.09454951, 0.05562446, 0.02922866, 0.008594955, 0.01466872, 
    0.01787139, 0.0968828, 0.1117553, 0.0523659, 0.01564552,
  2.808287e-05, 0.002145813, 0.06042678, 0.005272023, 0.107341, 0.1609636, 
    0.1274801, 0.05388085, 0.04394514, 0.1021033, 0.008593163, 0.01348878, 
    0.01358927, 0.03428802, 0.0945465, 0.09090187, 0.04895661, 0.09423009, 
    0.1740605, 0.05639961, 0.05981422, 0.01311183, 0.001766149, 0.1228254, 
    0.05745155, 0.08685367, 0.1152116, 0.1077918, 0.02518031,
  0.0007221036, 0.2123719, 0.3527522, 0.069961, 0.09518358, 0.1299446, 
    0.09851802, 0.06927595, 0.2279803, 0.0558659, 0.05956604, 0.01300342, 
    0.1355023, 0.1897791, 0.08197081, 0.05681812, 0.1014372, 0.1805142, 
    0.1053339, 0.03150824, 0.04760251, 0.05293217, 0.01905197, 0.2362144, 
    0.195476, 0.06385768, 0.05662973, 0.1966085, 0.00207524,
  0.0398645, 0.3638911, 0.3185783, 0.0006328349, 0.003580101, 0.004925439, 
    0.0198546, 0.08510333, 0.4350002, 0.3060071, 0.149426, 0.09515287, 
    0.2266015, 0.1874137, 0.07462278, 0.00152142, 0.002276625, 0.03308146, 
    0.03226984, 0.002433488, 0.02488862, 0.06616664, 0.0506713, 0.2913481, 
    0.1947344, 0.06183409, 0.09385774, 0.01859531, 0.00495961,
  0.03141965, 0.1204208, 0.002983795, 0.01287706, 0.01134496, 0.03224247, 
    0.1402432, 0.06678167, 0.039439, 0.0329995, 0.007126796, 0.05100972, 
    0.174913, 0.1000786, 0.08952221, 0.09959614, 0.06672533, 0.06985895, 
    0.1189534, 0.118705, 0.2447945, 0.04153023, 0.0003650019, 0.02292198, 
    0.04407236, 0.0342506, 0.08070368, 0.0632188, 0.2075653,
  0.07018337, 0.003301812, 0.0002913239, 0.000839502, 0.03404761, 
    0.002236589, 0.03486946, 0.06514599, 0.0803241, 0.006434808, 0.01963809, 
    0.0381975, 0.01507133, -0.0001113907, 0.02955035, 0.005060911, 
    0.009141345, 0.01329116, 0.07793743, 0.09168784, 0.18466, 0.0990724, 
    0.02726753, 0.02985968, 0.0217106, -4.533246e-06, 0.003872496, 
    0.007437197, 0.03019292,
  -2.605425e-05, -1.935233e-06, 6.01002e-05, 0.000403211, 0.005698193, 
    0.0103836, 7.012575e-06, -4.111494e-08, -2.263596e-05, 0.0937851, 
    0.1243484, 0.1005986, 0.06421234, 0.02560216, 0.030596, 0.02029456, 
    0.01960714, 0.04887085, 0.006904026, 0.007315175, -8.99724e-05, 
    0.01920668, 0.01977839, 0.03418035, 0.01760971, 0.01316223, 0.005862939, 
    -2.309117e-11, -2.686825e-05,
  3.019399e-05, 0.0003531223, -3.467394e-05, 0.001189559, 0.002244062, 
    -5.337517e-05, 0.003466548, -3.093177e-05, -4.260182e-05, 0.0009993589, 
    0.01589388, 0.03098153, 0.02618119, 0.04706667, 0.03342604, 0.00838495, 
    0.003158988, 0.001487474, 0.0002425773, 0, 0, 0.007215978, 0.01950831, 
    0.06190494, 0.02000213, 0.01716358, 0.004670221, 0, -2.648658e-05,
  -9.71741e-06, 0.002463761, -3.975294e-06, 0.001600983, 0, 0, 0, 0, 0, 0, 0, 
    -7.06685e-05, 0.001354095, 0, 0.01062453, -4.863534e-05, 0.0008462894, 0, 
    0, 6.906363e-06, -1.049738e-05, 0.002880475, 0.0003356875, 0.005166268, 
    0.008417885, 0.009862798, 0.004064833, 0.008777053, 0,
  0.005813634, 0.00100247, 0.003149924, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, -3.697359e-06, 8.125829e-05, -3.84582e-06, 0, 
    0.002915355, 0.003805568,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -9.366551e-05, -0.0001727986, 0, 0, 0, 
    -0.0001111364, 0.002879295, 0.002735368, 0.0004702761, 0, 0, 0, 
    1.136417e-06, 0, 0, 0, 0,
  0, 0, 0, 0.002606448, 0.0002082764, 0.0005174834, 0.000111836, 
    -8.701964e-06, 0.0002476332, 0.002417862, 0.0003803007, 0.004182982, 
    0.003890716, 0.000908475, 9.677213e-05, 0.000182516, 0.007850545, 
    0.01189903, 0.01694914, 0.008340104, 0.01393776, 0.003814568, 
    -7.926756e-06, 0.001023596, 0, 0, 0, 0.001493284, 0,
  0.04056008, 0.03885799, 0.03750912, 0.0106468, 0.03769756, 0.03319881, 
    0.03479358, 0.04590266, 0.02049792, 0.01456645, 0.003718711, 0.01920985, 
    0.02483036, 0.00134628, 0.005510727, 0.02455701, 0.05459892, 0.0303517, 
    0.05343572, 0.05681355, 0.05596664, 0.05312205, 0.04768086, 0.01446347, 
    0.01124112, 0.004668364, 0.01734621, 0.04419599, 0.04095393,
  0.06544193, 0.04085103, 0.02284942, 0.05355667, 0.08079004, 0.05087473, 
    0.03055369, 0.02439769, 0.01247053, 0.03207155, 0.07222778, 0.06505613, 
    0.02324466, 0.01320486, 0.029875, 0.05582129, 0.1425694, 0.09032136, 
    0.1593068, 0.1818933, 0.1872288, 0.06959879, 0.04185797, 0.04791368, 
    0.07573456, 0.1139509, 0.07539768, 0.1064922, 0.1218068,
  0.03362719, 0.03737651, 0.003730833, 0.08475195, 0.05026999, 0.1172017, 
    0.166228, 0.08123715, 0.05632417, 0.1600637, 0.173889, 0.09782238, 
    0.0367145, 0.07098966, 0.08320598, 0.1397136, 0.1582988, 0.1471127, 
    0.2299253, 0.1366375, 0.1652104, 0.07585712, 0.0312994, 0.01203168, 
    0.03844284, 0.1312037, 0.1438868, 0.1265105, 0.05695173,
  0.0001487666, 0.0006837437, 0.1296895, 0.003418163, 0.080742, 0.1340594, 
    0.1141405, 0.05130906, 0.05357423, 0.1001451, 0.01418306, 0.01257324, 
    0.008712052, 0.0503328, 0.09657127, 0.08224764, 0.03524512, 0.05921562, 
    0.1536716, 0.05373, 0.0650568, 0.002386143, 0.002450549, 0.1060421, 
    0.04505151, 0.09538232, 0.1096553, 0.1427206, 0.02488985,
  8.354471e-05, 0.2167331, 0.3258397, 0.04625822, 0.07011819, 0.08817737, 
    0.07555539, 0.05178574, 0.2000408, 0.04909672, 0.04746949, 0.0144539, 
    0.1163014, 0.1535273, 0.05414622, 0.04229669, 0.06498785, 0.1332618, 
    0.05390162, 0.0149318, 0.02471328, 0.03725974, 0.005466528, 0.1877942, 
    0.182112, 0.04217367, 0.04248668, 0.1314114, 0.0001992755,
  0.02313015, 0.3272346, 0.2574717, 0.0006320434, 0.004292853, 0.003459554, 
    0.008256165, 0.04649179, 0.3561434, 0.2575711, 0.1064737, 0.07737036, 
    0.1683348, 0.1672312, 0.05885669, 0.000982356, 0.002538341, 0.02443572, 
    0.0250286, 0.0003170519, 0.01411569, 0.05117246, 0.06201356, 0.2637425, 
    0.1536581, 0.05331955, 0.05878426, 0.004855219, 0.003782517,
  0.02646312, 0.07366373, 0.0001191223, 0.08060517, 0.007432353, 0.02222372, 
    0.08742005, 0.03481968, 0.02123559, 0.01889532, 0.003360871, 0.04438995, 
    0.160703, 0.08050915, 0.0690503, 0.08866507, 0.08648629, 0.0437978, 
    0.06046307, 0.06241701, 0.199016, 0.0237031, 0.001227549, 0.009933821, 
    0.03389584, 0.004824749, 0.06391294, 0.01688428, 0.1714428,
  0.1228941, 0.02037526, 0.003092251, 0.000130345, 0.05915733, 0.0003284689, 
    0.02165209, 0.02435521, 0.06591458, 0.007304425, 0.01872968, 0.03356834, 
    0.02734289, 0.003761609, 0.03204992, 0.001451769, 0.01044433, 
    0.003477238, 0.07092001, 0.08701567, 0.1699117, 0.07797489, 0.02726558, 
    0.05436873, 0.02814364, 0.08293957, 0.06367938, 0.03888096, 0.07658943,
  0.0129141, 0.007623015, 0.003641271, 0.005432676, 0.02352813, 0.05661905, 
    0.01085686, -1.968244e-05, 4.04557e-06, 0.1375965, 0.1765275, 0.1934884, 
    0.1454566, 0.1009692, 0.1014558, 0.08917625, 0.08210728, 0.06397281, 
    0.03706082, 0.03597309, 0.005241614, 0.08233354, 0.1656094, 0.1227286, 
    0.1275084, 0.1280349, 0.03402922, 0.002085761, 0.01268513,
  5.05989e-05, 0.0005204388, 0.005970816, 0.006352365, 0.007966707, 
    0.0001261899, 0.006957766, 0.000101149, -7.170378e-05, 0.005383173, 
    0.03437432, 0.04507741, 0.04418517, 0.1549246, 0.1365037, 0.0650266, 
    0.02162369, 0.03886305, 0.04513725, -8.481068e-05, 6.614178e-05, 
    0.01366588, 0.03176266, 0.1110813, 0.0539455, 0.05744764, 0.02166191, 
    0.01651238, 0.00267035,
  0.002118741, 0.005742295, -9.66009e-05, 0.001678122, -2.037715e-05, 0, 0, 
    0, 0, 0, 0, -0.0002024698, 0.01339096, 0.002999831, 0.01498579, 
    0.004564352, 0.00454629, 1.968837e-05, -4.093688e-05, 0.002931649, 
    0.0002009817, 0.005197454, 0.001730315, 0.01301226, 0.04830937, 
    0.03395068, 0.03178941, 0.0193606, 0.0001026555,
  0.01363548, 0.00609701, 0.00999532, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, -3.337623e-05, -3.003527e-05, -0.0002044526, 
    9.31871e-07, 0.004147476, 0.005037189,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.537926e-05, 
    -5.432936e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0001041952, -0.0002823269, 
    -4.185725e-05, 0, -3.876044e-10, 0.003370223, 0.01011869, 0.01852971, 
    0.02070612, 0.009022512, -6.531382e-07, -7.013985e-05, 0.000124547, 
    -2.20726e-06, 0, 0, 0,
  0.002000751, 0.001505339, 0, 0.006799038, 0.01489137, 0.01181913, 
    0.0181832, 0.0006353201, 0.006757968, 0.01341216, 0.02258821, 0.01732053, 
    0.0193562, 0.01376699, 0.004668769, 0.004603702, 0.03994789, 0.06183684, 
    0.0662685, 0.06144564, 0.0731599, 0.0150752, -0.0002309673, 0.003854458, 
    0.0003564929, 0.00357756, 0.003248567, 0.003285372, 0.0006752349,
  0.1286941, 0.1132046, 0.1222071, 0.03275544, 0.07857957, 0.135518, 
    0.1090766, 0.1170536, 0.03240661, 0.03752423, 0.06461477, 0.08543354, 
    0.08512143, 0.07465186, 0.06014847, 0.07725161, 0.1073484, 0.06595453, 
    0.05909108, 0.08210821, 0.1273726, 0.1082132, 0.0919184, 0.03227255, 
    0.03792039, 0.02664558, 0.03294001, 0.09712377, 0.109735,
  0.1341036, 0.1234684, 0.09758458, 0.13103, 0.1862142, 0.1020414, 
    0.07040783, 0.05252267, 0.05263256, 0.1198884, 0.1468627, 0.1075021, 
    0.06834773, 0.07307993, 0.06818755, 0.104247, 0.1759143, 0.1641555, 
    0.1645275, 0.1771515, 0.22887, 0.1195017, 0.08737142, 0.09061221, 
    0.1538246, 0.1916904, 0.1349768, 0.1673646, 0.178792,
  0.03363721, 0.02816953, 0.08862773, 0.07090446, 0.03787005, 0.1164115, 
    0.1483704, 0.08650079, 0.05700575, 0.1587428, 0.2108568, 0.1171252, 
    0.1086966, 0.07543425, 0.07721619, 0.1211704, 0.1415178, 0.1040759, 
    0.2027342, 0.1435599, 0.1345334, 0.03891171, 0.02882608, 0.01092327, 
    0.0194729, 0.113163, 0.1221207, 0.1122897, 0.04864574,
  1.010497e-06, 0.0005027971, 0.08618055, 0.002259749, 0.05899917, 0.1188019, 
    0.1034012, 0.0387266, 0.05377733, 0.07954635, 0.003529967, 0.01241704, 
    0.001615428, 0.05370069, 0.08774656, 0.06782851, 0.0246198, 0.04178866, 
    0.141628, 0.0599447, 0.04900001, -7.709364e-05, -0.0002729801, 0.0831416, 
    0.04189777, 0.07191435, 0.06670643, 0.08770333, 0.005048909,
  7.789885e-06, 0.2494907, 0.2841289, 0.04374648, 0.06895426, 0.06971363, 
    0.06555171, 0.04431768, 0.1871502, 0.05172597, 0.04295694, 0.01979842, 
    0.1146298, 0.1280038, 0.04589471, 0.04331809, 0.05105508, 0.121981, 
    0.03533027, 0.008272535, 0.005609036, 0.01180864, 0.0001123309, 
    0.1643209, 0.1668345, 0.0330271, 0.04285652, 0.08264918, 6.641025e-05,
  0.01530837, 0.3152786, 0.2230299, 0.0025733, 0.002173802, 0.004119746, 
    0.009550978, 0.04389685, 0.2881958, 0.2276597, 0.09509762, 0.06246158, 
    0.1447213, 0.165062, 0.05674234, 0.001812844, 0.004309447, 0.02528549, 
    0.01519778, 0.0001965027, 0.01511609, 0.03969168, 0.1104012, 0.2550042, 
    0.1291321, 0.05431205, 0.0446587, 0.002932872, 0.003003729,
  0.01732357, 0.04067668, 1.793707e-05, 0.06865541, 0.003617184, 0.01648418, 
    0.06341369, 0.02791856, 0.01226874, 0.01701172, 0.006009909, 0.04797929, 
    0.1386548, 0.05969629, 0.06107516, 0.09685809, 0.08535659, 0.03593998, 
    0.04501829, 0.05533988, 0.1674022, 0.02582167, 0.001286615, 0.004506181, 
    0.0104111, 0.00107648, 0.02890278, 0.002336221, 0.1505505,
  0.09842233, 0.01517229, 0.001629991, 8.237454e-05, 0.06618955, 
    1.367403e-05, 0.01552145, 0.009288256, 0.05446412, 0.008384223, 
    0.01694812, 0.03323951, 0.0169922, 0.003845167, 0.02930504, 7.679508e-05, 
    0.008514006, 0.000337179, 0.0528274, 0.09652364, 0.1767561, 0.06448336, 
    0.01996402, 0.03606353, 0.01830602, 0.09895945, 0.0502103, 0.02579639, 
    0.07600754,
  0.03989042, 0.01841626, 0.01792692, 0.02689666, 0.05385248, 0.07807945, 
    0.03047588, -2.994636e-05, 0.001842005, 0.1795486, 0.192864, 0.1786359, 
    0.1576858, 0.1211913, 0.09890367, 0.09270546, 0.07643201, 0.04211597, 
    0.05971571, 0.03760227, 0.02381947, 0.08836593, 0.1652769, 0.1375333, 
    0.1629599, 0.1571065, 0.1075678, 0.03758495, 0.03155422,
  0.04115546, 0.02771335, 0.04329954, 0.01703591, 0.02404572, 0.0360855, 
    0.01263441, 0.009148861, 0.02825167, 0.0205577, 0.05177303, 0.09132789, 
    0.1045202, 0.196171, 0.2390827, 0.1787633, 0.2071408, 0.2471264, 
    0.2234525, 0.01220385, 0.004395306, 0.04125144, 0.06817549, 0.1749986, 
    0.129806, 0.1379457, 0.1186962, 0.06553892, 0.05341752,
  0.02195252, 0.01604651, 0.001174946, 0.004856516, 0.000686656, 1.28449e-05, 
    -4.732012e-07, 0, 0, 0, 0.0004171191, 0.0001290648, 0.01268619, 
    0.01504511, 0.02136992, 0.02360737, 0.02412076, 0.03983587, 0.02918181, 
    0.006743069, 0.008666952, 0.009428595, 0.007867798, 0.07645985, 
    0.06778077, 0.06068353, 0.08858177, 0.07692217, 0.04039134,
  0.01925012, 0.007210007, 0.01517789, 0.001283132, 0.0002530008, 
    0.003531924, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0002863194, 
    -8.916531e-06, 0, 0, 0, -2.079869e-06, 0.001774194, 0.01966416, 
    0.004296916, 0.002315706, 0.006560824, 0.0163194,
  4.567989e-05, -6.605145e-05, -4.114518e-06, 0.000459246, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002374171,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.311202e-06, 
    -0.0001396749, 0.0003545429, -6.766642e-07, -1.27896e-05, -8.794742e-06, 
    5.729943e-06, -4.448487e-05, -3.231514e-06, -8.061807e-07, -5.227864e-07, 
    0, 0,
  0, 0, 0, 0, -1.595747e-05, 0, 9.215563e-09, 0, 0, 0, -1.160608e-08, 0, 
    -0.0002707554, 0.005024718, 0.002864863, -6.428599e-05, -0.0001341509, 
    0.03288633, 0.06333212, 0.07341347, 0.05817549, 0.02078957, 0.0187989, 
    0.006423049, 0.004510644, 0.0003508849, -2.064947e-06, 0, 0,
  0.03611628, 0.01876456, 0.00136014, 0.02730013, 0.03972976, 0.03875021, 
    0.04813337, 0.03494369, 0.03054223, 0.03693947, 0.06867515, 0.08467495, 
    0.04362964, 0.04389693, 0.07225443, 0.08323267, 0.1382303, 0.1088896, 
    0.1146662, 0.09905224, 0.147925, 0.06790175, 0.03115237, 0.05807327, 
    0.04768776, 0.02124416, 0.008722787, 0.01005127, 0.0384407,
  0.1355065, 0.1460051, 0.2052535, 0.1279671, 0.1563602, 0.222242, 0.1787378, 
    0.1699736, 0.09471903, 0.1035725, 0.1202568, 0.1483977, 0.1665299, 
    0.1590039, 0.1279585, 0.1677246, 0.197085, 0.1232455, 0.1071435, 
    0.1106473, 0.1541775, 0.1657853, 0.1765476, 0.07228559, 0.08470254, 
    0.07380424, 0.07750608, 0.2006657, 0.1694553,
  0.1217493, 0.1139914, 0.07940017, 0.1200015, 0.1681575, 0.07120718, 
    0.06686123, 0.07248102, 0.06907017, 0.1368748, 0.1546963, 0.1200874, 
    0.06490356, 0.0880352, 0.09980612, 0.09575661, 0.1634813, 0.1827786, 
    0.1680653, 0.1705539, 0.2545077, 0.1278756, 0.1115185, 0.1318833, 
    0.1863219, 0.2042446, 0.1436833, 0.168909, 0.1778233,
  0.02229544, 0.01223453, 0.07884476, 0.05964552, 0.02541742, 0.09544592, 
    0.1253429, 0.0567295, 0.03527912, 0.1256563, 0.213541, 0.1173364, 
    0.1209881, 0.07570392, 0.07475209, 0.09275582, 0.1083886, 0.1093348, 
    0.1630837, 0.1242509, 0.1064489, 0.03503331, 0.02545113, 0.009345091, 
    0.01908442, 0.09153695, 0.1092392, 0.1085486, 0.03270703,
  1.107419e-06, 0.0006902271, 0.04222292, 0.002095039, 0.0425272, 0.1267859, 
    0.1013804, 0.0315693, 0.05303867, 0.08663005, 0.001487104, 0.01565413, 
    -0.0002135257, 0.04014939, 0.07924883, 0.04926459, 0.02169299, 
    0.04127887, 0.1404125, 0.05463491, 0.01423974, 1.709999e-06, 
    -0.0001726529, 0.07686382, 0.04592704, 0.06776831, 0.03091061, 
    0.04926754, 6.519116e-05,
  2.319142e-06, 0.2538199, 0.2357048, 0.03811988, 0.07610226, 0.04497359, 
    0.05897958, 0.03523614, 0.1642257, 0.04458527, 0.04069681, 0.02148131, 
    0.1131141, 0.1048706, 0.03633981, 0.04475532, 0.03635826, 0.09214444, 
    0.01432014, 0.004496902, 0.002548506, 0.0005333182, 4.547614e-05, 
    0.1385544, 0.1447399, 0.02374408, 0.04264138, 0.04345066, 6.409036e-05,
  0.01180603, 0.2749378, 0.1816339, 0.007399517, 0.001510293, 0.005249072, 
    0.008519113, 0.02983623, 0.189728, 0.2029517, 0.0864682, 0.04446571, 
    0.1112152, 0.161672, 0.05336007, 0.002856186, 0.00549431, 0.02549351, 
    0.004699988, 0.0004723771, 0.01304205, 0.02810544, 0.1374187, 0.2179756, 
    0.09762459, 0.06426511, 0.02723486, 0.002983107, 0.005042689,
  0.003719195, 0.02403886, 1.095008e-05, 0.04741058, 0.002071158, 0.01038515, 
    0.04107728, 0.02332523, 0.008035023, 0.01541472, 0.008499878, 0.04337505, 
    0.1084538, 0.04938726, 0.06749205, 0.1066359, 0.07197148, 0.03777445, 
    0.03351251, 0.04654302, 0.1557689, 0.02101604, 0.001295877, 0.001415148, 
    0.001264283, 0.004604963, 0.01257596, 0.0002819074, 0.1111028,
  0.06197187, 0.004925722, 0.0006382095, 8.582494e-05, 0.05258115, 
    2.69421e-06, 0.01647396, 0.002789686, 0.05458158, 0.003696907, 
    0.009064866, 0.02993969, 0.02004008, 0.0004188649, 0.02635621, 
    0.001637457, 0.006012368, 1.152091e-05, 0.02654089, 0.09078582, 
    0.1645333, 0.05832301, 0.01055396, 0.02220284, 0.01972352, 0.08503095, 
    0.02309484, 0.01925669, 0.08005348,
  0.05270828, 0.04613548, 0.03928756, 0.03774385, 0.06154565, 0.07202919, 
    0.03634046, 0.003102193, 0.009382775, 0.1811824, 0.1747519, 0.1530303, 
    0.163629, 0.1110258, 0.08308116, 0.09240545, 0.05969194, 0.02825431, 
    0.03915935, 0.03470953, 0.03191648, 0.07162462, 0.1297212, 0.1283265, 
    0.1321437, 0.1541659, 0.07779264, 0.03696739, 0.0685651,
  0.1021367, 0.09941453, 0.1306536, 0.05061199, 0.08289492, 0.05615454, 
    0.02695448, 0.1525915, 0.1242542, 0.04030295, 0.1035883, 0.1250265, 
    0.1213655, 0.2074441, 0.2435682, 0.1764954, 0.1990534, 0.2503373, 
    0.2477629, 0.08587891, 0.02066156, 0.1253508, 0.1346042, 0.1652352, 
    0.1811988, 0.1869066, 0.1340206, 0.101055, 0.06941336,
  0.1019948, 0.07302976, 0.03925879, 0.04886421, 0.03164053, 0.01546801, 
    0.0009806727, 0, 0, -2.548166e-05, 0.003254166, 0.009202916, 0.01207966, 
    0.01541561, 0.03553082, 0.03094463, 0.0733704, 0.06923154, 0.1227121, 
    0.02963385, 0.03662648, 0.04356386, 0.02082042, 0.1078867, 0.1253106, 
    0.1115103, 0.1659265, 0.1309987, 0.08639254,
  0.06335886, 0.05377612, 0.05499285, 0.05281227, 0.02762995, 0.0178323, 
    0.01312269, 5.111111e-09, 0, 0, 0, 0, 0, 0, -7.744102e-05, 0.01073882, 
    -0.0001074484, 0.0324798, -9.63516e-06, 0.0007838184, -0.0004388343, 
    2.257717e-07, 0.0001382846, 0.06935578, 0.1247812, 0.02458827, 
    0.00189545, 0.01735602, 0.06047125,
  0.0256716, 0.05533892, 0.03009331, 0.05185953, 0.01816211, 0.02048291, 
    0.01637365, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.383482e-05, -8.716694e-06, 
    -1.043963e-05, -3.908834e-05, 2.419032e-05, -0.0008240728, -0.002106707, 
    0.03325609, 0, 0, 0.001443966, 0.02801158,
  0, 0, -4.253982e-11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, -9.246099e-08, -3.603001e-08, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0001206291, 0.003950194, 
    0.01316164, 0.004255193, 0.00627416, 0.0004533771, -7.632027e-05, 
    -5.061112e-05, 0.001179868, 0.006580589, 0.003167791, -0.002395712, 
    0.008442172, 0, 0,
  7.935386e-05, 0.0009484792, -0.0001220556, 0.005153832, 8.844228e-05, 
    -8.850358e-06, 0.001140076, -4.785915e-06, -8.28817e-08, 0.000166053, 
    0.001833452, -1.318667e-06, -0.0009234486, 0.01071377, 0.02245086, 
    0.0193318, 0.02127126, 0.07831328, 0.1418391, 0.1649166, 0.137053, 
    0.08903947, 0.05245544, 0.02333857, 0.04038443, 0.01673592, 0.01088956, 
    -0.0002893795, 0,
  0.08565338, 0.05347877, 0.03435596, 0.0749073, 0.07594915, 0.06083776, 
    0.08706024, 0.07227115, 0.07744645, 0.1265727, 0.1648158, 0.1950828, 
    0.1257367, 0.1281507, 0.1660874, 0.1953736, 0.2194673, 0.1424721, 
    0.1962248, 0.1606744, 0.2148118, 0.1613669, 0.125607, 0.1811495, 
    0.1206751, 0.06093396, 0.06236417, 0.0667641, 0.08529636,
  0.1628344, 0.174651, 0.2227917, 0.1498276, 0.1638797, 0.2274525, 0.1791732, 
    0.1831102, 0.1171443, 0.1332256, 0.1812695, 0.2200674, 0.1956893, 
    0.1729748, 0.1468045, 0.1876242, 0.1960485, 0.1225067, 0.1276261, 
    0.1378182, 0.184481, 0.161874, 0.1607897, 0.1542407, 0.1393055, 0.127305, 
    0.1090615, 0.2223334, 0.1971709,
  0.1065354, 0.09515365, 0.06208367, 0.1163953, 0.1512187, 0.05491192, 
    0.06342757, 0.06773695, 0.06729255, 0.1326281, 0.1518545, 0.1087031, 
    0.05406678, 0.07905479, 0.09158679, 0.08776209, 0.1606504, 0.1842285, 
    0.160068, 0.1704912, 0.2488384, 0.1039603, 0.1148832, 0.1512683, 
    0.1635142, 0.1862818, 0.1548392, 0.1580894, 0.1775115,
  0.01064922, 0.001130723, 0.05791263, 0.04920309, 0.01792535, 0.07151926, 
    0.1221075, 0.02669533, 0.04613429, 0.1074317, 0.2206106, 0.1110082, 
    0.08183284, 0.05122328, 0.08450813, 0.0856492, 0.08900848, 0.1071853, 
    0.135542, 0.1134318, 0.1097738, 0.02565182, 0.03229463, 0.01213455, 
    0.01935355, 0.08748484, 0.1023283, 0.08662131, 0.03801982,
  4.931836e-07, 0.0006796688, 0.01742143, 0.001497457, 0.0313371, 0.1316416, 
    0.108289, 0.03156076, 0.05117603, 0.08512788, 0.0009320377, 0.0129287, 
    7.877767e-05, 0.03979045, 0.07124366, 0.036313, 0.03290274, 0.04912642, 
    0.1283238, 0.04410655, 0.00279719, 3.781321e-06, -4.190794e-05, 
    0.05832691, 0.04164761, 0.06907216, 0.02051926, 0.01854891, 1.592408e-05,
  5.077979e-06, 0.2312545, 0.1963001, 0.03883602, 0.07120955, 0.02570029, 
    0.06211656, 0.03429944, 0.1293449, 0.0326763, 0.0403473, 0.01991778, 
    0.1104732, 0.0788216, 0.02664164, 0.04168847, 0.02622041, 0.05636244, 
    0.01040445, 0.003494704, 0.002256317, -0.0002626565, 6.544517e-05, 
    0.09881459, 0.1257583, 0.02274588, 0.03730543, 0.01351331, 1.80999e-05,
  0.008084041, 0.2366886, 0.1375783, 0.008653327, 0.002454271, 0.006359777, 
    0.008693783, 0.01705547, 0.1175047, 0.1726363, 0.08403444, 0.02941953, 
    0.07604083, 0.1462291, 0.05016917, 0.003332794, 0.005546263, 0.02221655, 
    0.003423275, 0.0009138405, 0.01199759, 0.01588527, 0.1323017, 0.1862639, 
    0.07123343, 0.07118052, 0.01819999, 0.002376687, 0.0125965,
  0.001096744, 0.01462584, 3.629735e-05, 0.03203728, 0.001588548, 
    0.006971323, 0.0271606, 0.01693484, 0.006682744, 0.01135314, 0.00707175, 
    0.04328013, 0.07209682, 0.04234354, 0.07700048, 0.1098199, 0.05509427, 
    0.04278306, 0.0162065, 0.02517211, 0.1353336, 0.01629021, 0.0005946183, 
    0.0007773875, 0.0002270206, 0.00122795, 0.007231014, 0.002267012, 
    0.08047599,
  0.02909062, 0.003079843, -4.649625e-06, 3.290678e-05, 0.04777148, 
    9.178038e-08, 0.008424497, 0.001073086, 0.04309976, 0.00226613, 
    0.003253574, 0.02659276, 0.03147386, 2.53495e-05, 0.01829014, 
    5.938036e-05, 0.002695287, 3.332011e-06, 0.03012891, 0.04859428, 0.15015, 
    0.05451415, 0.01022826, 0.01447438, 0.01407223, 0.05093495, 0.008160813, 
    0.01760176, 0.07880168,
  0.05841959, 0.05724794, 0.03283212, 0.02485869, 0.06086697, 0.06552582, 
    0.03740977, 0.005313685, 0.03169239, 0.1713913, 0.155847, 0.1303376, 
    0.1590581, 0.100529, 0.07185839, 0.08657008, 0.04517674, 0.01975105, 
    0.02934917, 0.02834586, 0.02405436, 0.05793022, 0.1198977, 0.1145497, 
    0.1152081, 0.1455992, 0.0662158, 0.0311683, 0.05060454,
  0.1057389, 0.111792, 0.190709, 0.1200107, 0.09203216, 0.06578799, 
    0.05357125, 0.2699169, 0.2179288, 0.09845059, 0.120386, 0.1167962, 
    0.1283074, 0.2139481, 0.2657317, 0.1602596, 0.1839416, 0.2378193, 
    0.2036941, 0.1481619, 0.05600727, 0.1811895, 0.1369972, 0.1456342, 
    0.1719661, 0.1851387, 0.1309842, 0.09730349, 0.05784452,
  0.1524023, 0.2091855, 0.1040354, 0.1532029, 0.04002731, 0.04758519, 
    0.03749893, -0.0001943191, -0.0001466369, 0.02416968, 0.04830913, 
    0.01606216, 0.01406168, 0.0303264, 0.08582771, 0.04564684, 0.1081743, 
    0.09509924, 0.2471102, 0.05851909, 0.1216715, 0.1119837, 0.1219819, 
    0.131633, 0.1278294, 0.1237153, 0.1840914, 0.1453012, 0.08232655,
  0.1898466, 0.1343232, 0.1905295, 0.1687784, 0.1149565, 0.08766627, 
    0.03205577, 0.02386392, 0.0008707992, -2.437574e-05, -1.100346e-07, 0, 
    -0.0007769963, 0.00183748, 0.02365914, 0.02652926, 0.02100458, 
    0.08561613, 0.0422851, 0.04090695, 0.05610493, 0.01938669, 0.05769816, 
    0.1182677, 0.1735721, 0.08294754, 0.006726562, 0.06981792, 0.1299546,
  0.08393186, 0.1345915, 0.08906561, 0.1454244, 0.1757784, 0.1006773, 
    0.02637232, 0.04394453, 0.01696778, -1.835481e-05, -5.001029e-06, 0, 0, 
    0, 0, 0.01224641, 0.0272269, 0.04548594, 0.04678377, 0.03891537, 
    0.06430665, 0.02829021, 0.04659965, 0.02300069, 0.04753284, 
    -0.0001314797, -1.631462e-06, 0.03708703, 0.07525535,
  0, 0.003703641, -0.0001252954, 0.002732932, 0.01916928, 0.02225086, 
    0.02112216, 0.01944596, 0.01148639, 0.004817366, 0.0003456301, 
    0.001139911, -4.740639e-05, 0, 0, 0, 9.132791e-07, 1.113344e-06, 
    -2.386146e-05, 0.01726156, 0.03917188, 0.03828497, -9.568497e-05, 
    -0.002147914, 0.0001018584, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0020066, 0.03957583, 0.04244142, 
    0.03714195, 0.01979265, 0.01934662, 0.007346662, 0.005989891, 
    0.0005997736, 0.009343283, 0.04876777, 0.05170619, 0.03014055, 
    0.03093502, 0.002161291, 0,
  0.02597301, 0.03205172, 0.03530956, 0.03192549, 0.000854363, 0.003099018, 
    0.01550176, -0.0001019659, -0.0006759431, 0.002852105, 0.002037584, 
    -9.275212e-05, -0.0002579843, 0.04668403, 0.04920987, 0.05223136, 
    0.08191186, 0.154001, 0.2014631, 0.2462851, 0.2593814, 0.262412, 
    0.2666046, 0.147134, 0.1292077, 0.04618509, 0.0433162, 0.01457885, 
    0.03045382,
  0.1399646, 0.1088933, 0.08390012, 0.1893141, 0.1365895, 0.1156705, 
    0.1341355, 0.1498563, 0.1391553, 0.2074476, 0.2402942, 0.2249115, 
    0.1706714, 0.1832691, 0.2193422, 0.259117, 0.2329959, 0.1582004, 
    0.2176782, 0.1879963, 0.2641523, 0.1805868, 0.2011418, 0.2308591, 
    0.1838208, 0.1929708, 0.1496913, 0.1145527, 0.1172639,
  0.1597999, 0.1853178, 0.2250192, 0.1631836, 0.1704724, 0.2055422, 
    0.1677256, 0.1663836, 0.1121587, 0.1421884, 0.1999491, 0.2191636, 
    0.1935558, 0.17411, 0.128108, 0.1693947, 0.1784941, 0.113961, 0.137207, 
    0.1755855, 0.193995, 0.1726401, 0.1501799, 0.1797779, 0.1547838, 
    0.1679302, 0.1796456, 0.2329278, 0.1951944,
  0.09755161, 0.07624517, 0.04881097, 0.1026512, 0.1269869, 0.04577361, 
    0.06020996, 0.05526699, 0.0652162, 0.1288184, 0.150127, 0.08669934, 
    0.04752139, 0.07445722, 0.08215749, 0.09219871, 0.1633205, 0.1780789, 
    0.1382167, 0.1755088, 0.2512147, 0.09584243, 0.1316583, 0.1586547, 
    0.1358259, 0.1794768, 0.1710782, 0.1425662, 0.1741755,
  0.01206621, -4.156143e-05, 0.04028557, 0.04550362, 0.01489777, 0.05325134, 
    0.08460283, 0.01055709, 0.04055932, 0.1027663, 0.2111211, 0.09323302, 
    0.05006213, 0.04780788, 0.08361997, 0.09168694, 0.07317407, 0.09005808, 
    0.1182063, 0.08231118, 0.10203, 0.02272859, 0.02747731, 0.006936314, 
    0.02854005, 0.08113142, 0.08654805, 0.06867995, 0.03617245,
  1.194624e-07, 0.0006412497, 0.003499137, 0.001039514, 0.02226827, 
    0.1203806, 0.106686, 0.02395158, 0.05238351, 0.0575955, 0.0008933598, 
    0.01031063, -6.978041e-05, 0.04261042, 0.04671702, 0.02388633, 
    0.02791088, 0.05258192, 0.09758905, 0.03980606, 0.0001677619, 
    3.022032e-06, 1.321453e-06, 0.04850001, 0.03720254, 0.06847897, 
    0.01331216, 0.003369284, 2.368699e-06,
  2.021293e-06, 0.2296152, 0.1728913, 0.06151669, 0.06504489, 0.01759498, 
    0.04693424, 0.03312565, 0.1129754, 0.02355615, 0.03721687, 0.01889102, 
    0.1125798, 0.06363808, 0.01919425, 0.02376218, 0.02477096, 0.03492287, 
    0.008982595, 0.002462103, 0.001154205, 0.0002245616, 2.372469e-05, 
    0.07335582, 0.1188383, 0.02206193, 0.04202453, 0.003862753, 1.330208e-05,
  0.005879792, 0.1911064, 0.1260986, 0.004074308, 0.00270236, 0.005349573, 
    0.005672744, 0.0144629, 0.08140229, 0.1715064, 0.07701232, 0.01840444, 
    0.04937843, 0.1391128, 0.05036704, 0.005055569, 0.004266135, 0.015795, 
    0.008642601, 0.0009512822, 0.01823886, 0.01493017, 0.1317115, 0.1609771, 
    0.06987713, 0.06990673, 0.0142831, 0.002627937, 0.01031972,
  0.001422965, 0.00124082, 0.0001324712, 0.02934314, 0.00143537, 0.005201736, 
    0.01704399, 0.01108943, 0.004958147, 0.008349305, 0.004919337, 
    0.05487864, 0.05200054, 0.05261798, 0.08783627, 0.1114095, 0.03814905, 
    0.03589189, 0.01014738, 0.02237481, 0.1225637, 0.01778639, 0.0001912766, 
    0.000537517, 0.0007050254, -1.870148e-06, 0.001769479, 0.009480172, 
    0.06242209,
  0.01802891, 0.0002374194, -1.266286e-05, 1.80585e-05, 0.04668472, 
    -5.770936e-07, 0.004013612, 0.0008312584, 0.02100444, 0.003890506, 
    0.001652096, 0.02622559, 0.01237182, 4.62748e-05, 0.008814366, 
    5.163747e-05, 0.001140456, 6.052732e-06, 0.01253496, 0.0154628, 
    0.1136416, 0.05024808, 0.006657877, 0.0108165, 0.0277102, 0.02480739, 
    0.000539359, 0.02669199, 0.04477622,
  0.05194316, 0.05820745, 0.02743204, 0.01811923, 0.06189635, 0.05772383, 
    0.04332886, 0.008618508, 0.06183454, 0.1500361, 0.1379321, 0.1252197, 
    0.1569501, 0.09361443, 0.05244274, 0.05169481, 0.01299267, 0.005811787, 
    0.02619918, 0.0219193, 0.02496568, 0.04315539, 0.1032002, 0.1058026, 
    0.09932537, 0.1247417, 0.0507515, 0.0311339, 0.03032385,
  0.0960309, 0.1022774, 0.1826009, 0.1403978, 0.08678024, 0.0837266, 
    0.1083833, 0.240873, 0.1968881, 0.1023605, 0.1247771, 0.1439835, 
    0.1305753, 0.2240399, 0.2835672, 0.16791, 0.1621038, 0.2241476, 
    0.1588177, 0.1462338, 0.1367313, 0.1857421, 0.134314, 0.1299972, 
    0.1595604, 0.1865432, 0.1310513, 0.08753407, 0.04212805,
  0.1732511, 0.2358079, 0.110934, 0.1381308, 0.02533734, 0.08105724, 
    0.1149757, 0.01628123, 0.02168869, 0.05459712, 0.09558977, 0.07140415, 
    0.1075147, 0.1200324, 0.1219004, 0.114448, 0.1528639, 0.1735506, 
    0.2720696, 0.1741658, 0.134922, 0.1230605, 0.1478287, 0.2245194, 
    0.1655426, 0.1259496, 0.1784755, 0.1603868, 0.1048559,
  0.2487921, 0.1948408, 0.2129747, 0.139568, 0.1240993, 0.12006, 0.09582788, 
    0.09607344, 0.09973302, 0.03041063, 0.02211737, 9.316559e-05, 0.0386055, 
    0.001268076, 0.01990674, 0.04478711, 0.0703166, 0.1540172, 0.103747, 
    0.09532461, 0.0954238, 0.1105592, 0.1206688, 0.1729766, 0.2013788, 
    0.09465835, 0.080577, 0.1702872, 0.2057771,
  0.1291793, 0.1947027, 0.1875201, 0.1877473, 0.2188912, 0.1734731, 
    0.09368705, 0.09566218, 0.09815811, 0.07433172, 0.0006667956, 0.01456415, 
    0.01102166, 0.0339619, 0.0753049, 0.09602011, 0.1239827, 0.07938848, 
    0.06060593, 0.1281453, 0.1603305, 0.0967, 0.1020446, 0.01674881, 
    0.07377283, 0.0003637328, 1.253167e-05, 0.1046612, 0.1003025,
  0.0003706317, 0.03683271, 0.1053633, 0.09736158, 0.09944186, 0.1259782, 
    0.1894891, 0.1968628, 0.1155558, 0.0561482, 0.07579518, 0.05819933, 
    0.02067478, 0.01966259, 0.01621029, 0.01057729, 0.009200287, 0.005133405, 
    0.03686086, 0.07993252, 0.07963457, 0.07150414, 0.02816295, 0.02707639, 
    0.00967097, -5.92645e-05, 0, 0, -0.0001570287,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.02379001, 0.05218612, 0.04934406, 
    0.05822233, 0.0477334, 0.04351093, 0.0148972, 0.01138476, 0.01066357, 
    0.05106927, 0.1812757, 0.1910079, 0.09734631, 0.08651949, 0.0159271, 
    0.0003125692,
  0.1155613, 0.120048, 0.1419488, 0.08984014, 0.001085354, 0.004986844, 
    0.04261287, -0.0008686026, -0.001364391, 0.02131876, 0.002081494, 
    -0.000476323, 0.0292218, 0.1412641, 0.1563046, 0.1197374, 0.1457102, 
    0.218867, 0.2357794, 0.2673164, 0.2790618, 0.2836197, 0.3255187, 
    0.2249811, 0.214183, 0.1590271, 0.1886215, 0.1589569, 0.05841611,
  0.2000004, 0.1650766, 0.1659757, 0.2579536, 0.1778067, 0.165694, 0.1773009, 
    0.2306566, 0.1739338, 0.2548603, 0.2578076, 0.2247399, 0.2126167, 
    0.2053607, 0.2509052, 0.2630011, 0.2489902, 0.1560666, 0.2221969, 
    0.2027944, 0.2822653, 0.2279869, 0.2441394, 0.2437254, 0.2275199, 
    0.2454462, 0.2108006, 0.2007495, 0.2120646,
  0.1598031, 0.1706063, 0.2327791, 0.172054, 0.1755334, 0.2167074, 0.1850123, 
    0.1770287, 0.1216675, 0.1676422, 0.2128666, 0.1933427, 0.1933382, 
    0.176354, 0.1269359, 0.1515026, 0.1940927, 0.1106262, 0.1598133, 
    0.1969393, 0.1913882, 0.1630864, 0.1527828, 0.1999206, 0.2230027, 
    0.2009485, 0.1925942, 0.2273504, 0.1979235,
  0.09836044, 0.07011889, 0.05405445, 0.09350446, 0.1082975, 0.04306141, 
    0.06739058, 0.05655173, 0.05474421, 0.1270416, 0.1379005, 0.07391201, 
    0.04377278, 0.06586409, 0.07791575, 0.1104108, 0.1482583, 0.1750346, 
    0.1379032, 0.1784014, 0.2610675, 0.09558181, 0.1349044, 0.1605842, 
    0.09638503, 0.1663271, 0.1673623, 0.1171121, 0.1564504,
  0.002815957, 0.0001892459, 0.03169028, 0.0427679, 0.01337398, 0.0451608, 
    0.05246379, 0.001130976, 0.03498931, 0.0903093, 0.1986936, 0.08410867, 
    0.03510427, 0.05022955, 0.07025155, 0.09191741, 0.05103841, 0.07156591, 
    0.1060754, 0.06095469, 0.1110036, 0.02262507, 0.02040276, 0.008141261, 
    0.03506352, 0.0787847, 0.07497031, 0.0532605, 0.03132263,
  7.315747e-08, 0.0007242036, 0.002136121, 0.0008558473, 0.01761737, 
    0.1167124, 0.1054939, 0.01935191, 0.05663903, 0.03912801, 0.0003780501, 
    0.007591708, 0.0003359059, 0.03707076, 0.03294663, 0.01695607, 
    0.02066563, 0.06503353, 0.07721549, 0.02790801, 2.519701e-05, 
    1.49988e-06, 6.751223e-08, 0.02591377, 0.02886527, 0.05543627, 
    0.008120777, 0.0003868539, 2.065126e-06,
  6.299165e-06, 0.2324302, 0.1688661, 0.07696797, 0.04703833, 0.01363387, 
    0.04754593, 0.0375142, 0.1099273, 0.02193086, 0.04122558, 0.02357811, 
    0.1241683, 0.05631903, 0.01444257, 0.01588888, 0.02968775, 0.03459152, 
    0.01174653, 0.001812666, 0.0008434334, -1.097193e-05, 0.0002422589, 
    0.05134675, 0.1192267, 0.0158576, 0.04431634, 0.002503951, 2.450557e-06,
  0.01096701, 0.1621311, 0.09605677, 0.008050212, 0.004014159, 0.004429172, 
    0.006928739, 0.01210795, 0.06947622, 0.1833307, 0.09729966, 0.01344582, 
    0.04819335, 0.1299578, 0.04809479, 0.01127117, 0.004029452, 0.00878852, 
    0.01155698, 0.001047585, 0.03681767, 0.02923127, 0.1363734, 0.1628081, 
    0.06772208, 0.07193132, 0.01335188, 0.004254734, 0.01060812,
  0.002015297, 0.0001227699, 0.0001283901, 0.0322037, 0.001186295, 
    0.004464721, 0.0138823, 0.006812281, 0.0042152, 0.006646438, 0.005557979, 
    0.04625701, 0.03672716, 0.04022724, 0.09620295, 0.09543419, 0.03599831, 
    0.01773612, 0.008346207, 0.02479007, 0.114523, 0.0121825, 0.0001880219, 
    0.0006220831, 0.001345769, 5.319728e-06, -0.0001148596, 0.04499607, 
    0.05522734,
  0.01287345, -2.159878e-05, -1.053571e-05, 3.979149e-05, 0.04430408, 
    -9.13031e-05, 0.001861046, 0.0006055536, 0.0109346, 0.00664937, 
    0.001656065, 0.02690213, 0.01410548, 0.000102772, 0.0005017831, 
    0.0004083678, 3.574916e-05, 2.137859e-06, 0.006902885, 0.0003738951, 
    0.06856814, 0.04837823, 0.00323385, 0.005791737, 0.01044177, 0.004708597, 
    -0.0006330611, 0.02204513, 0.01639426,
  0.04321469, 0.06171906, 0.03564755, 0.02201004, 0.07058623, 0.04457215, 
    0.04759326, 0.01304736, 0.08962731, 0.1406158, 0.1301915, 0.1124495, 
    0.1566088, 0.1016003, 0.03466477, 0.02543241, 0.0005061475, 0.001610819, 
    0.01505041, 0.02115519, 0.02197997, 0.03740683, 0.09470785, 0.08741377, 
    0.0869273, 0.08853817, 0.03907428, 0.02550374, 0.01381931,
  0.09194108, 0.1006534, 0.1821306, 0.1372186, 0.08391839, 0.1007897, 
    0.1847422, 0.1930894, 0.1685388, 0.1027717, 0.1266565, 0.1560601, 
    0.1194803, 0.2123542, 0.2887737, 0.1647833, 0.1626849, 0.1886609, 
    0.1295806, 0.14081, 0.1818242, 0.1788246, 0.1360362, 0.1253693, 
    0.1559439, 0.1590734, 0.1127218, 0.06960294, 0.03403013,
  0.1877575, 0.2310203, 0.1044469, 0.1294493, 0.0195368, 0.08527581, 
    0.1329605, 0.05276978, 0.06733479, 0.1112982, 0.1642206, 0.12048, 
    0.122361, 0.1425346, 0.1496527, 0.1539545, 0.1822942, 0.232499, 
    0.2644965, 0.1602598, 0.1394896, 0.1363177, 0.1527794, 0.2498413, 
    0.1827458, 0.1373381, 0.1640869, 0.1551938, 0.1458137,
  0.2796996, 0.2161187, 0.195035, 0.1322335, 0.1200203, 0.1468019, 0.1342309, 
    0.1463629, 0.1827319, 0.1348571, 0.1132971, 0.005667232, 0.07526319, 
    0.08197721, 0.01099254, 0.117764, 0.1273514, 0.2205312, 0.1121635, 
    0.08482216, 0.1383177, 0.1374844, 0.1213811, 0.189447, 0.1958618, 
    0.1328072, 0.06914357, 0.2018794, 0.2398206,
  0.1927703, 0.2599691, 0.2505173, 0.2074703, 0.2036749, 0.1856714, 
    0.1375612, 0.1290382, 0.1544898, 0.2691458, 0.05024781, 0.04194221, 
    0.03216159, 0.07408816, 0.1086186, 0.1723183, 0.1376044, 0.09174106, 
    0.06853876, 0.1307647, 0.1867791, 0.1607981, 0.1255943, 0.02453891, 
    0.05633871, 0.0001053625, -0.0001144033, 0.1449671, 0.1459176,
  0.09493648, 0.1442491, 0.1979941, 0.1806786, 0.1661572, 0.1759304, 
    0.2249842, 0.2140222, 0.1381408, 0.125271, 0.1490942, 0.1257714, 
    0.09164786, 0.09223723, 0.1222261, 0.06970726, 0.02867088, 0.07101004, 
    0.1066101, 0.1199577, 0.1335534, 0.1388904, 0.0843632, 0.03871873, 
    0.02621183, -0.0002319669, -0.0001249026, -0.001356168, 0.1113066,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.192887e-05, -2.192887e-05, 
    -2.192887e-05, -2.192887e-05, -2.192887e-05, -2.192887e-05, 
    -2.192887e-05, 0, 0, 0, 0, 0, 0, 0, 0,
  -0.0006693949, -7.566133e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0004582497, 
    0.05446088, 0.1260816, 0.1160819, 0.1526408, 0.1063471, 0.1150668, 
    0.05770069, 0.03270929, 0.02651222, 0.1070064, 0.2393116, 0.3117779, 
    0.2890614, 0.241807, 0.04183084, 0.005077882,
  0.1832468, 0.2472305, 0.2105217, 0.1763365, 0.01694132, 0.02812632, 
    0.1236013, -0.004725508, 0.0138695, 0.05141968, 0.02502978, -0.001638532, 
    0.08940328, 0.2275151, 0.249534, 0.2365257, 0.2054436, 0.2614269, 
    0.2700174, 0.2822252, 0.2807116, 0.285495, 0.3270958, 0.2438782, 
    0.2724729, 0.1724633, 0.1738098, 0.1775727, 0.1266137,
  0.2607745, 0.2482238, 0.2585173, 0.3221052, 0.239332, 0.2396914, 0.2110645, 
    0.3019959, 0.2341335, 0.2922634, 0.2966599, 0.2456214, 0.2079167, 
    0.2313288, 0.24981, 0.2727372, 0.2629797, 0.166519, 0.1997793, 0.2014765, 
    0.2777848, 0.2483106, 0.2306386, 0.2379654, 0.2549156, 0.2154811, 
    0.193126, 0.1990696, 0.2312049,
  0.1584485, 0.1735714, 0.237927, 0.1794414, 0.1746928, 0.2219294, 0.1791373, 
    0.192267, 0.1223504, 0.18603, 0.2101758, 0.1842437, 0.1859833, 0.1627706, 
    0.1159339, 0.1304756, 0.2087666, 0.09903155, 0.1779044, 0.1778381, 
    0.185407, 0.1803588, 0.1527442, 0.2329528, 0.2042227, 0.2134506, 
    0.2069343, 0.225728, 0.2089218,
  0.09295342, 0.0550711, 0.05721813, 0.09307986, 0.1042984, 0.04135438, 
    0.06476669, 0.03990794, 0.05925997, 0.1105844, 0.09689606, 0.04741885, 
    0.04131949, 0.07057426, 0.07646828, 0.09571299, 0.1373694, 0.1650413, 
    0.1484215, 0.1737911, 0.2286222, 0.08626992, 0.1419667, 0.1356126, 
    0.06397648, 0.1645994, 0.157347, 0.1091852, 0.1487421,
  0.001286092, 0.0001124725, 0.02970433, 0.04200844, 0.01102236, 0.0384589, 
    0.02758703, 0.0007642391, 0.03808314, 0.08836669, 0.1732338, 0.0730442, 
    0.02446044, 0.05123484, 0.05959282, 0.08930124, 0.04149946, 0.05956031, 
    0.1045973, 0.0487753, 0.1047049, 0.02888752, 0.01419512, 0.009516127, 
    0.03734128, 0.07352126, 0.08062572, 0.04552848, 0.02422095,
  2.345783e-07, 0.0006974985, 0.0008379482, 0.0007917614, 0.01482208, 
    0.1101433, 0.105574, 0.02152558, 0.06110144, 0.022337, 0.0004314828, 
    0.003932978, -0.0005569623, 0.04165953, 0.02680776, 0.01382653, 
    0.0291984, 0.06718445, 0.0721209, 0.01555808, 1.668339e-05, 4.23088e-07, 
    4.356071e-08, 0.01140974, 0.02310565, 0.04374636, 0.004166162, 
    0.0001891569, 4.643346e-07,
  0.0003682651, 0.2462779, 0.1789754, 0.08224647, 0.04980882, 0.01210152, 
    0.05746617, 0.03475376, 0.1101509, 0.01866971, 0.03658823, 0.03101193, 
    0.1250281, 0.06145044, 0.01196419, 0.01185102, 0.03499112, 0.03556225, 
    0.01101399, 0.001327838, 0.001456451, 0.0002766732, 0.001810576, 
    0.04073385, 0.129599, 0.01128117, 0.05333636, 0.001969357, -1.173896e-06,
  0.01892763, 0.1390315, 0.0830209, 0.01033525, 0.003551753, 0.003808525, 
    0.005278555, 0.01102463, 0.0664382, 0.1967442, 0.1166568, 0.01100688, 
    0.05571592, 0.1197787, 0.0470889, 0.00773033, 0.002612891, 0.002488059, 
    0.01083916, 0.0009098754, 0.04057691, 0.02898758, 0.1575273, 0.1698003, 
    0.06716851, 0.06524734, 0.01084564, 0.01174429, 0.01932656,
  0.001147649, -7.178699e-05, -0.000111046, 0.05726239, 0.0009795019, 
    0.004607435, 0.01369661, 0.004764149, 0.003228285, 0.005114341, 
    0.004650771, 0.03020442, 0.02578315, 0.05426272, 0.09817713, 0.09533916, 
    0.02644141, 0.00853255, 0.006110829, 0.03103023, 0.1042131, 0.007773899, 
    0.0002594583, 0.0006713316, 0.002766938, -1.710365e-06, -0.0002837511, 
    0.06115438, 0.04254729,
  0.007155115, -9.658206e-07, -2.07381e-06, 0.0001656547, 0.04375833, 
    0.000262919, 0.00101524, 0.0004764595, 0.007607829, 0.008357685, 
    0.001517453, 0.02903348, 0.01160138, 0.0001590859, 1.672935e-05, 
    0.0001849907, 2.814356e-05, -4.124461e-05, 0.001010368, -7.740643e-06, 
    0.02260393, 0.04664489, 0.001924773, 0.003688636, 0.007592673, 
    0.001142275, -0.0002807348, 0.01274216, 0.03058273,
  0.04016111, 0.05502482, 0.04520212, 0.03404495, 0.06875812, 0.03897724, 
    0.06991489, 0.01567064, 0.1011024, 0.1456714, 0.1308065, 0.1014515, 
    0.1363453, 0.1152332, 0.02622758, 0.01487479, 0.0001194779, 0.006605282, 
    0.009540349, 0.01407175, 0.02179297, 0.04515526, 0.08029716, 0.0742753, 
    0.0742194, 0.07427184, 0.02114555, 0.01545783, 0.004239996,
  0.0880567, 0.09172226, 0.195772, 0.1255105, 0.07934341, 0.09216387, 
    0.244105, 0.145967, 0.1408456, 0.09388553, 0.1325183, 0.1540396, 
    0.1113461, 0.1989487, 0.2862645, 0.1782529, 0.1613544, 0.1670111, 
    0.1203411, 0.1414265, 0.188408, 0.1857135, 0.1300074, 0.1344025, 
    0.1525741, 0.143322, 0.1084878, 0.06310133, 0.03991633,
  0.1917333, 0.2301164, 0.1117629, 0.1222394, 0.01835912, 0.08832353, 
    0.1852936, 0.116625, 0.1007104, 0.2146077, 0.2255907, 0.1534304, 
    0.1271939, 0.1665286, 0.1323416, 0.1676714, 0.1742802, 0.2386505, 
    0.2609393, 0.16219, 0.1481527, 0.1424326, 0.1581564, 0.2743948, 
    0.2114241, 0.1313247, 0.1620234, 0.1770457, 0.1633661,
  0.3091607, 0.2454057, 0.1837333, 0.1238729, 0.1112043, 0.1332508, 
    0.1918792, 0.1847283, 0.211842, 0.1770769, 0.1600772, 0.04520617, 
    0.0766445, 0.2512143, 0.01988145, 0.1538619, 0.1954081, 0.2694875, 
    0.1503921, 0.07264555, 0.1554791, 0.131587, 0.1413517, 0.1896759, 
    0.2355678, 0.1653539, 0.06053389, 0.1975094, 0.2944671,
  0.2079336, 0.280737, 0.271063, 0.2312602, 0.1864375, 0.1592383, 0.1440262, 
    0.1237891, 0.1709772, 0.2924118, 0.1294884, 0.1385041, 0.1515063, 
    0.2059493, 0.1543173, 0.1807618, 0.153332, 0.1081054, 0.07890845, 
    0.1179513, 0.2082405, 0.1462126, 0.1365263, 0.03912061, 0.1016265, 
    0.002592077, -0.001475962, 0.2559092, 0.1646219,
  0.182806, 0.1882205, 0.2532144, 0.2387999, 0.1732153, 0.1724043, 0.2419132, 
    0.23471, 0.1590795, 0.1591461, 0.1802513, 0.1326414, 0.09442346, 
    0.08883647, 0.1523984, 0.1264804, 0.08380415, 0.0963948, 0.1058287, 
    0.126295, 0.1558196, 0.1963419, 0.1473288, 0.1086252, 0.06356151, 
    0.006812074, -0.002526676, 0.01524522, 0.2642855,
  4.385775e-05, 4.385775e-05, 4.385775e-05, 4.385775e-05, 4.385775e-05, 
    4.385775e-05, 4.385775e-05, -5.752991e-05, -2.316121e-05, 1.120749e-05, 
    4.557618e-05, 7.994488e-05, 0.0001143136, 0.0001486823, 0.00103941, 
    0.001073779, 0.001108147, 0.001142516, 0.001176885, 0.001211253, 
    0.001245622, 0.000274128, 0.0002053906, 0.0001366532, 6.791584e-05, 
    -8.215586e-07, -6.955896e-05, -0.0001382964, 4.385775e-05,
  0.0004087718, -4.93201e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.006908392, 
    0.1161711, 0.1393966, 0.1509416, 0.2212201, 0.2267078, 0.2352135, 
    0.180472, 0.09794594, 0.06709323, 0.1851635, 0.2406261, 0.3269414, 
    0.3786019, 0.315355, 0.1457432, 0.01620016,
  0.1558997, 0.2884986, 0.2112469, 0.2820365, 0.05667741, 0.05846747, 
    0.1649935, 0.04597217, 0.06976837, 0.1111805, 0.06436595, 0.007972499, 
    0.1394702, 0.2404461, 0.340323, 0.2883886, 0.2200992, 0.2628474, 
    0.2940043, 0.2918086, 0.3142572, 0.3236616, 0.3174185, 0.2491182, 
    0.2838655, 0.1659608, 0.1643093, 0.1820417, 0.1336258,
  0.2554435, 0.276289, 0.2599545, 0.3222514, 0.2529692, 0.2412135, 0.2157209, 
    0.3126585, 0.2342999, 0.2842538, 0.3025262, 0.233955, 0.2261635, 
    0.2520855, 0.2678288, 0.2696944, 0.2796284, 0.1751276, 0.1971723, 
    0.2013282, 0.2724767, 0.2557016, 0.215868, 0.2516302, 0.2439723, 
    0.2192527, 0.173784, 0.2239358, 0.2288309,
  0.1633916, 0.1775661, 0.2530021, 0.1638468, 0.1742377, 0.2221048, 
    0.1766868, 0.1856713, 0.1057374, 0.1780212, 0.1981634, 0.1790279, 
    0.1753176, 0.1596614, 0.1247941, 0.1367972, 0.221912, 0.1023956, 
    0.1760484, 0.1900242, 0.1811847, 0.1548233, 0.1563402, 0.210655, 
    0.225107, 0.2002717, 0.2015373, 0.2072334, 0.2081946,
  0.0852604, 0.05478171, 0.05195306, 0.09642469, 0.08517445, 0.03974055, 
    0.06020989, 0.0496527, 0.0572492, 0.1013527, 0.09159721, 0.04248592, 
    0.0483636, 0.07127161, 0.0718968, 0.1044095, 0.1328126, 0.1581923, 
    0.1549369, 0.1859267, 0.2097548, 0.07799046, 0.1355134, 0.1093518, 
    0.04356846, 0.1353592, 0.1633572, 0.1041842, 0.1451752,
  4.761657e-05, 6.816247e-06, 0.02928995, 0.03972671, 0.01093458, 0.0338886, 
    0.02049569, 0.0001380098, 0.04213312, 0.08792829, 0.1597265, 0.06919596, 
    0.02909857, 0.047918, 0.04981249, 0.08456694, 0.03799438, 0.05044855, 
    0.1045016, 0.03457339, 0.1016095, 0.02771602, 0.01410501, 0.01153747, 
    0.03474453, 0.07154211, 0.07318008, 0.03787456, 0.01973645,
  2.198563e-07, 0.001027025, 0.0008074808, 0.0009156348, 0.0117274, 
    0.1021809, 0.106689, 0.01741206, 0.06698103, 0.009731249, 0.0005858314, 
    0.002140008, 0.002754965, 0.04259748, 0.03791201, 0.01768203, 0.03593734, 
    0.06934433, 0.05215893, 0.007587808, 0.0001482924, 3.898766e-07, 
    5.855029e-08, 0.001746607, 0.01920981, 0.04017273, 0.002801201, 
    0.0001934252, 4.477107e-07,
  1.146281e-05, 0.2471901, 0.1917421, 0.08467595, 0.04972751, 0.01370889, 
    0.05449306, 0.03672296, 0.1209838, 0.01953564, 0.03392714, 0.03281672, 
    0.1310011, 0.06151763, 0.0118612, 0.01227197, 0.04247821, 0.03972767, 
    0.008928647, 0.001681712, 0.002164073, 0.00238543, 0.004357819, 
    0.0399177, 0.1417196, 0.007515455, 0.0624518, 0.001877996, 2.069274e-06,
  0.04772951, 0.1264254, 0.08382378, 0.006568209, 0.003128973, 0.003993297, 
    0.005429414, 0.01062234, 0.0671361, 0.2111734, 0.09721474, 0.01106715, 
    0.06124593, 0.1195716, 0.04512846, 0.006946534, 0.004053978, 0.001959309, 
    0.0128858, 0.0006799826, 0.05836843, 0.02957021, 0.1791659, 0.1636487, 
    0.08867221, 0.06052911, 0.01354012, 0.02687268, 0.02921077,
  0.0007362512, 0.0006833752, 0.001027752, 0.08735959, 0.0008892011, 
    0.007000202, 0.01868177, 0.0050492, 0.003373794, 0.003954764, 
    0.004414617, 0.02017643, 0.02479295, 0.08874141, 0.1136551, 0.0933995, 
    0.02308633, 0.0009668152, 0.007536987, 0.03740212, 0.1247895, 
    0.007170376, 0.0003795447, 0.0009801572, 0.004674767, 7.662058e-06, 
    -6.346445e-05, 0.06149561, 0.03373359,
  0.0008427593, 0.0005312859, 1.623812e-07, 0.0003641892, 0.05552296, 
    0.0004587763, 0.0009920939, 0.0005374242, 0.006810164, 0.01593967, 
    0.002449651, 0.03280781, 0.01816101, 6.815367e-05, 1.17374e-05, 
    8.62962e-05, 0.0003046944, -3.06486e-05, 0.005225662, 6.972794e-07, 
    0.01045606, 0.04669817, 0.001922544, 0.004319254, 0.003671901, 
    0.001366197, -0.0001659419, 0.008812703, 0.03653834,
  0.02938022, 0.04758905, 0.0364954, 0.03709502, 0.07368337, 0.03787997, 
    0.09838051, 0.03462614, 0.1132166, 0.1601478, 0.139991, 0.09854195, 
    0.1303851, 0.1068092, 0.02675755, 0.009606476, 0.0002983925, 0.01202049, 
    0.003605668, 0.009872297, 0.01306325, 0.0408122, 0.07261701, 0.06080799, 
    0.06350216, 0.06396828, 0.02457129, 0.002346143, 0.006443332,
  0.0691835, 0.08174413, 0.1828758, 0.1196227, 0.07581691, 0.08226842, 
    0.2534864, 0.1071017, 0.1184394, 0.08838314, 0.1274448, 0.1516057, 
    0.1163482, 0.1803082, 0.2855488, 0.1822106, 0.162022, 0.1548998, 0.13616, 
    0.1272952, 0.1919306, 0.1999517, 0.127546, 0.142517, 0.1558522, 
    0.1206251, 0.08090068, 0.05671803, 0.03439207,
  0.1750759, 0.2305175, 0.1146264, 0.1114615, 0.02204369, 0.09913154, 
    0.1996501, 0.1643361, 0.1713608, 0.25064, 0.2325571, 0.1783616, 
    0.1352971, 0.1572876, 0.1261398, 0.1670738, 0.1675813, 0.2180229, 
    0.2527013, 0.173499, 0.1548111, 0.1438224, 0.1524962, 0.2995695, 
    0.2227042, 0.1550808, 0.1664995, 0.1549185, 0.1515523,
  0.2924018, 0.2421075, 0.1826234, 0.1194769, 0.1027039, 0.1220167, 0.197161, 
    0.2250719, 0.2661247, 0.198663, 0.1593318, 0.1226348, 0.1212773, 
    0.3013536, 0.0489159, 0.1671645, 0.1743288, 0.2962892, 0.1635756, 
    0.06601164, 0.142976, 0.129498, 0.1593615, 0.21476, 0.2262724, 0.1727962, 
    0.05781024, 0.1852153, 0.2830158,
  0.2021886, 0.2608561, 0.2587216, 0.2245532, 0.1742844, 0.1362322, 
    0.1433886, 0.1210042, 0.1620603, 0.2713791, 0.1762352, 0.2069598, 
    0.2576338, 0.2592923, 0.1934966, 0.1789517, 0.1445258, 0.1049705, 
    0.07737871, 0.09163858, 0.1999556, 0.1349667, 0.1297371, 0.05383036, 
    0.0960296, 0.009372747, 0.0004867523, 0.288139, 0.1592266,
  0.2085054, 0.2173855, 0.2821301, 0.2414617, 0.1720314, 0.170316, 0.2461324, 
    0.2429959, 0.1646454, 0.2093231, 0.1819341, 0.1237941, 0.1002154, 
    0.07484241, 0.1379043, 0.1053545, 0.08650596, 0.09460824, 0.09684918, 
    0.1296829, 0.1784738, 0.1970746, 0.2044214, 0.1850542, 0.1498985, 
    0.04551854, 0.001352777, 0.151758, 0.306823,
  0.0001984276, 0.0001812432, 0.0001640589, 0.0001468745, 0.0001296902, 
    0.0001125058, 9.532146e-05, 0.0005063417, 0.0008418875, 0.001177433, 
    0.001512979, 0.001848525, 0.002184071, 0.002519616, -0.001342519, 
    -0.00115006, -0.0009576, -0.0007651406, -0.0005726811, -0.0003802217, 
    -0.0001877622, 0.002069614, 0.001558793, 0.001047972, 0.0005371513, 
    2.63304e-05, -0.0004844905, -0.0009953113, 0.000212175,
  0.01354727, -0.000234678, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0003262977, 
    0.02085651, 0.1749489, 0.1475596, 0.1467393, 0.2175361, 0.2681531, 
    0.334772, 0.2528671, 0.213099, 0.1573875, 0.235164, 0.2439423, 0.3327569, 
    0.3816194, 0.3295436, 0.2327451, 0.04597342,
  0.1399082, 0.2916878, 0.2205909, 0.325289, 0.1131745, 0.1103, 0.1757626, 
    0.1512238, 0.1546081, 0.1880801, 0.1259178, 0.07374505, 0.1707083, 
    0.2405961, 0.349179, 0.3300413, 0.2275151, 0.2838098, 0.3048407, 
    0.2859569, 0.2804678, 0.3010924, 0.3130435, 0.2368218, 0.305425, 
    0.169744, 0.155468, 0.1888068, 0.1482318,
  0.2749183, 0.2783204, 0.2626536, 0.3379407, 0.2444215, 0.2225311, 0.221352, 
    0.3019579, 0.2462724, 0.2845137, 0.3184359, 0.2388288, 0.230178, 
    0.2490721, 0.2775742, 0.2376903, 0.2953808, 0.1971272, 0.1913263, 
    0.1897866, 0.2518762, 0.2581295, 0.2041857, 0.2736074, 0.2467998, 
    0.2066068, 0.1754809, 0.2024266, 0.231535,
  0.1722211, 0.1797009, 0.2555496, 0.1470671, 0.1709819, 0.2334987, 
    0.1736378, 0.1957908, 0.103355, 0.1888981, 0.1756676, 0.1683101, 
    0.1519462, 0.1477879, 0.1322795, 0.1139195, 0.2135212, 0.1051476, 
    0.1848954, 0.1629646, 0.1836818, 0.1664285, 0.1889339, 0.200738, 
    0.2040318, 0.1930456, 0.1983024, 0.1960022, 0.2177688,
  0.07558002, 0.05024734, 0.05233218, 0.09667115, 0.09172999, 0.05665128, 
    0.05781702, 0.04300871, 0.06510276, 0.09728787, 0.07618064, 0.0390261, 
    0.04446832, 0.07497189, 0.05883269, 0.102022, 0.144132, 0.1299285, 
    0.1628927, 0.1751296, 0.2058711, 0.0735643, 0.1161386, 0.106058, 
    0.03522602, 0.1154161, 0.1515685, 0.09533908, 0.135106,
  5.699803e-05, 6.188912e-06, 0.03115333, 0.03862225, 0.01007031, 0.037053, 
    0.02106822, 4.565159e-05, 0.04573834, 0.08562402, 0.1439864, 0.05196962, 
    0.0333887, 0.04696478, 0.04602412, 0.07985663, 0.04737417, 0.04490349, 
    0.1007466, 0.03361876, 0.1100384, 0.02113197, 0.01631436, 0.009528202, 
    0.04067043, 0.07635545, 0.06630625, 0.03401566, 0.01601398,
  4.330614e-07, 0.001159639, 0.0005144454, 0.001395237, 0.0130085, 0.1057033, 
    0.1187015, 0.02987623, 0.0758635, 0.007749607, 0.0009850035, 0.002274689, 
    0.00214638, 0.03199933, 0.03319623, 0.02215432, 0.04263203, 0.08294103, 
    0.04904975, 0.005937253, 7.020086e-05, 8.041375e-07, 9.588003e-08, 
    0.0008176573, 0.01615766, 0.05566447, 0.003867856, 0.0003441015, 
    2.640364e-06,
  8.457055e-05, 0.2501263, 0.2041779, 0.1095244, 0.05827301, 0.02701094, 
    0.05682406, 0.05519318, 0.1383881, 0.02196196, 0.04127228, 0.03364887, 
    0.1445365, 0.08026172, 0.02714845, 0.01822529, 0.05636154, 0.05259066, 
    0.008837728, 0.002202298, 0.003397634, 0.00737931, 0.002965756, 
    0.0515369, 0.1712572, 0.007734883, 0.07686563, 0.003544541, -2.116487e-06,
  0.08538005, 0.1487778, 0.1058073, 0.006151757, 0.003497737, 0.004945768, 
    0.006943437, 0.014043, 0.07649821, 0.2041469, 0.1064126, 0.0134373, 
    0.08310613, 0.1345806, 0.04461738, 0.006414387, 0.008123568, 0.001655305, 
    0.006572885, 0.0009944468, 0.05192006, 0.03049646, 0.175532, 0.1874457, 
    0.1081218, 0.05966119, 0.01166785, 0.0314359, 0.03948875,
  0.009860381, 0.01226958, 0.01069748, 0.1197165, 0.001172984, 0.01044214, 
    0.03392754, 0.008081733, 0.005412527, 0.004416368, 0.006164676, 
    0.02055612, 0.03628576, 0.1033133, 0.1276795, 0.1029606, 0.0329204, 
    0.00120188, 0.01895649, 0.04474094, 0.1467475, 0.009607795, 0.0008067438, 
    0.001693419, 0.00675816, 1.361623e-05, 1.231899e-06, 0.04574587, 
    0.04797101,
  -1.488355e-06, 0.0001427941, 1.984335e-07, 0.0001250546, 0.08751255, 
    0.002221183, 0.001374843, 0.001386632, 0.007857691, 0.02627087, 
    0.002643532, 0.03813158, 0.02653411, 8.679573e-05, 5.188082e-05, 
    9.824431e-06, 0.00152683, 0.0005447185, 0.0004212873, 2.163599e-06, 
    0.007604342, 0.04395454, 0.002264189, 0.005553582, 0.004132624, 
    0.001999645, -5.71045e-05, 0.001763661, 0.02768158,
  0.008242782, 0.02695146, 0.01184672, 0.02603755, 0.07776043, 0.04385655, 
    0.08174326, 0.03495969, 0.1248228, 0.1750854, 0.1541705, 0.094616, 
    0.1218808, 0.1041312, 0.02038751, 0.006081034, -2.47124e-05, 0.01722841, 
    3.310797e-05, 0.004476885, 0.009976503, 0.02413849, 0.05517534, 
    0.04736994, 0.05634835, 0.05950464, 0.0115225, 0.0001056219, 0.004612464,
  0.05415812, 0.06070402, 0.1703384, 0.1161109, 0.07512844, 0.06051371, 
    0.2475784, 0.07319526, 0.09657491, 0.09251687, 0.1280632, 0.1413141, 
    0.1168882, 0.1615096, 0.2623867, 0.1830214, 0.1740484, 0.1475236, 
    0.1244405, 0.1050728, 0.1922217, 0.2008341, 0.1307291, 0.153573, 
    0.1519739, 0.1148483, 0.06974214, 0.05584017, 0.03731065,
  0.1614396, 0.2460016, 0.1064415, 0.09413229, 0.03103297, 0.1102879, 
    0.1929386, 0.1860607, 0.2504511, 0.256311, 0.2276057, 0.2022101, 
    0.1442297, 0.1613467, 0.1388352, 0.1755438, 0.1784264, 0.2013425, 
    0.2470909, 0.1779233, 0.161163, 0.1469235, 0.1497855, 0.2802362, 
    0.2224374, 0.1789918, 0.150553, 0.1663463, 0.1629536,
  0.2856389, 0.243414, 0.1764039, 0.1221438, 0.09210999, 0.1169846, 
    0.1954165, 0.2213223, 0.2971701, 0.1931799, 0.1394288, 0.1380497, 
    0.1664417, 0.2970424, 0.06301936, 0.1684564, 0.1522089, 0.312224, 
    0.1539819, 0.0529312, 0.1362957, 0.1251014, 0.1836229, 0.2223174, 
    0.2301993, 0.1762991, 0.05847967, 0.1733519, 0.2747944,
  0.1821362, 0.2609398, 0.2536709, 0.2126751, 0.1701925, 0.116694, 0.1291735, 
    0.1225067, 0.154705, 0.2515907, 0.2056727, 0.1886497, 0.2598605, 
    0.2806626, 0.187617, 0.1851822, 0.1419497, 0.1006579, 0.08919093, 
    0.07464392, 0.1820591, 0.1296728, 0.1210212, 0.07100923, 0.08696872, 
    0.06269551, 0.01648022, 0.2910411, 0.167099,
  0.2052865, 0.2123683, 0.2866193, 0.2456205, 0.1715847, 0.1702088, 
    0.2451941, 0.2515638, 0.1636685, 0.2101935, 0.1711159, 0.1065112, 
    0.08735719, 0.05633428, 0.1280255, 0.09853135, 0.08187684, 0.09015312, 
    0.08390703, 0.1292274, 0.1695873, 0.1970629, 0.1971371, 0.2457394, 
    0.1871129, 0.1014837, 0.0986674, 0.1555883, 0.3290365,
  0.01256921, 0.01144051, 0.0103118, 0.0091831, 0.008054395, 0.006925691, 
    0.005796986, 0.01005492, 0.01317882, 0.01630273, 0.01942663, 0.02255054, 
    0.02567444, 0.02879835, 0.0344607, 0.03532274, 0.03618479, 0.03704683, 
    0.03790887, 0.03877092, 0.03963296, 0.03713481, 0.03427757, 0.03142032, 
    0.02856308, 0.02570583, 0.02284859, 0.01999135, 0.01347218,
  0.03691494, 0.007345036, -7.958776e-05, 0, 0, -1.95097e-05, 0, 0, 0, 0, 
    -9.757422e-05, 0.03074171, 0.04542438, 0.2263226, 0.1541917, 0.1523049, 
    0.242752, 0.2930972, 0.3808028, 0.3799103, 0.3163534, 0.2924886, 
    0.2635588, 0.2367327, 0.3293951, 0.3801928, 0.3302243, 0.2898322, 0.082076,
  0.1716296, 0.2904692, 0.2091455, 0.3433236, 0.1904704, 0.153412, 0.1982428, 
    0.2387891, 0.254401, 0.2283493, 0.2065291, 0.1240662, 0.1638207, 
    0.2338507, 0.3603419, 0.358731, 0.2773457, 0.2967704, 0.3057684, 
    0.283627, 0.339519, 0.3114665, 0.3101268, 0.2476054, 0.2644386, 
    0.2182738, 0.1646003, 0.2059061, 0.1677825,
  0.2976517, 0.3016182, 0.2510979, 0.3319805, 0.2456095, 0.2289201, 
    0.2079193, 0.299781, 0.2796022, 0.3078732, 0.3441429, 0.2351589, 
    0.2095366, 0.2690733, 0.3038706, 0.2409956, 0.2864323, 0.1899109, 
    0.2068014, 0.1966214, 0.2236592, 0.2238514, 0.1808121, 0.2819964, 
    0.1916232, 0.2219155, 0.1832801, 0.1946929, 0.2361069,
  0.165398, 0.1788681, 0.262241, 0.1479529, 0.1722154, 0.2143862, 0.1765961, 
    0.1869737, 0.1196328, 0.1647142, 0.1681971, 0.1775202, 0.1378747, 
    0.1457117, 0.1347106, 0.100431, 0.2240802, 0.1191958, 0.1918346, 
    0.1695314, 0.1697395, 0.1616579, 0.1858574, 0.1759289, 0.2168818, 
    0.2005984, 0.2092108, 0.1822247, 0.2132328,
  0.06586222, 0.04530433, 0.05250648, 0.1078736, 0.1065711, 0.06048687, 
    0.05854166, 0.0409602, 0.06794637, 0.1026757, 0.06891339, 0.0627088, 
    0.05526977, 0.07618631, 0.06686195, 0.1044891, 0.1512008, 0.109568, 
    0.1789132, 0.1697083, 0.219591, 0.08184116, 0.09903838, 0.1078225, 
    0.04175184, 0.09137007, 0.1572456, 0.09414881, 0.1285229,
  0.001846261, 1.880645e-06, 0.03657262, 0.03649344, 0.01260311, 0.03720815, 
    0.02887621, 1.833381e-05, 0.05010847, 0.08456594, 0.1660152, 0.04472625, 
    0.03711345, 0.04407188, 0.04672974, 0.06627113, 0.06140584, 0.04277327, 
    0.08928055, 0.05906748, 0.1214206, 0.02319333, 0.0173594, 0.007409702, 
    0.05958379, 0.0809367, 0.07361753, 0.04362527, 0.0139245,
  3.486031e-07, 0.006278882, 0.0003297005, 0.001716776, 0.0143193, 0.1102096, 
    0.1120108, 0.02905549, 0.08883126, 0.007605764, 0.001770214, 0.004027333, 
    0.01124338, 0.02819083, 0.03152516, 0.02739603, 0.04840935, 0.09092249, 
    0.0518207, 0.00486336, 2.765407e-05, 1.132734e-06, 1.453886e-07, 
    0.001037019, 0.01501722, 0.03363004, 0.005201186, 0.0007480555, 
    4.091716e-06,
  -3.637634e-05, 0.2373001, 0.2231782, 0.1479732, 0.0677293, 0.03296741, 
    0.05977168, 0.05996808, 0.1557967, 0.02362821, 0.03467343, 0.03489076, 
    0.1587558, 0.0909438, 0.0270971, 0.03142661, 0.06189955, 0.06564328, 
    0.009747555, 0.00202347, 0.003590599, 0.0073834, 0.01022192, 0.07443879, 
    0.1987988, 0.01189625, 0.08064492, 0.004289481, 1.953258e-05,
  0.1033029, 0.1877041, 0.1365944, 0.00909154, 0.003482545, 0.003866894, 
    0.005101329, 0.0136032, 0.1022752, 0.2432493, 0.1194128, 0.01825924, 
    0.09653367, 0.1483497, 0.04478061, 0.005256951, 0.009312686, 0.001695707, 
    0.00663965, 0.0009937859, 0.04116518, 0.03771493, 0.2017773, 0.2125598, 
    0.1400481, 0.05871559, 0.01016473, 0.03425355, 0.05185585,
  0.03642678, 0.009840677, 0.01492109, 0.1563766, 0.001302827, 0.01302102, 
    0.05126351, 0.01043588, 0.005172664, 0.00475011, 0.005845215, 0.01962722, 
    0.04160772, 0.1059027, 0.1413234, 0.1096537, 0.04097651, 0.001713816, 
    0.02315742, 0.05063868, 0.1764339, 0.009928337, 0.00077422, 0.003459504, 
    0.00483095, 1.116252e-05, 0.001832183, 0.03341984, 0.0745559,
  9.146782e-06, 5.835362e-06, 2.877316e-07, 0.002667085, 0.09943331, 
    0.002049807, 0.008319998, 0.001338592, 0.02579751, 0.02058161, 
    0.00251753, 0.0385684, 0.02876935, 8.098898e-05, 0.0001540616, 
    7.930544e-06, 0.008359203, 0.0003450234, 2.298603e-05, -1.919853e-06, 
    0.002750945, 0.04596628, 0.003893102, 0.008367386, 0.00873073, 
    0.003835263, -0.0002169582, 0.00537689, 0.01199707,
  0.000495685, 0.00604592, 0.00167929, 0.01839809, 0.07845785, 0.04271526, 
    0.0605227, 0.03226858, 0.1292343, 0.1856493, 0.1486648, 0.1022331, 
    0.1329185, 0.1017537, 0.02426179, 0.006341385, 0.0001722707, 0.01779233, 
    0.0001358301, 0.007276401, 0.006064285, 0.02562917, 0.03828251, 
    0.04486432, 0.04878429, 0.05505582, 0.004759716, 0.0002628418, 0.001302872,
  0.04344381, 0.04518301, 0.1608503, 0.1107327, 0.0798872, 0.04411216, 
    0.2262019, 0.05079508, 0.07976858, 0.0857167, 0.1182713, 0.1412888, 
    0.1137543, 0.1524743, 0.2453638, 0.181345, 0.1715528, 0.1376469, 
    0.1306809, 0.1043002, 0.2129278, 0.1879364, 0.12847, 0.1741435, 
    0.1443534, 0.116488, 0.06492455, 0.05563113, 0.03596104,
  0.15165, 0.2369023, 0.1109117, 0.07894587, 0.02353544, 0.09883803, 
    0.1762835, 0.230468, 0.2719181, 0.2637301, 0.2267192, 0.2106268, 
    0.1399231, 0.1585909, 0.1731353, 0.1896916, 0.1604858, 0.2032023, 
    0.2461372, 0.1727564, 0.1667562, 0.1668607, 0.1532262, 0.3045973, 
    0.2317061, 0.1739512, 0.1418531, 0.1469034, 0.1710941,
  0.295059, 0.2529491, 0.1608594, 0.1154104, 0.08857444, 0.1186045, 
    0.2084186, 0.2364388, 0.2815765, 0.1737591, 0.1541144, 0.1448794, 
    0.1678427, 0.285262, 0.06260037, 0.1650856, 0.1477072, 0.3280852, 
    0.1661518, 0.04076205, 0.1362444, 0.1268044, 0.2533021, 0.2282037, 
    0.2457819, 0.1850357, 0.07349643, 0.1630266, 0.2975145,
  0.1734826, 0.2699634, 0.2588745, 0.206287, 0.1726651, 0.1017898, 0.1171884, 
    0.1319982, 0.1507583, 0.2450507, 0.2015637, 0.1642455, 0.2492924, 
    0.2711027, 0.234495, 0.1894944, 0.1363337, 0.09618436, 0.09631825, 
    0.06584269, 0.1670032, 0.1232385, 0.1212534, 0.06860468, 0.08818031, 
    0.1878738, 0.06251855, 0.2722149, 0.1807175,
  0.2191162, 0.2027122, 0.3072951, 0.2547186, 0.1766064, 0.1805022, 
    0.2414901, 0.2413674, 0.1661347, 0.2247485, 0.1756534, 0.109498, 
    0.07847249, 0.04843816, 0.1258336, 0.1059869, 0.07957535, 0.07857179, 
    0.07512867, 0.1213097, 0.1571416, 0.1989799, 0.2055383, 0.2490754, 
    0.2127192, 0.1478527, 0.20006, 0.1450631, 0.3487562,
  0.02753257, 0.0255592, 0.02358584, 0.02161248, 0.01963911, 0.01766575, 
    0.01569238, 0.02684464, 0.03062025, 0.03439585, 0.03817146, 0.04194707, 
    0.04572268, 0.04949829, 0.04624642, 0.04677605, 0.04730568, 0.0478353, 
    0.04836493, 0.04889455, 0.04942418, 0.05293445, 0.05060258, 0.04827071, 
    0.04593883, 0.04360697, 0.0412751, 0.03894322, 0.02911126,
  0.06373479, 0.03909881, 0.02206558, 0.001182602, -5.393467e-06, 
    -0.001262875, -0.0009178801, -0.0008870203, 0.0001016367, 2.942268e-05, 
    0.01375753, 0.04240868, 0.06615587, 0.2614735, 0.169748, 0.2127745, 
    0.2820015, 0.3734984, 0.4134063, 0.4373541, 0.4016268, 0.3323204, 
    0.2862723, 0.2509492, 0.3393095, 0.4015564, 0.364309, 0.2950874, 0.1105619,
  0.2108283, 0.3727297, 0.1902685, 0.3644409, 0.2693445, 0.1652908, 
    0.2032054, 0.3050427, 0.2888863, 0.285352, 0.2625604, 0.1350616, 
    0.1544782, 0.2537419, 0.3871686, 0.3314564, 0.2719247, 0.3045045, 
    0.3009026, 0.2996274, 0.3399001, 0.3066186, 0.2970568, 0.2235889, 
    0.2985871, 0.2110612, 0.1742482, 0.2602098, 0.1530751,
  0.3310899, 0.3572819, 0.3316239, 0.3629214, 0.3135085, 0.2357569, 
    0.2040189, 0.2900607, 0.3025221, 0.3510017, 0.3392609, 0.2469391, 0.228, 
    0.280189, 0.2901725, 0.2016262, 0.2668183, 0.1858843, 0.1785713, 
    0.195324, 0.2289628, 0.208885, 0.2059995, 0.2600308, 0.2235718, 
    0.2550602, 0.204321, 0.1960598, 0.2224475,
  0.1950867, 0.1676756, 0.2450085, 0.1583283, 0.1759859, 0.2431125, 
    0.1997039, 0.2202769, 0.1522574, 0.1826623, 0.1630901, 0.1872157, 
    0.1329582, 0.1417807, 0.1289679, 0.08583184, 0.2272355, 0.124578, 
    0.1826442, 0.162098, 0.1733573, 0.1747807, 0.1744169, 0.1670198, 0.23493, 
    0.2069677, 0.2163195, 0.1838914, 0.1946672,
  0.06614749, 0.04579075, 0.04564405, 0.1284413, 0.1111839, 0.06945316, 
    0.06194009, 0.06081845, 0.06721935, 0.11052, 0.0673632, 0.04329117, 
    0.06481972, 0.08399171, 0.06340317, 0.1083409, 0.1648741, 0.1091914, 
    0.172499, 0.167041, 0.2172253, 0.08868408, 0.08993194, 0.1097217, 
    0.05299072, 0.09105895, 0.1584003, 0.09765107, 0.1237458,
  0.01810426, -2.004732e-05, 0.03970392, 0.03509204, 0.0174081, 0.0398331, 
    0.03732095, -1.136535e-05, 0.0547593, 0.08314557, 0.1659394, 0.04572855, 
    0.04640656, 0.04453753, 0.05477142, 0.0571735, 0.06003881, 0.0387291, 
    0.08186787, 0.05260831, 0.1260014, 0.03078307, 0.02102411, 0.006114093, 
    0.0759747, 0.1060893, 0.08314881, 0.06783763, 0.01590475,
  2.449684e-07, 0.02205341, 0.0005223459, 0.003722333, 0.0158869, 0.09681271, 
    0.09993617, 0.02211637, 0.1167749, 0.00417733, 0.001611745, 0.004330585, 
    0.01505777, 0.03282082, 0.02202255, 0.02571168, 0.0585691, 0.08742054, 
    0.05295972, 0.006848196, 2.301945e-06, 1.906291e-05, 1.454567e-07, 
    0.001249137, 0.0246377, 0.03910628, 0.004766688, 0.002273618, 2.108294e-06,
  0.000160726, 0.2105365, 0.2449307, 0.1749431, 0.06222247, 0.02800359, 
    0.05889513, 0.07424599, 0.1319931, 0.01712658, 0.03712082, 0.03839634, 
    0.156299, 0.07037064, 0.02135305, 0.03202911, 0.05298316, 0.06591816, 
    0.009876832, 0.002324959, 0.005209067, 0.01079808, 0.009853714, 
    0.07488422, 0.1885077, 0.02125171, 0.08771686, 0.003158589, 2.77542e-05,
  0.07368507, 0.1784258, 0.1458134, 0.01767748, 0.002441808, 0.004252731, 
    0.006273657, 0.011837, 0.1158706, 0.2739163, 0.1158585, 0.01802402, 
    0.08078548, 0.1144319, 0.03237845, 0.004543849, 0.007678313, 0.00239011, 
    0.002026503, 0.001967015, 0.03071793, 0.03432664, 0.1726568, 0.2407916, 
    0.1635848, 0.05680987, 0.01245092, 0.0211298, 0.03571796,
  0.0298939, 0.002954815, 0.004099767, 0.2100459, 0.001175395, 0.008876559, 
    0.05545899, 0.01294987, 0.005508614, 0.00580496, 0.007010559, 0.01714578, 
    0.02665742, 0.09259401, 0.130478, 0.1075291, 0.03486158, 0.0002796043, 
    0.02841282, 0.04585098, 0.1826705, 0.00886766, 0.001481375, 0.004536549, 
    0.002667733, 8.003932e-06, 0.002064471, 0.02121913, 0.06397322,
  3.255388e-06, 1.897685e-06, 2.783514e-07, 0.0003367877, 0.05958788, 
    0.001515248, 0.03372171, 0.001031874, 0.05425767, 0.01120161, 
    0.002503779, 0.0389409, 0.02865685, 0.0001223425, 9.751746e-05, 
    0.0007046754, 0.01487209, 0.0009220152, 1.024855e-05, 0.0002493442, 
    0.0008189622, 0.0388209, 0.004871076, 0.01303969, 0.00996566, 
    0.007529742, 2.968537e-06, 0.0001638655, 0.001567487,
  -2.465734e-05, 0.001388849, 0.0005498665, 0.01511912, 0.08001246, 
    0.0293767, 0.02189513, 0.02666813, 0.1318899, 0.1889449, 0.1556497, 
    0.1053496, 0.1327389, 0.08720995, 0.03169845, 0.01322059, 0.004264735, 
    0.01709903, 0.0006145404, 0.003008802, 0.001668797, 0.02605954, 
    0.03141289, 0.05872964, 0.05095006, 0.05790658, 0.005190119, 
    0.0004746377, 0.0007876242,
  0.04228019, 0.03233151, 0.1608875, 0.1052951, 0.0900078, 0.03748875, 
    0.2214354, 0.03778103, 0.06285878, 0.09727685, 0.1066167, 0.1283657, 
    0.1187987, 0.1502164, 0.2368218, 0.1776325, 0.1810332, 0.1319761, 
    0.1241572, 0.1121911, 0.2128708, 0.1882437, 0.1132834, 0.1619527, 
    0.1397919, 0.1203046, 0.06378962, 0.05861738, 0.03649245,
  0.1570838, 0.2316861, 0.0974216, 0.067147, 0.0250697, 0.08823653, 
    0.1875013, 0.2486339, 0.2597551, 0.2748962, 0.2136039, 0.208542, 
    0.1440745, 0.1663529, 0.2106594, 0.1971873, 0.1744928, 0.2302343, 
    0.255761, 0.1814304, 0.1754836, 0.1733406, 0.1703951, 0.2733183, 
    0.2513473, 0.1990318, 0.154053, 0.1416606, 0.1594762,
  0.295265, 0.2753383, 0.1792685, 0.1159091, 0.09706823, 0.1317955, 
    0.2167619, 0.2439037, 0.2668293, 0.1890474, 0.1467536, 0.142772, 
    0.1484099, 0.2954306, 0.05217859, 0.1675204, 0.1674853, 0.3521094, 
    0.190431, 0.02990701, 0.1845847, 0.1401919, 0.2695975, 0.2199934, 
    0.2109557, 0.1871903, 0.1377316, 0.178204, 0.3249623,
  0.1829374, 0.227594, 0.2510986, 0.193383, 0.1472326, 0.08584996, 0.1033757, 
    0.1258568, 0.1455437, 0.2472827, 0.2094581, 0.181868, 0.2243259, 
    0.2663912, 0.2537315, 0.183921, 0.1771906, 0.09548954, 0.1246721, 
    0.09779968, 0.1506136, 0.1275759, 0.1259977, 0.06328852, 0.09169015, 
    0.2568599, 0.1235598, 0.2771994, 0.1879762,
  0.2453833, 0.2553382, 0.3671751, 0.2729279, 0.1693179, 0.1784483, 
    0.2396528, 0.2319747, 0.1804201, 0.2223863, 0.1724335, 0.1045072, 
    0.06578498, 0.04379331, 0.109345, 0.09739949, 0.07138988, 0.07441069, 
    0.07267369, 0.1173561, 0.1430943, 0.1943793, 0.2138716, 0.2265471, 
    0.2036242, 0.1805845, 0.229248, 0.125594, 0.3523249,
  0.07186773, 0.06564563, 0.05942353, 0.05320143, 0.04697933, 0.04075723, 
    0.03453514, 0.04933641, 0.05266127, 0.05598613, 0.059311, 0.06263586, 
    0.06596072, 0.06928559, 0.05993903, 0.06309835, 0.06625767, 0.06941699, 
    0.07257631, 0.07573564, 0.07889496, 0.09978849, 0.09952641, 0.09926432, 
    0.09900223, 0.09874015, 0.09847806, 0.09821597, 0.0768454,
  0.08012234, 0.04464604, 0.03877037, 0.009576204, 0.004693232, 0.02645295, 
    0.01564357, 0.01630091, 0.005544887, 0.0006240147, 0.02422315, 
    0.04933656, 0.07268126, 0.2520733, 0.2384382, 0.3173385, 0.3408171, 
    0.4403479, 0.4556291, 0.4708441, 0.5009226, 0.3790201, 0.2914814, 
    0.2469625, 0.3232999, 0.4179058, 0.3806984, 0.3023163, 0.1295856,
  0.2559651, 0.3949221, 0.276728, 0.3464353, 0.3172658, 0.1653941, 0.2154878, 
    0.3404848, 0.336123, 0.3251744, 0.3542626, 0.1420168, 0.1524859, 
    0.2824294, 0.4632371, 0.3676095, 0.2807022, 0.3792493, 0.3111567, 
    0.2462874, 0.3075958, 0.324515, 0.3050908, 0.2240594, 0.3233465, 
    0.1750549, 0.1424634, 0.3133323, 0.1945512,
  0.3351161, 0.3537861, 0.3188368, 0.3926296, 0.2852071, 0.2618671, 
    0.2534328, 0.3193449, 0.3305848, 0.3299359, 0.3514369, 0.2655664, 
    0.255757, 0.2756076, 0.3013161, 0.223003, 0.2692339, 0.2060344, 
    0.2096098, 0.1930875, 0.2322659, 0.225218, 0.1685606, 0.2678109, 
    0.1642623, 0.2645025, 0.2253671, 0.2054496, 0.2306413,
  0.1952088, 0.1627567, 0.2424718, 0.1736486, 0.1877057, 0.2427443, 
    0.2083912, 0.2212579, 0.16331, 0.1825773, 0.1538716, 0.1878779, 0.144879, 
    0.1518742, 0.1175435, 0.08789567, 0.2264193, 0.1253062, 0.1823588, 
    0.1577336, 0.1808375, 0.1872126, 0.1615123, 0.1663096, 0.2224499, 
    0.2041777, 0.2169189, 0.184019, 0.1695872,
  0.08197373, 0.04976726, 0.04081182, 0.1297375, 0.1148102, 0.07701453, 
    0.07318683, 0.0712698, 0.07765026, 0.1355636, 0.07966837, 0.04511872, 
    0.1015848, 0.09200937, 0.09002413, 0.1189283, 0.1657198, 0.1010504, 
    0.1792994, 0.1519604, 0.2249314, 0.0711339, 0.1059336, 0.1176646, 
    0.07227757, 0.105707, 0.161082, 0.09869521, 0.1298696,
  0.02301771, -6.546803e-05, 0.04112499, 0.03336757, 0.04081926, 0.04442533, 
    0.04372841, -4.905105e-05, 0.05757535, 0.08802283, 0.1265444, 0.05576704, 
    0.06031785, 0.05040466, 0.05886043, 0.06344858, 0.06040303, 0.03472561, 
    0.09332684, 0.0581496, 0.1263372, 0.03337645, 0.02280496, 0.006785151, 
    0.08079278, 0.07364079, 0.06280836, 0.08375446, 0.01753923,
  1.618678e-07, 0.08026469, 0.00318384, 0.008725869, 0.0168582, 0.07711684, 
    0.07518092, 0.01193427, 0.1137919, 0.001886113, 0.003763122, 0.006115734, 
    0.0186629, 0.03553642, 0.02588114, 0.02168327, 0.06166828, 0.08800726, 
    0.05187413, 0.01347895, 0.0005156269, 0.001342693, 1.268945e-07, 
    0.000167823, 0.02583466, 0.04163781, 0.00516428, 0.007262364, 
    -2.754516e-06,
  4.997647e-05, 0.1588053, 0.2515469, 0.1755206, 0.04783522, 0.02491979, 
    0.05337008, 0.08144706, 0.1155801, 0.01195044, 0.03783322, 0.04055564, 
    0.1472461, 0.06298491, 0.02022963, 0.03375322, 0.04476834, 0.0594991, 
    0.01148714, 0.001516539, 0.009529601, 0.007972045, 0.004348621, 
    0.05509216, 0.1477722, 0.03150191, 0.09712398, 0.00220171, 1.81348e-05,
  0.03532555, 0.09941565, 0.07324532, 0.0306094, 0.003225541, 0.004738845, 
    0.007502867, 0.01126757, 0.09963539, 0.2346348, 0.1075521, 0.01949581, 
    0.07217255, 0.09573197, 0.03053592, 0.005513886, 0.01189898, 0.003580551, 
    0.002728393, 0.00327577, 0.02484881, 0.02778642, 0.1552787, 0.1706233, 
    0.1464226, 0.04821932, 0.01698696, 0.01697228, 0.03050531,
  0.01115077, 2.322476e-05, -1.4032e-05, 0.2479769, 0.000776688, 0.007954454, 
    0.05047769, 0.01530287, 0.005199952, 0.006105209, 0.0128432, 0.01179256, 
    0.02455699, 0.09026877, 0.1058549, 0.09538124, 0.02913417, 0.0007097546, 
    0.03375117, 0.04924172, 0.1541563, 0.009432253, 0.00351374, 0.009726426, 
    0.001742879, 2.325601e-05, 0.001176408, 0.008396429, 0.02034246,
  1.053699e-06, 6.296857e-07, 1.524146e-07, -5.953726e-05, 0.008249511, 
    0.0001577852, 0.04415526, 0.0004042611, 0.03977692, 0.004657181, 
    0.002477627, 0.04178307, 0.02674032, 0.0002033069, 0.0007101365, 
    0.005595834, 0.0189236, 0.008723894, 1.9186e-05, 1.20948e-05, 
    0.005242684, 0.03667269, 0.006552381, 0.0223976, 0.01457641, 0.009375157, 
    -4.360581e-06, 1.739341e-05, 4.875267e-05,
  -1.972638e-05, 0.0007818525, 0.000380011, 0.009636614, 0.08255671, 
    0.01989557, 0.007929641, 0.02119484, 0.1153363, 0.1711721, 0.1700519, 
    0.1012636, 0.1226988, 0.08277592, 0.04988998, 0.01145954, 0.01223753, 
    0.02619024, 0.001842632, 0.001630261, 0.003341655, 0.02643558, 
    0.03868412, 0.07670654, 0.05698247, 0.07022862, 0.0111932, 0.00113189, 
    0.0008551643,
  0.0464079, 0.03302819, 0.1525455, 0.1042286, 0.08796074, 0.01928227, 
    0.2154528, 0.04108084, 0.05190938, 0.1084851, 0.1008102, 0.1239294, 
    0.127568, 0.1393175, 0.2268437, 0.187999, 0.1772972, 0.1430977, 
    0.1173261, 0.112089, 0.2156432, 0.1956382, 0.1129737, 0.1573276, 
    0.1465083, 0.1241328, 0.07005716, 0.05986064, 0.04417748,
  0.1451765, 0.2225724, 0.1002991, 0.06325776, 0.02789541, 0.1050147, 
    0.2236666, 0.2578768, 0.2439376, 0.26865, 0.2042663, 0.2197548, 
    0.1467283, 0.2122725, 0.2407473, 0.2176781, 0.1832829, 0.2067385, 
    0.2567286, 0.1826935, 0.162024, 0.1868386, 0.17134, 0.3117245, 0.2446047, 
    0.2073244, 0.1692081, 0.1582191, 0.1688144,
  0.3081437, 0.2463486, 0.1852389, 0.1221562, 0.09999873, 0.1232323, 
    0.2384715, 0.2529672, 0.2449635, 0.2099749, 0.1356475, 0.130589, 
    0.1417173, 0.3044043, 0.05008917, 0.1688172, 0.1850105, 0.3781328, 
    0.1945977, 0.04437982, 0.1831739, 0.1480239, 0.2518732, 0.2078634, 
    0.2249389, 0.1917216, 0.1749655, 0.1742636, 0.3023184,
  0.2052481, 0.2405162, 0.26969, 0.1946345, 0.1495546, 0.1260948, 0.1038026, 
    0.1181191, 0.1326207, 0.2480094, 0.2353043, 0.1881021, 0.1945885, 
    0.2720807, 0.2474746, 0.1733171, 0.2518784, 0.09335743, 0.1731637, 
    0.1370579, 0.1431908, 0.1589963, 0.1131454, 0.06943393, 0.09395575, 
    0.2768914, 0.1805962, 0.2795547, 0.2291254,
  0.2811552, 0.2634069, 0.3943903, 0.3252929, 0.2064109, 0.1871431, 
    0.2628843, 0.2365602, 0.1922169, 0.2216074, 0.1736333, 0.09892979, 
    0.054253, 0.04201574, 0.09969106, 0.1189346, 0.08338221, 0.08165781, 
    0.08868945, 0.1199788, 0.1279357, 0.2016532, 0.2266818, 0.2164282, 
    0.1955446, 0.2119479, 0.2511488, 0.09521623, 0.3720949,
  0.1588344, 0.1500731, 0.1413118, 0.1325504, 0.1237891, 0.1150278, 
    0.1062664, 0.1210103, 0.1229471, 0.1248839, 0.1268207, 0.1287575, 
    0.1306943, 0.1326311, 0.1032827, 0.1145811, 0.1258796, 0.137178, 
    0.1484764, 0.1597748, 0.1710732, 0.1809911, 0.1765172, 0.1720434, 
    0.1675695, 0.1630956, 0.1586217, 0.1541478, 0.1658435,
  0.1115285, 0.07558514, 0.03658155, 0.0357632, 0.03741563, 0.07417171, 
    0.05808174, 0.05864962, 0.02109387, 0.01070894, 0.0278801, 0.04987457, 
    0.08973407, 0.222999, 0.2919254, 0.3341527, 0.3248609, 0.4427405, 
    0.4403827, 0.4965041, 0.5395277, 0.3890195, 0.2861217, 0.2779882, 
    0.3418256, 0.4021147, 0.4156418, 0.3045173, 0.1633067,
  0.265734, 0.3593561, 0.1756666, 0.3739535, 0.3680498, 0.1548699, 0.2429076, 
    0.3305929, 0.3825259, 0.3454846, 0.3726175, 0.1325422, 0.1495267, 
    0.3296073, 0.4238841, 0.4055131, 0.3219489, 0.3332893, 0.3394667, 
    0.2703428, 0.32221, 0.2946998, 0.310121, 0.2523211, 0.2860102, 0.1991692, 
    0.1769574, 0.3022055, 0.2385698,
  0.3397857, 0.3970529, 0.3952593, 0.3880483, 0.3251166, 0.3111551, 0.275796, 
    0.3587246, 0.3781435, 0.3399295, 0.3215639, 0.2919479, 0.2704706, 
    0.321683, 0.2962915, 0.2475581, 0.2817146, 0.208319, 0.2087005, 
    0.2104187, 0.2320437, 0.1986857, 0.2440006, 0.2439688, 0.1762996, 
    0.2848565, 0.2294542, 0.192636, 0.2359861,
  0.1878056, 0.1581351, 0.2364814, 0.1687729, 0.1840179, 0.2384198, 
    0.2055496, 0.2125535, 0.1695163, 0.1752692, 0.1652481, 0.1963169, 
    0.1651751, 0.1629389, 0.1073154, 0.1266734, 0.2583378, 0.151341, 
    0.2007971, 0.1943252, 0.1973709, 0.2030746, 0.1584371, 0.1782884, 
    0.2388679, 0.2001356, 0.2335778, 0.1848442, 0.1682044,
  0.08948366, 0.05836318, 0.05830992, 0.1392481, 0.1130915, 0.08252882, 
    0.08760341, 0.08190016, 0.09504476, 0.1875972, 0.1084268, 0.05845008, 
    0.0918722, 0.1113836, 0.1107398, 0.1367024, 0.1661582, 0.1199143, 
    0.1896073, 0.1627088, 0.2169848, 0.08006268, 0.1131751, 0.1348032, 
    0.09473147, 0.1273025, 0.1915321, 0.09991718, 0.1315816,
  0.0249658, 0.0009979814, 0.04866491, 0.0322624, 0.02217616, 0.04437808, 
    0.03756534, 0.0005900127, 0.05507879, 0.07377437, 0.05633899, 0.03066012, 
    0.0966686, 0.05989388, 0.04930128, 0.07332449, 0.06434095, 0.03668817, 
    0.09270056, 0.04811312, 0.1415585, 0.04231369, 0.02621703, 0.006619893, 
    0.09592723, 0.06032817, 0.05626336, 0.0826119, 0.03368262,
  1.107753e-07, 0.05086086, 0.09136654, 0.01672976, 0.02649702, 0.06454921, 
    0.08126651, 0.01284933, 0.1128071, 0.001845703, 0.01980729, 0.02459199, 
    0.02617405, 0.03653564, 0.03282594, 0.03299883, 0.06171535, 0.1082141, 
    0.0466349, 0.02759709, 0.008177399, 0.01178919, 1.394817e-07, 
    9.583958e-05, 0.02989981, 0.03802656, 0.01460187, 0.02218028, 3.144554e-05,
  5.232283e-05, 0.1266454, 0.1983212, 0.1854658, 0.0485164, 0.02673454, 
    0.04606932, 0.08477773, 0.1058865, 0.01202329, 0.05097158, 0.04010949, 
    0.1338843, 0.05411562, 0.02117619, 0.03717683, 0.04130732, 0.05249622, 
    0.01592297, 0.005370045, 0.01472669, 0.00758828, 0.001270502, 0.05409972, 
    0.1250885, 0.03681831, 0.1117261, 0.004293449, 2.434851e-06,
  0.01648727, 0.06051203, 0.04515947, 0.05616689, 0.003817338, 0.006511418, 
    0.009606054, 0.01132962, 0.08740595, 0.217375, 0.1058498, 0.02595274, 
    0.06469723, 0.07833992, 0.03173596, 0.009448131, 0.01422716, 0.006659168, 
    0.004625644, 0.003628996, 0.0256495, 0.02167498, 0.131908, 0.1431776, 
    0.1356723, 0.04599943, 0.01937561, 0.01229092, 0.02865537,
  0.00115843, -6.968351e-06, -2.815608e-05, 0.2742184, 0.001619285, 
    0.008619373, 0.04271913, 0.02214536, 0.00537045, 0.005989831, 0.02156339, 
    0.01161791, 0.02532192, 0.08947439, 0.09958005, 0.08789422, 0.01856962, 
    0.001444708, 0.03825432, 0.06243482, 0.1340387, 0.009782952, 0.007739105, 
    0.01681937, 0.002840596, 1.515648e-05, 2.634904e-05, 0.001846774, 
    0.007523595,
  8.452694e-07, 2.817376e-07, 8.472692e-08, -1.250968e-05, 0.0005909585, 
    2.154436e-06, 0.02818492, 0.0001755186, 0.04176089, 0.02119738, 
    0.003121148, 0.0466542, 0.02559348, 0.004321151, 0.006108643, 0.01212672, 
    0.02419553, 0.03005081, 3.975181e-05, -2.197265e-05, 0.0007347632, 
    0.03158824, 0.008045716, 0.03861066, 0.01970303, 0.01292741, 
    1.531896e-05, 9.989189e-06, 1.147959e-05,
  -2.214428e-05, -5.229981e-05, 0.008350464, 0.008805783, 0.08495515, 
    0.01478513, -0.0009923136, 0.01527244, 0.08369312, 0.1623341, 0.1744659, 
    0.09495141, 0.1126324, 0.09017143, 0.0699288, 0.02066709, 0.02133973, 
    0.04603641, 0.01517187, 0.007626208, 0.01422979, 0.03371078, 0.05585367, 
    0.06962583, 0.06965069, 0.06273045, 0.01690438, 0.003037052, 0.0007788419,
  0.04804047, 0.03935513, 0.1477139, 0.1109752, 0.05986081, 0.01363235, 
    0.2073493, 0.0392843, 0.04016027, 0.116599, 0.1019241, 0.1308413, 
    0.1326306, 0.1421963, 0.2257533, 0.2304728, 0.1761791, 0.1369324, 
    0.111089, 0.1325939, 0.2391493, 0.211001, 0.1249897, 0.152473, 0.1620293, 
    0.1496353, 0.07873796, 0.05812534, 0.06398419,
  0.1458153, 0.2098296, 0.1117091, 0.08648658, 0.02705175, 0.1241956, 
    0.2557825, 0.2570705, 0.2240778, 0.2255089, 0.1870833, 0.2117935, 
    0.1517521, 0.2388413, 0.2752613, 0.2863416, 0.2222764, 0.2687863, 
    0.2414482, 0.1873224, 0.1682527, 0.2484578, 0.2006958, 0.3283963, 
    0.296274, 0.2263032, 0.2016196, 0.1779412, 0.1853169,
  0.2642119, 0.255714, 0.1793193, 0.1510469, 0.1376918, 0.1569696, 0.2820856, 
    0.2778884, 0.252021, 0.1729392, 0.1328755, 0.1333341, 0.141467, 
    0.3119976, 0.07498612, 0.2189825, 0.2451694, 0.3944231, 0.2902341, 
    0.07838167, 0.1920254, 0.1814983, 0.3399251, 0.2644609, 0.2292081, 
    0.2173844, 0.2245706, 0.1945724, 0.2951257,
  0.2541001, 0.2307976, 0.28973, 0.2050779, 0.1597099, 0.137378, 0.09760258, 
    0.1144079, 0.1279686, 0.2653751, 0.3194319, 0.2501227, 0.237464, 
    0.3348704, 0.2964255, 0.2033841, 0.3006839, 0.1075771, 0.2334114, 
    0.1443101, 0.1598426, 0.2002022, 0.09787709, 0.05646574, 0.1136434, 
    0.2840276, 0.2127893, 0.2915429, 0.2886517,
  0.2719783, 0.3093336, 0.4303466, 0.3449391, 0.2312439, 0.2176847, 
    0.2828099, 0.2545963, 0.1959156, 0.2153736, 0.1682451, 0.09832077, 
    0.07742134, 0.06340624, 0.1142126, 0.1353648, 0.109121, 0.102635, 
    0.07076029, 0.08946823, 0.1459704, 0.2225224, 0.2387618, 0.2192827, 
    0.1910235, 0.235684, 0.2671266, 0.09730322, 0.364706,
  0.2562161, 0.2474208, 0.2386255, 0.2298302, 0.2210349, 0.2122397, 
    0.2034444, 0.2240391, 0.2289038, 0.2337684, 0.2386331, 0.2434978, 
    0.2483624, 0.2532271, 0.2511455, 0.2646914, 0.2782374, 0.2917834, 
    0.3053294, 0.3188754, 0.3324214, 0.3358026, 0.3261872, 0.3165718, 
    0.3069565, 0.2973411, 0.2877257, 0.2781104, 0.2632523,
  0.1241159, 0.09782873, 0.04910697, 0.05908907, 0.04088603, 0.1130701, 
    0.1100107, 0.09358508, 0.04671053, 0.02397315, 0.02991696, 0.08240125, 
    0.1351675, 0.2411416, 0.3528912, 0.3517396, 0.330273, 0.4040359, 
    0.4018969, 0.5051081, 0.5641004, 0.3762639, 0.2777096, 0.2683557, 
    0.3631105, 0.4167355, 0.4122544, 0.3040366, 0.1396785,
  0.2705712, 0.3656105, 0.2073485, 0.3536453, 0.3910676, 0.1600993, 
    0.3292008, 0.333577, 0.4013692, 0.3490194, 0.3694585, 0.119898, 
    0.1489684, 0.3569598, 0.3760269, 0.4123996, 0.3220961, 0.2960434, 
    0.3103439, 0.2582093, 0.3287519, 0.2722396, 0.3053569, 0.2670468, 
    0.3423101, 0.1894941, 0.1614254, 0.2448412, 0.20355,
  0.3246454, 0.3690901, 0.4238087, 0.3538936, 0.3067684, 0.319244, 0.2804257, 
    0.3844035, 0.3687423, 0.3785163, 0.345787, 0.3263365, 0.2816618, 
    0.3020112, 0.3147182, 0.258965, 0.2889113, 0.2257504, 0.2079944, 
    0.2007399, 0.2133834, 0.2349012, 0.3222047, 0.2445316, 0.1863668, 
    0.3155892, 0.2934506, 0.223107, 0.2203538,
  0.2179789, 0.1822225, 0.2444241, 0.1737163, 0.1820572, 0.238588, 0.2199419, 
    0.2297014, 0.176769, 0.1790663, 0.1868138, 0.2233037, 0.1872409, 
    0.1746571, 0.1005108, 0.1532, 0.2565957, 0.1681813, 0.2245005, 0.2138173, 
    0.2040881, 0.2204287, 0.1642291, 0.1783773, 0.2419196, 0.2176028, 
    0.2400314, 0.2055613, 0.1748487,
  0.1108128, 0.06971522, 0.06314487, 0.1312961, 0.1233445, 0.0983758, 
    0.08967479, 0.1049034, 0.138523, 0.2065634, 0.1526638, 0.07925996, 
    0.0845523, 0.1115649, 0.1312262, 0.1623918, 0.1889108, 0.1277867, 
    0.1942516, 0.1542929, 0.2315111, 0.1045854, 0.1255265, 0.1621384, 
    0.1176943, 0.1377477, 0.1985408, 0.09731372, 0.1273309,
  0.03104589, 0.001978204, 0.0785413, 0.03185532, 0.02414698, 0.05625004, 
    0.04148782, 0.002077999, 0.05899838, 0.06204347, 0.005963771, 0.0191681, 
    0.1206802, 0.05394513, 0.05361443, 0.08071687, 0.08240587, 0.04155514, 
    0.09567602, 0.07241224, 0.1427555, 0.05601966, 0.03405031, 0.005115119, 
    0.09711602, 0.06226542, 0.05700596, 0.08182158, 0.05419013,
  2.002854e-06, 0.02072987, 0.08275471, 0.01761031, 0.03318184, 0.0568784, 
    0.07927405, 0.02911886, 0.1197243, 0.002266008, 0.004259715, 0.02302739, 
    0.02528146, 0.04857346, 0.147345, 0.05251471, 0.05682065, 0.1193916, 
    0.05271567, 0.03313263, 0.03495027, 0.02731172, -4.061287e-06, 
    5.108078e-05, 0.03837705, 0.03394149, 0.03680557, 0.041724, 0.001743667,
  -2.261619e-05, 0.1072775, 0.1751081, 0.1874203, 0.05118973, 0.03174572, 
    0.04341406, 0.08654471, 0.1001032, 0.01690865, 0.06321561, 0.04298169, 
    0.131043, 0.04960636, 0.02062563, 0.03280051, 0.03466644, 0.04304551, 
    0.02426964, 0.01131812, 0.0171178, 0.007596903, 0.0001837714, 0.05558017, 
    0.1102089, 0.04952507, 0.1332945, 0.008131736, 0.0003220534,
  0.008467642, 0.05035201, 0.03388987, 0.1690485, 0.004074109, 0.007860497, 
    0.01124895, 0.01243106, 0.1046602, 0.2191108, 0.1092641, 0.03012262, 
    0.05977745, 0.06457599, 0.03131936, 0.01158159, 0.01844224, 0.01169438, 
    0.007293109, 0.006764224, 0.02941431, 0.02710687, 0.105694, 0.1241625, 
    0.1287261, 0.04338558, 0.02257773, 0.01086466, 0.02689091,
  0.0003808662, -5.282366e-06, -5.173576e-06, 0.2348544, 0.002306823, 
    0.009145579, 0.03504797, 0.02336922, 0.006355233, 0.0091713, 0.03542984, 
    0.01997878, 0.02992898, 0.0858689, 0.09659274, 0.08288543, 0.01216432, 
    0.004102786, 0.04575247, 0.06370448, 0.1289689, 0.01032911, 0.02111971, 
    0.01526104, 0.008663264, 2.171295e-05, 2.678765e-06, 9.250663e-05, 
    0.003547722,
  7.446048e-07, 1.337868e-07, 8.107004e-08, -5.15764e-06, 4.323209e-05, 
    1.576995e-06, 0.007766304, 0.0001386723, 0.0292261, 0.01496475, 
    0.004180118, 0.06210101, 0.04112592, 0.02470909, 0.01380473, 0.01660887, 
    0.02800175, 0.04023102, 3.281287e-05, -4.791633e-05, 1.239798e-05, 
    0.03091686, 0.01304114, 0.04763038, 0.02126103, 0.02033163, 0.000575419, 
    5.025227e-06, 4.522362e-06,
  -1.299598e-05, -4.99943e-05, 0.004502568, 0.007109019, 0.08214559, 
    0.01324352, -0.00335254, 0.01380469, 0.05562477, 0.1581081, 0.1712636, 
    0.1004541, 0.1041312, 0.08511341, 0.07593866, 0.0234491, 0.04405012, 
    0.08525046, 0.001059751, 0.004652938, 0.01615782, 0.03608438, 0.07588415, 
    0.07355075, 0.06629708, 0.05743344, 0.03788072, 0.003875083, 0.001009184,
  0.03677181, 0.03675985, 0.1466589, 0.1135691, 0.03188578, 0.0123169, 
    0.2002203, 0.02721726, 0.03643747, 0.08695546, 0.09890713, 0.1348781, 
    0.1520952, 0.1356084, 0.2240854, 0.2415239, 0.1984511, 0.157505, 
    0.1139361, 0.1391499, 0.2124034, 0.2118904, 0.1556012, 0.1713025, 
    0.1740613, 0.1599974, 0.09212772, 0.06646077, 0.09273821,
  0.1578104, 0.26285, 0.1042453, 0.06710773, 0.04413704, 0.162546, 0.247971, 
    0.2477974, 0.1969589, 0.15881, 0.1639617, 0.2143552, 0.154605, 0.2974952, 
    0.2900439, 0.3659293, 0.2375899, 0.2851528, 0.2368632, 0.1772046, 
    0.1446626, 0.1987862, 0.2425119, 0.3265932, 0.295626, 0.2468372, 
    0.2105232, 0.209249, 0.197654,
  0.2712643, 0.2890731, 0.219483, 0.1355669, 0.1121439, 0.1391629, 0.2528012, 
    0.2668885, 0.2622573, 0.1292923, 0.1521876, 0.1354976, 0.1360828, 
    0.3188973, 0.08193032, 0.1778336, 0.2156396, 0.3900872, 0.2492468, 
    0.08187626, 0.158982, 0.1552607, 0.2785475, 0.263416, 0.2085036, 
    0.216407, 0.2742245, 0.218888, 0.316555,
  0.2717709, 0.2161372, 0.2497713, 0.2106365, 0.1869665, 0.1573485, 
    0.1391133, 0.119417, 0.1339874, 0.2863979, 0.3522578, 0.2765886, 
    0.2234741, 0.2613527, 0.2682252, 0.172908, 0.217486, 0.08911331, 
    0.1410726, 0.1175053, 0.1904363, 0.1498033, 0.08645557, 0.04890336, 
    0.1088555, 0.2968505, 0.2065625, 0.2561798, 0.2646829,
  0.3050238, 0.3009926, 0.4070676, 0.2923517, 0.228706, 0.211789, 0.2732256, 
    0.2823692, 0.2293251, 0.2362458, 0.1786852, 0.08457123, 0.05229579, 
    0.04460747, 0.07456154, 0.1117273, 0.07429207, 0.08483896, 0.09192573, 
    0.1022279, 0.1587634, 0.2387981, 0.2492196, 0.2238992, 0.1904581, 
    0.2486307, 0.2850908, 0.09959764, 0.3396249,
  0.3003374, 0.2942557, 0.288174, 0.2820924, 0.2760107, 0.269929, 0.2638474, 
    0.2967347, 0.3071111, 0.3174874, 0.3278638, 0.3382402, 0.3486166, 
    0.358993, 0.3698438, 0.3775077, 0.3851716, 0.3928355, 0.4004994, 
    0.4081633, 0.4158272, 0.3869256, 0.374967, 0.3630084, 0.3510498, 
    0.3390912, 0.3271325, 0.3151739, 0.3052027,
  0.1187288, 0.1074577, 0.08235607, 0.06622731, 0.07275726, 0.1401535, 
    0.1424669, 0.1406285, 0.07933349, 0.04925855, 0.04244346, 0.1243944, 
    0.190364, 0.2341074, 0.3536809, 0.3328874, 0.3660788, 0.3818895, 
    0.3928165, 0.4650162, 0.5891513, 0.3972763, 0.2584405, 0.2533069, 
    0.3780769, 0.4207706, 0.3835281, 0.2612276, 0.1331264,
  0.2301874, 0.3562208, 0.2089755, 0.3284802, 0.3896208, 0.1625284, 
    0.3585513, 0.3482662, 0.4151465, 0.370714, 0.3566335, 0.1290785, 
    0.1391788, 0.353269, 0.4443009, 0.4520142, 0.3427914, 0.2889598, 
    0.3078441, 0.257919, 0.3056754, 0.2870437, 0.3519464, 0.2967146, 
    0.3874807, 0.1865828, 0.1687798, 0.2597941, 0.1918692,
  0.3166665, 0.3558236, 0.3363879, 0.3383337, 0.3025998, 0.3438282, 
    0.2594714, 0.4231352, 0.3439316, 0.3690326, 0.3476832, 0.3244495, 
    0.3051105, 0.3015006, 0.3379617, 0.2517264, 0.251437, 0.2525543, 
    0.2083491, 0.2094126, 0.2190639, 0.2763503, 0.3193454, 0.2493729, 
    0.2449653, 0.2784383, 0.2873437, 0.2264128, 0.1862128,
  0.2128511, 0.200554, 0.259377, 0.1777638, 0.180564, 0.228879, 0.2477051, 
    0.2373276, 0.2101512, 0.1871098, 0.198239, 0.2125552, 0.1979291, 
    0.1750054, 0.1199728, 0.199792, 0.3014948, 0.2174322, 0.2816505, 
    0.1883957, 0.2200233, 0.2235042, 0.1642709, 0.1735888, 0.2840698, 
    0.2336865, 0.2316543, 0.2108271, 0.2003601,
  0.1170941, 0.08036495, 0.07159425, 0.1552484, 0.1244432, 0.1094873, 
    0.1169931, 0.1155793, 0.1521057, 0.2060979, 0.1646734, 0.1147389, 
    0.08037269, 0.1248057, 0.1445888, 0.1795965, 0.1932685, 0.1312398, 
    0.2069052, 0.1614027, 0.2302351, 0.1166788, 0.1281831, 0.1950625, 
    0.09302304, 0.128461, 0.1941443, 0.09977312, 0.1321955,
  0.03163881, 0.003074436, 0.06902228, 0.04159846, 0.02549168, 0.07302133, 
    0.04942985, 0.006344186, 0.06394006, 0.05551757, 0.005507939, 
    0.004953906, 0.08079559, 0.07046764, 0.07312845, 0.08823971, 0.09937209, 
    0.04883312, 0.0995738, 0.08207557, 0.133895, 0.06029189, 0.05397445, 
    0.004911886, 0.08929671, 0.06520694, 0.0606165, 0.07075347, 0.05823323,
  0.0006494098, 0.005534005, 0.0154521, 0.02122164, 0.02880144, 0.05436908, 
    0.08257412, 0.02428706, 0.1046227, 0.002358235, 0.002087923, 0.005988027, 
    0.02163208, 0.03904616, 0.1542896, 0.05131245, 0.05999494, 0.1350732, 
    0.0478121, 0.05984643, 0.07778454, 0.07050819, 0.0001221274, 
    3.478094e-05, 0.0599976, 0.03909732, 0.04123122, 0.05434472, 0.02415506,
  0.0002797328, 0.08815442, 0.1543266, 0.1966984, 0.04752647, 0.03133534, 
    0.0414783, 0.07827711, 0.09289736, 0.01807346, 0.05854604, 0.04200221, 
    0.1241184, 0.04568652, 0.0194514, 0.02566829, 0.02831198, 0.03448876, 
    0.02274262, 0.01353943, 0.01744248, 0.01025364, 7.547079e-05, 0.05248161, 
    0.105641, 0.06253528, 0.1369043, 0.01249069, 0.001637233,
  0.007227293, 0.05342491, 0.02710566, 0.2157979, 0.005435344, 0.009262872, 
    0.01304793, 0.01200084, 0.113708, 0.2022471, 0.1096423, 0.02875051, 
    0.0539139, 0.05848473, 0.02911019, 0.01198489, 0.0196114, 0.01409577, 
    0.007684393, 0.00790251, 0.03526002, 0.03041914, 0.08378807, 0.1076865, 
    0.1257633, 0.03983644, 0.0230928, 0.01324657, 0.02564013,
  0.0001901797, -3.111358e-06, -1.765443e-06, 0.1660744, 0.002675385, 
    0.01222914, 0.03053158, 0.01700675, 0.007136603, 0.01487885, 0.04601274, 
    0.02751796, 0.03280434, 0.07694148, 0.0872542, 0.07093709, 0.01608292, 
    0.008226127, 0.05290801, 0.06597355, 0.1197958, 0.01222252, 0.03791853, 
    0.008814919, 0.01563769, 0.0003162401, 1.397194e-06, 2.164857e-05, 
    0.002320428,
  7.033308e-07, 7.910075e-08, 6.360068e-08, -3.398856e-06, 1.740001e-05, 
    1.360554e-07, 0.0004855072, 0.0001770819, 0.01093246, 0.007928241, 
    0.01637724, 0.0826512, 0.06435102, 0.04091758, 0.04163212, 0.04813483, 
    0.02788338, 0.04547511, 0.002636764, -1.010368e-05, 8.734659e-06, 
    0.04354753, 0.01792919, 0.04289955, 0.02123357, 0.03870358, 0.0110228, 
    2.365358e-06, 2.013464e-06,
  3.3396e-07, -2.978946e-05, 0.00214561, 0.003735109, 0.07968245, 0.01143335, 
    -0.002889974, 0.008851749, 0.04505282, 0.1493501, 0.1724108, 0.1105001, 
    0.1100938, 0.08951534, 0.07260332, 0.04611237, 0.05923025, 0.1021081, 
    0.001401882, 0.01357063, 0.01842302, 0.04571686, 0.07072075, 0.08319777, 
    0.07223749, 0.04558904, 0.04522814, 0.006502082, 0.002692183,
  0.0221907, 0.03862967, 0.1452888, 0.1098984, 0.02423516, 0.005147101, 
    0.1857562, 0.03011135, 0.03103542, 0.08268397, 0.1042574, 0.1205302, 
    0.1485499, 0.1377426, 0.2433367, 0.2524073, 0.2009818, 0.1560292, 
    0.1592602, 0.1285797, 0.1840126, 0.2115282, 0.1725336, 0.1785284, 
    0.1988198, 0.165493, 0.1127735, 0.08125168, 0.08670171,
  0.1625762, 0.260795, 0.1148324, 0.06289182, 0.044687, 0.14738, 0.207732, 
    0.2507106, 0.172274, 0.1214589, 0.1368628, 0.2036109, 0.1302743, 
    0.3153393, 0.286734, 0.3630011, 0.2752144, 0.2732937, 0.2317959, 
    0.1854095, 0.124585, 0.1364764, 0.1998361, 0.3202454, 0.2785605, 
    0.2516429, 0.2259222, 0.2127204, 0.2115,
  0.2947408, 0.2970923, 0.2349925, 0.1575644, 0.1297395, 0.1692121, 
    0.1743177, 0.2670664, 0.262155, 0.138448, 0.1848192, 0.1506154, 
    0.1220864, 0.3264796, 0.1010216, 0.1475626, 0.1925305, 0.3797944, 
    0.1911258, 0.08072537, 0.1467776, 0.1379959, 0.2489003, 0.2601508, 
    0.199523, 0.1860834, 0.2948616, 0.2650535, 0.3270166,
  0.2748975, 0.2609854, 0.2303907, 0.1893243, 0.1734068, 0.1710778, 
    0.1246315, 0.1331825, 0.1407052, 0.303432, 0.3062766, 0.2280871, 
    0.2090687, 0.2666788, 0.2249855, 0.1418114, 0.1675375, 0.07268118, 
    0.04430435, 0.04651983, 0.1290837, 0.1110184, 0.09076496, 0.07717966, 
    0.1161416, 0.3096277, 0.193895, 0.2082658, 0.2701569,
  0.2921016, 0.2172035, 0.3643517, 0.2966233, 0.2372986, 0.1920085, 0.237374, 
    0.2318059, 0.1854654, 0.2538921, 0.2107706, 0.09564906, 0.04903848, 
    0.04853868, 0.05467185, 0.08448982, 0.03433287, 0.03991424, 0.0559436, 
    0.06084103, 0.1167096, 0.1850877, 0.25247, 0.231501, 0.1936923, 
    0.2762624, 0.3034773, 0.1140499, 0.3229428,
  0.3328915, 0.3284591, 0.3240268, 0.3195945, 0.3151622, 0.3107299, 
    0.3062975, 0.3506283, 0.3644005, 0.3781726, 0.3919448, 0.405717, 
    0.4194891, 0.4332613, 0.4404404, 0.4440921, 0.4477438, 0.4513955, 
    0.4550472, 0.458699, 0.4623507, 0.4246754, 0.4116839, 0.3986923, 
    0.3857008, 0.3727093, 0.3597177, 0.3467262, 0.3364373,
  0.1172309, 0.1252135, 0.1149773, 0.077517, 0.1032816, 0.1636969, 0.152192, 
    0.1662359, 0.0948798, 0.05835759, 0.08634517, 0.1409658, 0.2160132, 
    0.2053128, 0.2725137, 0.3535245, 0.4067131, 0.3768077, 0.3566764, 
    0.4629675, 0.6203037, 0.3981185, 0.2409669, 0.2782625, 0.3857657, 
    0.4315102, 0.375361, 0.217299, 0.1534753,
  0.3176701, 0.3086618, 0.2129756, 0.3031251, 0.3353792, 0.1363724, 
    0.3620686, 0.3835113, 0.4238371, 0.3691548, 0.3423027, 0.1066879, 
    0.1446829, 0.3831142, 0.5349118, 0.4446278, 0.4014514, 0.3245799, 
    0.3718462, 0.3116693, 0.3225894, 0.3098081, 0.3623979, 0.3034977, 
    0.3421018, 0.3093789, 0.1654681, 0.2997524, 0.2028177,
  0.4077412, 0.4006351, 0.3089169, 0.3549631, 0.3194332, 0.3306739, 
    0.3290105, 0.4602134, 0.3883362, 0.3950036, 0.3929125, 0.3435021, 
    0.3580706, 0.3169379, 0.3495308, 0.2959216, 0.3100822, 0.2858858, 
    0.2497243, 0.2684168, 0.2392898, 0.3586826, 0.3253179, 0.3453719, 
    0.3472539, 0.298361, 0.293873, 0.2274964, 0.2184737,
  0.2463512, 0.2314498, 0.3112165, 0.206994, 0.2091318, 0.2454451, 0.2883002, 
    0.2928168, 0.2424981, 0.219872, 0.2210227, 0.2645603, 0.2502428, 
    0.2257674, 0.1734106, 0.2353235, 0.3488763, 0.2705075, 0.347836, 
    0.2465093, 0.25111, 0.2302549, 0.1978012, 0.1733912, 0.2793082, 
    0.2331487, 0.2579425, 0.2392578, 0.2552179,
  0.1399176, 0.1061709, 0.1039371, 0.2061607, 0.1457357, 0.1647864, 
    0.1425368, 0.1569207, 0.1774629, 0.2418131, 0.1714791, 0.1214226, 
    0.1055422, 0.144917, 0.1755967, 0.2033301, 0.2073243, 0.1420074, 
    0.2419285, 0.1829309, 0.2334066, 0.1327672, 0.1800714, 0.207699, 
    0.07089883, 0.1392598, 0.1776147, 0.1233965, 0.1597055,
  0.04115435, 0.01574742, 0.04737271, 0.05838053, 0.03035884, 0.0835173, 
    0.06284337, 0.03800248, 0.07860602, 0.07262351, 0.01632238, 0.0001807874, 
    0.04371227, 0.1057049, 0.1108059, 0.1473562, 0.1051994, 0.06649089, 
    0.1197645, 0.09128388, 0.1368393, 0.07470764, 0.08664212, 0.004096061, 
    0.07480031, 0.07273626, 0.08670476, 0.06718203, 0.06608511,
  0.00552281, 0.004924721, 0.004397388, 0.01963668, 0.0298251, 0.06048235, 
    0.09976197, 0.03877002, 0.11614, 0.002281304, 0.001326291, 0.003700286, 
    0.02253486, 0.03700778, 0.1065965, 0.05395596, 0.07512863, 0.1324963, 
    0.03762832, 0.05233816, 0.06607224, 0.0943405, 0.01678801, 1.518424e-05, 
    0.07544117, 0.05156132, 0.03066892, 0.07601978, 0.08503109,
  0.008341751, 0.07293046, 0.1338329, 0.184038, 0.04006079, 0.02938584, 
    0.03956846, 0.07059146, 0.07780718, 0.01786108, 0.04712936, 0.03712191, 
    0.1127008, 0.03755501, 0.01827114, 0.02138252, 0.02263097, 0.02833229, 
    0.02243285, 0.01484718, 0.01999842, 0.01618655, 0.0001285183, 0.04785956, 
    0.09858654, 0.05095244, 0.1146166, 0.01876832, 0.005872508,
  0.008563805, 0.051032, 0.02179702, 0.1474772, 0.008648471, 0.01253187, 
    0.01499544, 0.01138995, 0.1144239, 0.1888493, 0.09508628, 0.02394872, 
    0.04668789, 0.04564065, 0.02715172, 0.01289686, 0.01917441, 0.01491525, 
    0.008032375, 0.007401139, 0.03454051, 0.03074053, 0.06193107, 0.09708012, 
    0.1177435, 0.03594364, 0.02306902, 0.01456897, 0.02282581,
  9.557931e-05, -1.242869e-06, -6.538169e-07, 0.114691, 0.002779408, 
    0.01989685, 0.02874945, 0.01802793, 0.009475904, 0.01886976, 0.05674633, 
    0.02622266, 0.035441, 0.06601743, 0.08199567, 0.06055452, 0.02442447, 
    0.01442543, 0.0595785, 0.07257707, 0.1025108, 0.01464197, 0.04453434, 
    0.01116878, 0.02708951, 0.005643754, 2.132129e-05, 5.947541e-07, 
    0.001523318,
  6.420598e-07, 4.998884e-08, 2.188643e-08, -1.601578e-06, 2.736739e-06, 
    2.0796e-07, 0.0004065103, 0.0002056719, 0.004475655, 0.01644842, 
    0.02299932, 0.1026186, 0.06610816, 0.03440921, 0.04067378, 0.07666259, 
    0.04785435, 0.09111042, 0.01868282, 0.0003595032, 3.900498e-06, 
    0.05748582, 0.0291526, 0.03054164, 0.02144199, 0.0336678, 0.06186152, 
    -4.242177e-06, 1.191843e-06,
  3.823006e-07, 8.516834e-06, 0.004200801, 0.002523496, 0.07131317, 
    0.0102012, -0.002376694, 0.004667224, 0.03408445, 0.158939, 0.1706295, 
    0.1717803, 0.1534555, 0.133517, 0.07702168, 0.08598469, 0.0709006, 
    0.1103198, 0.01216808, 0.02380626, 0.01586396, 0.07353207, 0.06640708, 
    0.1113693, 0.09369057, 0.05437722, 0.05610932, 0.02383729, 0.002558168,
  0.01147524, 0.03828357, 0.1270258, 0.1073578, 0.01414436, 0.002413842, 
    0.1697304, 0.02405104, 0.02656643, 0.07669514, 0.1197403, 0.1099822, 
    0.1492306, 0.1737794, 0.2578099, 0.2878683, 0.2201822, 0.175293, 
    0.1914496, 0.1522633, 0.1856985, 0.221568, 0.1928044, 0.1795481, 
    0.2187438, 0.1777163, 0.124195, 0.1073167, 0.08050074,
  0.1531396, 0.2696955, 0.1162481, 0.05764805, 0.05227004, 0.15241, 
    0.1926348, 0.2381693, 0.1450497, 0.08320918, 0.1053298, 0.2052805, 
    0.1505904, 0.3448414, 0.3157853, 0.3815973, 0.2776484, 0.2760929, 
    0.2455223, 0.2346522, 0.1148727, 0.1311857, 0.192304, 0.3204227, 
    0.295952, 0.2887517, 0.2615177, 0.2488268, 0.2200613,
  0.2764944, 0.3283307, 0.2313617, 0.2037931, 0.133433, 0.1547527, 0.1914422, 
    0.2682289, 0.206462, 0.156499, 0.1699855, 0.1987274, 0.1003283, 
    0.3071726, 0.2135556, 0.1804101, 0.2759762, 0.3755035, 0.2398833, 
    0.08985136, 0.1254077, 0.1541723, 0.2228454, 0.2744413, 0.2352328, 
    0.1690947, 0.350943, 0.3109146, 0.3462155,
  0.3185399, 0.3227622, 0.236336, 0.227655, 0.2676709, 0.2349821, 0.1718615, 
    0.1623701, 0.1528472, 0.331051, 0.2613222, 0.2115945, 0.2305324, 
    0.2527766, 0.233551, 0.1620839, 0.1806762, 0.06137029, 0.03801968, 
    0.04187258, 0.09828457, 0.1085414, 0.05385705, 0.1004181, 0.08614833, 
    0.3197277, 0.1678929, 0.1675808, 0.4144922,
  0.2701684, 0.2667931, 0.3907854, 0.2780297, 0.278027, 0.2407357, 0.2874679, 
    0.239752, 0.2227553, 0.2153047, 0.3000819, 0.1369674, 0.05339229, 
    0.05302884, 0.05972192, 0.08525708, 0.02964241, 0.03244774, 0.03587664, 
    0.02843269, 0.0842841, 0.1234575, 0.2326093, 0.2293202, 0.1749421, 
    0.2991175, 0.2970263, 0.1273635, 0.3343173,
  0.3681359, 0.3673311, 0.3665263, 0.3657216, 0.3649168, 0.364112, 0.3633072, 
    0.3797287, 0.3941486, 0.4085687, 0.4229886, 0.4374086, 0.4518286, 
    0.4662485, 0.4629462, 0.4615766, 0.4602069, 0.4588373, 0.4574676, 
    0.456098, 0.4547284, 0.4400899, 0.4278443, 0.4155988, 0.4033532, 
    0.3911076, 0.3788621, 0.3666165, 0.3687798,
  0.1230053, 0.1438777, 0.1658755, 0.09019867, 0.1243777, 0.1831322, 
    0.1710857, 0.2162101, 0.1213265, 0.06348587, 0.14676, 0.1688931, 
    0.2190827, 0.168832, 0.2549674, 0.3381093, 0.3710027, 0.4530183, 
    0.3778999, 0.450872, 0.6399788, 0.4470937, 0.2555293, 0.3001754, 
    0.3639278, 0.4484664, 0.3572499, 0.2412312, 0.1617904,
  0.3473516, 0.3723748, 0.2368429, 0.2654744, 0.3073051, 0.1562015, 
    0.3302549, 0.4389026, 0.4192573, 0.365621, 0.3366671, 0.09142157, 
    0.1699399, 0.3791597, 0.5871518, 0.4364353, 0.4682948, 0.4148442, 
    0.454247, 0.4123474, 0.3795299, 0.3510824, 0.3427078, 0.335264, 
    0.3341081, 0.3153762, 0.2155732, 0.3871923, 0.2005158,
  0.4810467, 0.4303166, 0.355205, 0.3543347, 0.3235589, 0.300733, 0.3746413, 
    0.4547074, 0.4235511, 0.4638378, 0.4048218, 0.3875513, 0.3877863, 
    0.3685223, 0.351624, 0.3463324, 0.4116276, 0.2867891, 0.2864662, 
    0.3275377, 0.3240687, 0.4331399, 0.3539107, 0.3930577, 0.3837281, 
    0.4535703, 0.3197651, 0.3127446, 0.3167838,
  0.2713941, 0.2933666, 0.3616256, 0.262251, 0.2437484, 0.3051923, 0.3250754, 
    0.3060196, 0.2571942, 0.2658608, 0.2600713, 0.3070634, 0.2910048, 
    0.3180172, 0.1931298, 0.2794198, 0.3548535, 0.2926868, 0.3500799, 
    0.3103723, 0.2887407, 0.3372376, 0.296387, 0.1817206, 0.3047458, 
    0.2354397, 0.2460654, 0.2632747, 0.2509434,
  0.1684631, 0.1715734, 0.1687156, 0.2236923, 0.2017664, 0.1802837, 
    0.1651208, 0.2026427, 0.2645587, 0.3143765, 0.2086375, 0.1809803, 
    0.1061395, 0.1747221, 0.1961063, 0.2051455, 0.228771, 0.2026488, 
    0.2331938, 0.2049579, 0.2718801, 0.1579592, 0.2471621, 0.2424621, 
    0.07250147, 0.1215134, 0.1622668, 0.1150133, 0.2011424,
  0.09447844, 0.01140751, 0.03665562, 0.06465857, 0.04784591, 0.09723371, 
    0.06679857, 0.1526055, 0.1705128, 0.1192628, 0.02189129, -2.473858e-05, 
    0.02767282, 0.1471962, 0.09284286, 0.1560655, 0.1304917, 0.1399557, 
    0.2152647, 0.1451227, 0.1511221, 0.08953611, 0.1218981, 0.003706869, 
    0.07765411, 0.0899408, 0.1412046, 0.06296195, 0.07850593,
  0.03215609, 0.005018935, 0.0008132788, 0.02615266, 0.04259375, 0.07648382, 
    0.08953533, 0.05436233, 0.1554003, 0.002468449, 0.0004516183, 
    0.002820665, 0.03822585, 0.04177006, 0.1133886, 0.05464097, 0.1185407, 
    0.1338267, 0.03675616, 0.04274185, 0.04847022, 0.1015391, 0.08395769, 
    2.168697e-05, 0.07386316, 0.07592223, 0.03254898, 0.05113291, 0.0988988,
  0.01300215, 0.0565246, 0.1104885, 0.1675873, 0.03840938, 0.03105661, 
    0.03845115, 0.0597489, 0.06046893, 0.02105366, 0.04260724, 0.04933963, 
    0.110954, 0.03403061, 0.01950262, 0.02295, 0.02132424, 0.02604014, 
    0.02853278, 0.02261633, 0.02175715, 0.02805018, 0.002040575, 0.04391749, 
    0.0923959, 0.0325949, 0.09354563, 0.03171561, 0.02257635,
  0.01301224, 0.04487961, 0.01844461, 0.08670318, 0.01644416, 0.01851936, 
    0.01959295, 0.01328497, 0.1026743, 0.1738182, 0.07397139, 0.02353331, 
    0.04071941, 0.04275858, 0.02718242, 0.01656307, 0.01950455, 0.01603686, 
    0.009129145, 0.007664464, 0.03168917, 0.03191479, 0.04328665, 0.08402687, 
    0.1119701, 0.03560423, 0.02375173, 0.01459004, 0.02395175,
  3.009074e-05, -2.172527e-07, -3.318747e-07, 0.07049582, 0.006200967, 
    0.02890687, 0.02969275, 0.02254522, 0.0165067, 0.03245363, 0.05527083, 
    0.02438598, 0.03918822, 0.0532607, 0.07845652, 0.0521451, 0.04029274, 
    0.0293761, 0.06458067, 0.07744364, 0.0948179, 0.02020878, 0.05130554, 
    0.0184985, 0.03786953, 0.02652527, 0.003287006, 4.389589e-08, 0.000984531,
  5.60738e-07, 3.452985e-08, 5.256129e-09, 3.904601e-06, 5.376486e-07, 
    -6.155271e-06, 0.000249644, 3.095936e-05, 0.001286767, 0.04368671, 
    0.03874519, 0.1073761, 0.05866507, 0.03061742, 0.0333188, 0.08111843, 
    0.08268392, 0.1318843, 0.07008931, 0.006564035, 1.588889e-06, 0.06616215, 
    0.06346049, 0.05298178, 0.02975327, 0.04658695, 0.06991977, 0.001518482, 
    6.552567e-07,
  3.26158e-07, 1.945383e-06, 0.002643891, 0.00241408, 0.0598092, 0.00465246, 
    -0.002030902, 0.0009682513, 0.02513949, 0.1836817, 0.1967, 0.1716691, 
    0.1945265, 0.1614904, 0.155075, 0.1569326, 0.1222646, 0.143252, 
    0.08153795, 0.03599319, 0.01585947, 0.1051393, 0.09483316, 0.1646996, 
    0.1369408, 0.08920665, 0.07251208, 0.05028249, 0.003045183,
  0.007198332, 0.03590687, 0.09185518, 0.1230889, 0.009671867, 0.003189095, 
    0.1519902, 0.01844495, 0.02334125, 0.07856791, 0.1321056, 0.09915014, 
    0.2187132, 0.2164332, 0.2916402, 0.3089005, 0.2364797, 0.2359667, 
    0.306134, 0.1653271, 0.1496456, 0.2332987, 0.1905937, 0.1544378, 
    0.2546113, 0.1751247, 0.153487, 0.1537744, 0.08496224,
  0.1469426, 0.2984532, 0.09831439, 0.0914505, 0.04116172, 0.1595043, 
    0.2205986, 0.2274744, 0.1189495, 0.06011587, 0.08949423, 0.1986759, 
    0.1800559, 0.4142615, 0.4168144, 0.4304809, 0.2884953, 0.3039447, 
    0.2880739, 0.2525521, 0.1065376, 0.1162077, 0.2040384, 0.3344364, 
    0.353854, 0.2842987, 0.3178013, 0.264473, 0.2172383,
  0.3021986, 0.3627427, 0.2027524, 0.1559488, 0.1525365, 0.1683761, 
    0.2141719, 0.2049049, 0.173688, 0.09383107, 0.1901345, 0.2048199, 
    0.08278216, 0.2747314, 0.3127359, 0.2278829, 0.3134808, 0.380776, 
    0.2620382, 0.04333872, 0.1182905, 0.1359217, 0.2067282, 0.3246313, 
    0.2874325, 0.168898, 0.2966847, 0.3660159, 0.3625473,
  0.3488726, 0.3347057, 0.2627788, 0.2797538, 0.3394329, 0.1879426, 
    0.2275006, 0.1885317, 0.1620798, 0.3538876, 0.26651, 0.2842714, 
    0.2177769, 0.218067, 0.2315865, 0.145852, 0.1770268, 0.04843588, 
    0.0290542, 0.03764094, 0.1084079, 0.0989329, 0.03588046, 0.1006756, 
    0.09530782, 0.3293796, 0.1537355, 0.141857, 0.4835211,
  0.336309, 0.3341812, 0.3729744, 0.2831566, 0.2362385, 0.2545013, 0.2619533, 
    0.1986323, 0.1884566, 0.2321989, 0.1869209, 0.1111037, 0.08005654, 
    0.07417095, 0.08449542, 0.07534149, 0.04865788, 0.05296613, 0.05622848, 
    0.04725666, 0.07584578, 0.1394377, 0.216339, 0.2177814, 0.1614107, 
    0.2957857, 0.2816522, 0.153614, 0.311287,
  0.400963, 0.403028, 0.4050929, 0.4071579, 0.4092228, 0.4112878, 0.4133527, 
    0.4218818, 0.4350815, 0.4482812, 0.4614809, 0.4746806, 0.4878803, 
    0.50108, 0.4833129, 0.4781638, 0.4730147, 0.4678656, 0.4627165, 
    0.4575675, 0.4524184, 0.4474204, 0.4373049, 0.4271894, 0.4170738, 
    0.4069583, 0.3968427, 0.3867272, 0.3993111,
  0.1305353, 0.1695595, 0.2032683, 0.1436257, 0.1437864, 0.2033997, 
    0.2082612, 0.2547526, 0.1492471, 0.06679299, 0.1770974, 0.2048776, 
    0.2412588, 0.1293559, 0.2016321, 0.4078169, 0.3669179, 0.4709224, 
    0.4161581, 0.4484441, 0.6635427, 0.4895991, 0.2831874, 0.3027278, 
    0.3565431, 0.4531414, 0.3318759, 0.2421284, 0.1567074,
  0.3320605, 0.3325208, 0.2049456, 0.2181089, 0.266455, 0.1858193, 0.2874797, 
    0.4361016, 0.4038728, 0.3552133, 0.3405902, 0.09809235, 0.1532621, 
    0.3944522, 0.5901346, 0.443017, 0.4430845, 0.5161629, 0.4906215, 
    0.4190578, 0.4450354, 0.4132887, 0.3256924, 0.3365227, 0.3417079, 
    0.3249222, 0.2242141, 0.4561282, 0.2215899,
  0.4875347, 0.4214141, 0.3405522, 0.361153, 0.3189859, 0.3056203, 0.3529531, 
    0.426193, 0.4650138, 0.4267234, 0.3949965, 0.4390254, 0.4790892, 
    0.4085537, 0.3237311, 0.3611077, 0.3927987, 0.3678766, 0.298866, 
    0.3552298, 0.3563446, 0.5283667, 0.4746964, 0.3615909, 0.4144726, 
    0.4954965, 0.4411769, 0.3682307, 0.418553,
  0.3002555, 0.3104476, 0.3315676, 0.2942747, 0.2574813, 0.3166344, 
    0.3476885, 0.3099466, 0.2664362, 0.2690842, 0.2666923, 0.2868243, 
    0.2849112, 0.3014245, 0.2160696, 0.2902645, 0.3486785, 0.2564475, 
    0.3313386, 0.3311916, 0.3923364, 0.3817981, 0.3295569, 0.1875479, 
    0.2724366, 0.2363925, 0.2799031, 0.2617366, 0.2509827,
  0.2377028, 0.2157363, 0.2321986, 0.2376007, 0.2300876, 0.243258, 0.2167376, 
    0.2463435, 0.2650847, 0.3219936, 0.2021529, 0.1730127, 0.07965507, 
    0.2143603, 0.2345731, 0.1929615, 0.2104453, 0.2082167, 0.1981924, 
    0.2055426, 0.2754948, 0.1867737, 0.263428, 0.2930721, 0.04633377, 
    0.07875384, 0.1344399, 0.113193, 0.2334494,
  0.1792142, 0.04243279, 0.04015446, 0.07917897, 0.05235574, 0.136349, 
    0.07700583, 0.1586335, 0.249207, 0.1168871, 0.01521566, -2.173841e-05, 
    0.02832628, 0.1267396, 0.1167416, 0.09769166, 0.1272074, 0.09393159, 
    0.1939109, 0.119434, 0.183961, 0.1057422, 0.1287573, 0.004789217, 
    0.08762423, 0.1006659, 0.1620529, 0.09120397, 0.1022545,
  0.1768157, 0.001347473, 0.0004380976, 0.03351569, 0.08794513, 0.0798405, 
    0.08572047, 0.09341342, 0.1720351, 0.002638653, 0.000129848, 0.001490073, 
    0.06729268, 0.06591052, 0.1022996, 0.04758383, 0.1125739, 0.1489286, 
    0.04821286, 0.05837106, 0.05574959, 0.09024435, 0.141892, 0.0001157876, 
    0.06233375, 0.07822189, 0.04461749, 0.05029839, 0.1549541,
  0.02614252, 0.0503745, 0.07570051, 0.1767298, 0.06485027, 0.04157875, 
    0.04367021, 0.05158506, 0.05806776, 0.02835179, 0.0507487, 0.05978027, 
    0.1015345, 0.03702729, 0.02366181, 0.02745136, 0.02647805, 0.02936104, 
    0.04795431, 0.07218777, 0.04297896, 0.08510462, 0.02519225, 0.03938638, 
    0.08420694, 0.01466156, 0.1005155, 0.09085343, 0.09162336,
  0.02247793, 0.03566656, 0.0127089, 0.04419957, 0.04595669, 0.0479595, 
    0.04072456, 0.01874927, 0.08430427, 0.1490761, 0.06134764, 0.02644687, 
    0.04021662, 0.04585168, 0.03596815, 0.0259665, 0.02342005, 0.02153591, 
    0.01493083, 0.009487321, 0.03115857, 0.03707421, 0.02960255, 0.06434025, 
    0.09264816, 0.03814455, 0.02867664, 0.0192528, 0.02974221,
  2.013801e-06, 2.683207e-07, -7.964947e-08, 0.04287839, 0.01202696, 
    0.2007178, 0.03734908, 0.0338838, 0.02411512, 0.06582797, 0.05930285, 
    0.03132547, 0.04155014, 0.05519143, 0.0838956, 0.06034433, 0.07074822, 
    0.0552621, 0.08833615, 0.1059144, 0.1031651, 0.09469331, 0.04418448, 
    0.02520623, 0.06664208, 0.09795534, 0.03613197, -1.84741e-06, 0.0004677666,
  4.500315e-07, 2.714717e-08, 1.40899e-09, -2.895302e-07, -1.940485e-06, 
    0.000161386, 2.281068e-05, -1.835917e-05, 0.0004730343, 0.09933737, 
    0.05716027, 0.1185708, 0.06239776, 0.04026869, 0.05291592, 0.1008306, 
    0.06040855, 0.1567913, 0.1828541, 0.02003578, 3.093978e-06, 0.07269572, 
    0.1057462, 0.062871, 0.07962537, 0.08762777, 0.1150215, 0.08227795, 
    4.484278e-07,
  3.197044e-07, 9.00681e-07, 0.002566891, 0.002755297, 0.05207329, 0.0030295, 
    -0.001699186, -6.882134e-05, 0.02051031, 0.1788995, 0.1981951, 0.226476, 
    0.2395347, 0.1367719, 0.1517847, 0.1496237, 0.1568833, 0.1706184, 
    0.2536774, 0.06545756, 0.01374982, 0.143107, 0.08276489, 0.130442, 
    0.1707952, 0.114197, 0.1423295, 0.2028273, 0.01342969,
  0.005260601, 0.01804647, 0.05577976, 0.1254599, 0.001340376, 0.002494024, 
    0.1310111, 0.01520208, 0.02127853, 0.07073054, 0.1382505, 0.09606022, 
    0.241618, 0.211492, 0.2751062, 0.2747237, 0.2260481, 0.267109, 0.325811, 
    0.1572396, 0.1273076, 0.2490723, 0.1492571, 0.1419357, 0.2451771, 
    0.185738, 0.2017769, 0.1724286, 0.07868004,
  0.1732936, 0.262352, 0.08304191, 0.02160808, 0.04022384, 0.1699248, 
    0.2064444, 0.2373639, 0.09824518, 0.0413042, 0.08904283, 0.1873882, 
    0.1744439, 0.3666111, 0.3661848, 0.3712791, 0.3001783, 0.3302533, 
    0.3150752, 0.2458301, 0.09229336, 0.1312082, 0.206211, 0.3632858, 
    0.4221218, 0.4216972, 0.3648365, 0.2272428, 0.2131679,
  0.2988843, 0.358481, 0.2014234, 0.130086, 0.1124404, 0.1629352, 0.2355446, 
    0.171669, 0.131628, 0.06727803, 0.1838377, 0.1823269, 0.0512393, 
    0.2505143, 0.3494941, 0.2399035, 0.3086168, 0.4026246, 0.1826473, 
    0.02634905, 0.09434927, 0.1273636, 0.2428242, 0.3137276, 0.4325703, 
    0.1367009, 0.1908972, 0.2869077, 0.3407937,
  0.332055, 0.2788523, 0.2561016, 0.235476, 0.2968394, 0.2230303, 0.2027036, 
    0.167151, 0.1576324, 0.3694616, 0.2809038, 0.321154, 0.2516298, 
    0.2944922, 0.2176249, 0.1771252, 0.2012701, 0.04258877, 0.02961937, 
    0.05761596, 0.09152416, 0.09413887, 0.05460446, 0.1127638, 0.07484145, 
    0.3363247, 0.1419287, 0.1038703, 0.4200908,
  0.3415317, 0.3378414, 0.3803023, 0.304823, 0.2613922, 0.2444774, 0.2548916, 
    0.2139256, 0.2270971, 0.2357941, 0.1510488, 0.07305305, 0.1263034, 
    0.07950908, 0.09947015, 0.09306293, 0.06426531, 0.07494411, 0.06497858, 
    0.07685214, 0.1168074, 0.1781138, 0.2035816, 0.2158875, 0.1623821, 
    0.2726505, 0.2556635, 0.1572527, 0.3121437,
  0.4257114, 0.4279828, 0.4302543, 0.4325257, 0.4347971, 0.4370686, 0.43934, 
    0.4300043, 0.441374, 0.4527438, 0.4641136, 0.4754834, 0.4868532, 
    0.498223, 0.4882156, 0.4812576, 0.4742995, 0.4673415, 0.4603834, 
    0.4534253, 0.4464673, 0.4462695, 0.4395864, 0.4329032, 0.42622, 
    0.4195369, 0.4128537, 0.4061705, 0.4238943,
  0.1477159, 0.1868984, 0.2621172, 0.2223468, 0.170968, 0.2293777, 0.2517152, 
    0.2940844, 0.1523587, 0.1230008, 0.2247009, 0.2274145, 0.2898166, 
    0.1017976, 0.163688, 0.3770165, 0.3440557, 0.4820373, 0.4326555, 
    0.415615, 0.6926585, 0.5406148, 0.3152727, 0.2486875, 0.3799488, 
    0.4812111, 0.3237949, 0.2370175, 0.1639252,
  0.3169163, 0.2591903, 0.1763823, 0.1531464, 0.2229622, 0.2144614, 
    0.2148325, 0.4198264, 0.3935608, 0.3468335, 0.3333027, 0.08879979, 
    0.1552803, 0.3198785, 0.4896753, 0.4379825, 0.3936699, 0.4862703, 
    0.4841138, 0.4051269, 0.4760063, 0.4437656, 0.3817935, 0.3566667, 
    0.3407023, 0.3162458, 0.3725047, 0.4542035, 0.2164542,
  0.4308454, 0.3649477, 0.3272439, 0.3551678, 0.3127238, 0.3043157, 
    0.3320487, 0.3925228, 0.4156374, 0.4210852, 0.384269, 0.441478, 
    0.5246547, 0.4152258, 0.3233014, 0.3724217, 0.4064383, 0.4498438, 
    0.4060124, 0.3824078, 0.373217, 0.4822209, 0.4706781, 0.3537574, 
    0.3606382, 0.525521, 0.4980045, 0.3373321, 0.3551564,
  0.3513726, 0.3169263, 0.3168969, 0.3103623, 0.2758858, 0.2920556, 
    0.3488477, 0.3066386, 0.2648174, 0.2711753, 0.2816913, 0.3183995, 
    0.3273686, 0.2153463, 0.1987997, 0.2580768, 0.3417418, 0.2188666, 
    0.2748851, 0.3226296, 0.3887552, 0.3644156, 0.2888947, 0.1904858, 
    0.1983686, 0.2350748, 0.2507642, 0.2759879, 0.309309,
  0.3065786, 0.2448507, 0.2626639, 0.192572, 0.1925108, 0.1853033, 0.2067515, 
    0.2808957, 0.2504731, 0.2766839, 0.2098076, 0.226748, 0.04258315, 
    0.1925691, 0.3040926, 0.1338901, 0.2373278, 0.1978748, 0.1810587, 
    0.2482612, 0.2934192, 0.2847142, 0.2581121, 0.3498718, 0.05351498, 
    0.0564747, 0.1292605, 0.1655214, 0.2676726,
  0.2202115, 0.07724395, 0.01073465, 0.06621113, 0.09019545, 0.1460089, 
    0.08222792, 0.2008599, 0.187714, 0.07951995, 0.009305784, -2.370516e-05, 
    0.02140165, 0.07586299, 0.07814164, 0.09850469, 0.0913262, 0.06885344, 
    0.1337015, 0.1286137, 0.1918934, 0.1027915, 0.1072285, 0.01066613, 
    0.08845764, 0.08676044, 0.1688414, 0.1129271, 0.1741053,
  0.2774065, 0.0001539104, 0.0001584673, 0.06232874, 0.06215102, 0.08237547, 
    0.06817351, 0.08149075, 0.1676374, 0.01929635, 4.57559e-05, 0.0005825654, 
    0.03580221, 0.07723824, 0.09360972, 0.04450024, 0.0702737, 0.1263763, 
    0.04334193, 0.03594183, 0.04135538, 0.09070754, 0.2492813, 0.0004271555, 
    0.05459379, 0.07765155, 0.05137678, 0.06805322, 0.1297454,
  0.2429053, 0.0455577, 0.04973257, 0.1338813, 0.08859102, 0.09050153, 
    0.1009218, 0.05473595, 0.08344612, 0.04440621, 0.05682544, 0.04384946, 
    0.09763514, 0.04136325, 0.03131789, 0.08297177, 0.1505791, 0.05921642, 
    0.07027199, 0.09234388, 0.08718999, 0.1165595, 0.2224332, 0.02477595, 
    0.05850572, 0.004013975, 0.1091926, 0.10858, 0.2831551,
  0.04346335, 0.01893778, 0.006368563, 0.02077989, 0.2451181, 0.1808624, 
    0.1216688, 0.03634394, 0.05684998, 0.1270999, 0.1133874, 0.06605069, 
    0.05982541, 0.0738844, 0.04945484, 0.05619061, 0.05465118, 0.0784523, 
    0.03171839, 0.02292731, 0.04355092, 0.05273357, 0.02865759, 0.04177994, 
    0.05623224, 0.0467402, 0.04081125, 0.03104803, 0.08701775,
  -1.691968e-06, 3.867396e-07, 9.837087e-09, 0.02862157, 0.01540187, 
    0.08711192, 0.09003823, 0.1403804, 0.03373266, 0.2052484, 0.08494274, 
    0.05414013, 0.06968241, 0.06607901, 0.0764253, 0.05115222, 0.06243637, 
    0.1173481, 0.1408007, 0.2403997, 0.098402, 0.1102971, 0.09478611, 
    0.03027512, 0.06027078, 0.1424715, 0.3863605, -8.616472e-05, 0.0001631731,
  3.683013e-07, 2.306035e-08, 9.277823e-10, -1.136301e-07, 2.460757e-07, 
    0.001515712, -1.031527e-05, -0.0002889338, 0.0003152583, 0.1413879, 
    0.1118859, 0.1250612, 0.08983711, 0.04280075, 0.03837209, 0.05123461, 
    0.0317695, 0.05961775, 0.280041, 0.1807942, 6.169317e-05, 0.07727198, 
    0.03270013, 0.03800313, 0.06496581, 0.09325653, 0.1036845, 0.0365511, 
    3.488686e-07,
  2.581731e-07, -1.648041e-06, 0.002191739, 0.004943298, 0.048536, 
    0.002500353, -0.00147576, -0.0002674889, 0.01688897, 0.1613575, 
    0.2138866, 0.1984617, 0.2684523, 0.1802643, 0.2067456, 0.1994008, 
    0.1884845, 0.224607, 0.3420552, 0.10202, 0.01455585, 0.172626, 
    0.08298323, 0.1214717, 0.1380614, 0.1424693, 0.1884797, 0.2379673, 
    0.009762804,
  0.003029746, 0.01253964, 0.04008065, 0.1210609, 0.009249139, 0.001831413, 
    0.1163354, 0.0181318, 0.02025757, 0.0652907, 0.1403034, 0.0953472, 
    0.2288737, 0.2188583, 0.2574936, 0.2877689, 0.2265441, 0.2329305, 
    0.3520221, 0.1572765, 0.1207235, 0.2338203, 0.1307276, 0.1279828, 
    0.2577752, 0.2324595, 0.2913215, 0.2580982, 0.08769228,
  0.1507812, 0.2597288, 0.05786754, 0.01557132, 0.05566663, 0.1480236, 
    0.1767347, 0.2154734, 0.07833607, 0.04045897, 0.08873272, 0.2127195, 
    0.1742489, 0.3100623, 0.2678454, 0.3070723, 0.266959, 0.3400989, 
    0.2810066, 0.2655669, 0.1011666, 0.1237823, 0.2004966, 0.3760568, 
    0.4636158, 0.5661694, 0.3602227, 0.184158, 0.1869983,
  0.2571618, 0.3383413, 0.2080189, 0.1263632, 0.1187427, 0.177549, 0.2131254, 
    0.1328499, 0.1000427, 0.05041149, 0.1098028, 0.1386938, 0.04521829, 
    0.2288731, 0.3335712, 0.2403619, 0.3101862, 0.370934, 0.1422339, 
    0.02834755, 0.08166611, 0.1576365, 0.2862445, 0.2726803, 0.4673258, 
    0.1097169, 0.1453153, 0.1991042, 0.3123612,
  0.3147078, 0.2137218, 0.2410648, 0.2087068, 0.2422057, 0.2303937, 
    0.1841089, 0.1208068, 0.2042665, 0.2835655, 0.3000142, 0.3084469, 
    0.2495875, 0.3055263, 0.2108118, 0.1833481, 0.2276103, 0.07666151, 
    0.03806272, 0.1000145, 0.1014906, 0.08730172, 0.06127556, 0.1105403, 
    0.04807567, 0.3316435, 0.1472393, 0.06710329, 0.4326934,
  0.3421515, 0.3805921, 0.3893444, 0.2721998, 0.3227707, 0.2846528, 
    0.2898739, 0.2249862, 0.2568127, 0.2037177, 0.1545991, 0.1094012, 
    0.1002075, 0.1137102, 0.121441, 0.1227185, 0.1068129, 0.09052712, 
    0.1415995, 0.1636883, 0.1538872, 0.1974204, 0.2057548, 0.2211239, 
    0.1668013, 0.2457241, 0.2618253, 0.146131, 0.2992589,
  0.4513431, 0.4535102, 0.4556772, 0.4578443, 0.4600114, 0.4621785, 
    0.4643456, 0.4484296, 0.4581556, 0.4678817, 0.4776078, 0.4873338, 
    0.4970599, 0.5067859, 0.5028664, 0.4951833, 0.4875001, 0.4798169, 
    0.4721337, 0.4644506, 0.4567674, 0.456395, 0.4521851, 0.4479751, 
    0.4437652, 0.4395552, 0.4353452, 0.4311353, 0.4496094,
  0.1757396, 0.2471377, 0.3098411, 0.2482672, 0.2052982, 0.2396761, 
    0.2762713, 0.3206433, 0.1637988, 0.1454148, 0.2624581, 0.3047836, 
    0.3468721, 0.06846137, 0.1703007, 0.3400465, 0.3458812, 0.4491938, 
    0.4141753, 0.3990388, 0.7467006, 0.5476857, 0.3444947, 0.2333324, 
    0.3778136, 0.5211676, 0.3089167, 0.2380604, 0.230542,
  0.3018369, 0.2087882, 0.1866591, 0.1118203, 0.1842801, 0.2420938, 
    0.1295202, 0.3929314, 0.3963754, 0.3664311, 0.3069552, 0.0724904, 
    0.1570456, 0.2407344, 0.3791057, 0.4445534, 0.3634778, 0.4404221, 
    0.4558561, 0.4424838, 0.4931856, 0.4881592, 0.3997854, 0.398753, 
    0.3571614, 0.3133057, 0.3394893, 0.3951879, 0.235945,
  0.3506056, 0.3205062, 0.2509395, 0.2970464, 0.2876658, 0.3138434, 
    0.3250975, 0.3313002, 0.3561404, 0.3923873, 0.388033, 0.4673059, 0.54713, 
    0.4094822, 0.332934, 0.3660372, 0.4279296, 0.4706883, 0.4693135, 
    0.4013826, 0.3863834, 0.4400693, 0.4213924, 0.3011826, 0.343368, 
    0.4886238, 0.4856805, 0.3469788, 0.2985819,
  0.3151824, 0.3056203, 0.3502105, 0.2696347, 0.2735101, 0.279954, 0.3505503, 
    0.3140029, 0.2856938, 0.2822529, 0.2953869, 0.3756417, 0.3054118, 
    0.1682854, 0.1583399, 0.2335536, 0.3031516, 0.1849562, 0.2621786, 
    0.2800824, 0.3253801, 0.3205299, 0.2611389, 0.2174673, 0.1474053, 
    0.1911993, 0.2341611, 0.3110348, 0.3256876,
  0.3461821, 0.2622924, 0.2046841, 0.1640326, 0.1965046, 0.1962878, 
    0.1618068, 0.2239791, 0.2607367, 0.2337141, 0.1227692, 0.1123161, 
    0.01917531, 0.1060209, 0.3440737, 0.08700718, 0.2300639, 0.147541, 
    0.1644312, 0.2273011, 0.3144296, 0.3045715, 0.1720702, 0.3980907, 
    0.03006997, 0.05549579, 0.1418732, 0.2320532, 0.3016883,
  0.1526192, 0.07284243, 0.00534006, 0.0522886, 0.09022447, 0.09083481, 
    0.05393088, 0.08861827, 0.08821169, 0.03488541, 0.008424459, 
    -3.145977e-05, 0.01667492, 0.04775694, 0.07238095, 0.07988441, 
    0.06352723, 0.04282399, 0.1226751, 0.1061155, 0.1258567, 0.04812769, 
    0.05746347, 0.01983684, 0.07439534, 0.05819569, 0.09919602, 0.08835483, 
    0.1614851,
  0.16174, 1.250698e-05, 1.733184e-05, 0.05419364, 0.01261919, 0.08248058, 
    0.03828939, 0.02942724, 0.09036318, 0.00363442, 1.567903e-05, 
    0.0002343376, 0.01799874, 0.09000819, 0.04770124, 0.0248454, 0.04874406, 
    0.06936529, 0.01901285, 0.0139076, 0.01569633, 0.02863965, 0.1289317, 
    0.04477972, 0.05839322, 0.04629089, 0.02755856, 0.0129928, 0.04761029,
  0.3788763, 0.0578333, 0.04010343, 0.1235941, 0.03059676, 0.02787375, 
    0.05117349, 0.04526525, 0.05200256, 0.01985672, 0.04506784, 0.02297989, 
    0.08906326, 0.05217015, 0.01958407, 0.02727957, 0.03047823, 0.01574053, 
    0.0127775, 0.02290264, 0.02851376, 0.05835694, 0.37892, 0.01181285, 
    0.04351744, 0.0008643041, 0.05348881, 0.02756354, 0.09578507,
  0.1786701, 0.01007132, 0.002017407, 0.01172146, 0.07855515, 0.03866072, 
    0.05139001, 0.02481933, 0.03118097, 0.09071783, 0.05782482, 0.1382605, 
    0.03323336, 0.04191879, 0.03255943, 0.1212613, 0.1615133, 0.1733017, 
    0.1365564, 0.164227, 0.09256712, 0.1641419, 0.04534131, 0.02701401, 
    0.02868064, 0.04737563, 0.06850444, 0.1058135, 0.2338688,
  -3.621836e-07, 3.758818e-07, 1.936849e-08, 0.0197738, 0.01487672, 
    0.02095623, 0.03504509, 0.0242673, 0.01079051, 0.06352194, 0.05937758, 
    0.04299356, 0.03351308, 0.0301041, 0.03902315, 0.02723541, 0.02178794, 
    0.04730937, 0.08920117, 0.1127526, 0.06973879, 0.01813595, 0.2377285, 
    0.05604006, 0.00971368, 0.04284588, 0.1988025, 0.01917376, 5.860981e-05,
  3.239086e-07, 2.039962e-08, 8.143614e-10, -9.145369e-08, -3.258338e-05, 
    0.001019199, -8.119004e-05, 0.01936838, 0.0001681243, 0.233691, 
    0.1186878, 0.1136557, 0.07369444, 0.02534206, 0.0106673, 0.01402359, 
    0.01189483, 0.01768834, 0.1777059, 0.1886789, 0.0004392787, 0.06858298, 
    0.01423123, 0.01271414, 0.02679927, 0.038564, 0.05944652, 0.01009378, 
    2.765019e-07,
  1.692855e-07, -5.918014e-05, 0.0004733287, 0.002937906, 0.03402754, 
    0.002621075, -0.001357083, -0.000199342, 0.01789513, 0.1272655, 
    0.2099105, 0.1478258, 0.2683325, 0.1901198, 0.1679081, 0.2463129, 
    0.2347683, 0.2668476, 0.224871, 0.1168492, 0.01299665, 0.173486, 
    0.06979404, 0.1159054, 0.07699934, 0.0792745, 0.1028561, 0.1431248, 
    0.009516571,
  0.00125749, 0.005955991, 0.02844789, 0.1175003, 0.001774095, 0.0009961766, 
    0.1141642, 0.01424524, 0.01714767, 0.06152131, 0.1347974, 0.08398651, 
    0.2059382, 0.1960379, 0.261643, 0.2485045, 0.2308897, 0.2028177, 
    0.2685977, 0.1508834, 0.1156222, 0.2373412, 0.1059258, 0.1207069, 
    0.2596873, 0.2185072, 0.2710923, 0.2435496, 0.0773216,
  0.1185755, 0.2325896, 0.04233781, 0.01530961, 0.03868319, 0.1194744, 
    0.1368629, 0.1948589, 0.05836561, 0.03521728, 0.090524, 0.2220361, 
    0.2103216, 0.3296297, 0.2082031, 0.2583545, 0.2299614, 0.3404842, 
    0.2552048, 0.2473166, 0.08946073, 0.1237797, 0.1629048, 0.3672454, 
    0.4472119, 0.5754228, 0.3251697, 0.1845007, 0.1751702,
  0.2047674, 0.3341645, 0.1725748, 0.1084463, 0.1444337, 0.2257361, 
    0.1730419, 0.1142242, 0.0713084, 0.03332388, 0.05722879, 0.09032914, 
    0.04336324, 0.1955763, 0.2225755, 0.1966469, 0.3037629, 0.346853, 
    0.1376974, 0.02961642, 0.07361957, 0.1545902, 0.2578607, 0.2546091, 
    0.3935609, 0.1076812, 0.1080276, 0.1247513, 0.2492354,
  0.2746948, 0.17082, 0.2678649, 0.168765, 0.2283274, 0.2337674, 0.1998225, 
    0.1025289, 0.1936011, 0.2226675, 0.2830317, 0.2932885, 0.2276168, 
    0.3129497, 0.2501963, 0.2086583, 0.2196899, 0.1334873, 0.05074899, 
    0.1697847, 0.1726821, 0.07773823, 0.09287783, 0.1341149, 0.05986121, 
    0.3241624, 0.170202, 0.0340368, 0.368965,
  0.4028035, 0.4005051, 0.4106854, 0.2395813, 0.3238655, 0.3261511, 
    0.3655421, 0.2845001, 0.3085239, 0.2304823, 0.1566057, 0.1264235, 
    0.08678819, 0.1387949, 0.1458236, 0.1510971, 0.1449444, 0.1256195, 
    0.1696125, 0.1840417, 0.1640464, 0.2277084, 0.2069829, 0.2327674, 
    0.16909, 0.2434203, 0.238912, 0.1376305, 0.3143006,
  0.4753781, 0.4742626, 0.4731471, 0.4720316, 0.470916, 0.4698005, 0.468685, 
    0.4332013, 0.4420595, 0.4509176, 0.4597758, 0.4686339, 0.4774921, 
    0.4863502, 0.4935679, 0.4884287, 0.4832896, 0.4781504, 0.4730112, 
    0.467872, 0.4627328, 0.4653755, 0.462772, 0.4601686, 0.4575652, 
    0.4549617, 0.4523583, 0.4497549, 0.4762705,
  0.2376152, 0.3482167, 0.3100131, 0.2827251, 0.2229742, 0.2167436, 
    0.2724674, 0.3686457, 0.191595, 0.1933455, 0.2481779, 0.3122748, 
    0.4513888, 0.04046221, 0.1972432, 0.3078263, 0.3187897, 0.4032573, 
    0.3787849, 0.3923173, 0.7624537, 0.6293417, 0.3346522, 0.2265582, 
    0.3573452, 0.5360622, 0.3285258, 0.2080436, 0.2932541,
  0.2360123, 0.1503293, 0.1631404, 0.06814732, 0.1459128, 0.2570561, 
    0.06409393, 0.3562924, 0.4022209, 0.3750392, 0.2722874, 0.07572469, 
    0.1519637, 0.1698374, 0.3149153, 0.4050891, 0.3437859, 0.383811, 
    0.4228559, 0.479065, 0.4856546, 0.5307841, 0.4145141, 0.4387789, 
    0.335375, 0.3066221, 0.3284771, 0.3008258, 0.2783524,
  0.29489, 0.2779837, 0.202778, 0.2429416, 0.2702098, 0.3147719, 0.2758721, 
    0.2908755, 0.308183, 0.3362549, 0.3799081, 0.4476745, 0.5064347, 
    0.3629611, 0.3063928, 0.3456859, 0.4192047, 0.4259406, 0.4505523, 
    0.4202409, 0.4368261, 0.4072542, 0.363872, 0.2744736, 0.3049768, 
    0.4455017, 0.3960589, 0.3056866, 0.2568837,
  0.274645, 0.2898296, 0.3470826, 0.2494226, 0.2696425, 0.2907335, 0.3446701, 
    0.3073989, 0.3147507, 0.2983922, 0.2707331, 0.3367076, 0.2596049, 
    0.1546927, 0.1091106, 0.1871218, 0.2572071, 0.1859914, 0.2442953, 
    0.2259047, 0.2593499, 0.3174704, 0.2441582, 0.2037377, 0.1301675, 
    0.1461753, 0.2073773, 0.3007285, 0.3094581,
  0.3348802, 0.2111469, 0.145082, 0.1447081, 0.1894824, 0.2094286, 0.1099362, 
    0.1622587, 0.1973605, 0.20556, 0.07897872, 0.05475079, 0.01416233, 
    0.05874895, 0.3399938, 0.08136486, 0.1872653, 0.1147838, 0.1280707, 
    0.189261, 0.3129038, 0.2291994, 0.1199013, 0.4119241, 0.01881067, 
    0.05508911, 0.1432317, 0.1831455, 0.2583121,
  0.05747651, 0.08692454, 0.005003827, 0.02984551, 0.05190081, 0.06507991, 
    0.01688066, 0.02673584, 0.05120898, 0.02529283, 0.003760367, 
    -5.457639e-06, 0.01686628, 0.03283982, 0.05229481, 0.04055221, 
    0.05174965, 0.03982348, 0.1535518, 0.09364694, 0.06697037, 0.01531401, 
    0.02966248, 0.02402749, 0.04975374, 0.03991318, 0.07322422, 0.03796132, 
    0.07909498,
  0.05717186, -0.0007218391, -1.196998e-06, 0.007882609, -0.001597289, 
    0.03739036, 0.01926631, 0.009649804, 0.04343021, 0.0006494189, 
    4.976274e-06, 6.484166e-05, 0.01694137, 0.04933006, 0.0172059, 
    0.01217211, 0.01747728, 0.03097599, 0.003940941, 0.004657558, 
    0.001475576, 0.003814264, 0.03029069, 0.1457607, 0.04242798, 0.03696854, 
    0.001543356, 0.00131189, 0.01280998,
  0.1322223, 0.07176859, 0.0282358, 0.1185246, 0.01191502, 0.01121747, 
    0.01487041, 0.01143364, 0.01995148, 0.0009568133, 0.02509292, 
    0.008840183, 0.06930096, 0.007739589, 0.007528866, 0.004230645, 
    0.008611945, 0.005621758, 0.00216684, 0.005288336, 0.006034035, 
    0.0100412, 0.1191667, 0.008421893, 0.03832096, 0.0002930845, 0.02666043, 
    0.006021193, 0.02550998,
  0.02452321, 0.007799224, 0.001215022, 0.003645128, 0.01195017, 0.007073314, 
    0.006525983, 0.002340355, 0.03743497, 0.06560835, 0.02756291, 0.02004987, 
    0.02240534, 0.03267302, 0.004982379, 0.01280472, 0.02895087, 0.05080312, 
    0.1462199, 0.3392215, 0.1389803, 0.1256196, 0.1789936, 0.02603816, 
    0.01852767, 0.02505167, 0.01738623, 0.0113444, 0.03533889,
  -1.61839e-08, 3.660015e-07, 1.981274e-08, 0.01905369, 0.01535914, 
    0.004763674, 0.01168751, 0.004370623, 0.001109968, 0.01056917, 
    0.01699537, 0.009676595, 0.0229312, 0.007861677, 0.01717775, 0.01303689, 
    0.003954511, 0.0106304, 0.03089497, 0.04385265, 0.03369235, 0.003684717, 
    0.2859643, 0.06912979, 0.0005174682, 0.01096224, 0.07550643, 0.1147912, 
    0.0001053185,
  3.034053e-07, 1.873332e-08, 7.835134e-10, -1.073216e-07, -2.348623e-05, 
    5.288759e-05, -3.94327e-05, 0.003370561, 8.691251e-05, 0.249342, 
    0.06861871, 0.04484077, 0.02073309, 0.001862987, 0.001342335, 
    0.002131123, 0.006869083, 0.01226849, 0.06563312, 0.0785905, 0.008106242, 
    0.05711886, 0.004387098, 0.001654111, 0.00960347, 0.007846732, 
    0.08566547, 0.004027158, 2.42238e-07,
  1.201903e-07, -6.034762e-05, 5.854768e-05, 0.001906226, 0.02304695, 
    0.003478233, -0.001206901, -8.755154e-05, 0.01941076, 0.1097957, 
    0.1974038, 0.1318434, 0.2745204, 0.1975588, 0.1127462, 0.1780044, 
    0.196711, 0.1502606, 0.0847918, 0.06114894, 0.009569012, 0.1825373, 
    0.06398711, 0.07448858, 0.05860316, 0.06999442, 0.04835937, 0.05385813, 
    0.01308487,
  -0.0006300742, 0.002323277, 0.02310475, 0.1178779, -1.742484e-05, 
    0.0002210793, 0.1063457, 0.007605566, 0.01395243, 0.0630959, 0.128092, 
    0.07664872, 0.1493217, 0.174545, 0.2459419, 0.2372995, 0.2314359, 
    0.186608, 0.171246, 0.15036, 0.09834515, 0.2366391, 0.0964727, 0.104537, 
    0.2313924, 0.1694868, 0.1793578, 0.1868508, 0.05756415,
  0.09853456, 0.2027205, 0.02886688, 0.01183535, 0.08787178, 0.07152685, 
    0.108864, 0.1560036, 0.04601353, 0.02726416, 0.08464805, 0.2053749, 
    0.1774146, 0.2858551, 0.1449843, 0.2173498, 0.2159953, 0.3330611, 
    0.217108, 0.2269857, 0.0805434, 0.1288907, 0.1283894, 0.3525434, 
    0.4064573, 0.4819821, 0.3021787, 0.1897972, 0.1814159,
  0.1923945, 0.3335409, 0.1515943, 0.1026726, 0.1680162, 0.183612, 0.1591367, 
    0.08042493, 0.04786561, 0.0221161, 0.03568408, 0.06074521, 0.02656859, 
    0.1452221, 0.1612445, 0.1858623, 0.2706396, 0.3267797, 0.1115912, 
    0.028721, 0.06730586, 0.1238996, 0.2513849, 0.2453003, 0.2947351, 
    0.1242797, 0.08303364, 0.08483303, 0.2072121,
  0.2382256, 0.1482677, 0.279182, 0.1734012, 0.2624474, 0.2512296, 0.1798985, 
    0.09214083, 0.1429405, 0.1765832, 0.2620573, 0.2965713, 0.2028048, 
    0.3307008, 0.3235223, 0.2947085, 0.2388863, 0.1498029, 0.07324998, 
    0.2609774, 0.1569152, 0.07347707, 0.07216091, 0.1391699, 0.09195253, 
    0.3288015, 0.1888136, 0.01079874, 0.2807994,
  0.46107, 0.4524928, 0.4511905, 0.2619102, 0.3324275, 0.3534785, 0.4039408, 
    0.3074325, 0.2997132, 0.2331628, 0.1928762, 0.1485504, 0.1035138, 
    0.1575762, 0.1800847, 0.1787556, 0.156906, 0.1596819, 0.2011971, 
    0.2167655, 0.1760727, 0.2366399, 0.2215841, 0.2201772, 0.139694, 
    0.2623002, 0.2473823, 0.1159222, 0.2883422,
  0.3653514, 0.3618405, 0.3583296, 0.3548187, 0.3513078, 0.3477969, 0.344286, 
    0.3395079, 0.3497638, 0.3600196, 0.3702754, 0.3805313, 0.3907871, 
    0.4010429, 0.3787993, 0.3775104, 0.3762215, 0.3749326, 0.3736437, 
    0.3723548, 0.3710659, 0.4142657, 0.4088096, 0.4033536, 0.3978976, 
    0.3924415, 0.3869855, 0.3815295, 0.3681601,
  0.2853765, 0.3674977, 0.2741406, 0.2581165, 0.2162563, 0.1928195, 
    0.2339728, 0.3151321, 0.19577, 0.1489532, 0.2408452, 0.2995441, 
    0.5139453, 0.0156113, 0.24659, 0.3185735, 0.33102, 0.3664897, 0.3465275, 
    0.3962751, 0.7739366, 0.6924903, 0.3154736, 0.2255386, 0.4147133, 
    0.5597916, 0.3041481, 0.1865824, 0.2792722,
  0.1784233, 0.1017623, 0.1665669, 0.04371315, 0.114923, 0.2476717, 
    0.01984356, 0.3292302, 0.3810158, 0.351026, 0.2417075, 0.09074923, 
    0.1346885, 0.1297702, 0.2539954, 0.3553434, 0.2922653, 0.324201, 
    0.3781146, 0.4447527, 0.4846991, 0.5314112, 0.416781, 0.4468871, 0.31561, 
    0.3240418, 0.3267758, 0.2129376, 0.316754,
  0.2462896, 0.2300523, 0.1638357, 0.2081805, 0.2376376, 0.2738768, 
    0.2213407, 0.244922, 0.2636176, 0.2688517, 0.342473, 0.4078738, 
    0.4386221, 0.317389, 0.2733794, 0.3224464, 0.3955626, 0.4326223, 
    0.4165945, 0.3833964, 0.3975828, 0.3926398, 0.3147173, 0.2510439, 
    0.2692073, 0.3993201, 0.3291667, 0.2519192, 0.2213065,
  0.2400617, 0.2529052, 0.2945268, 0.21706, 0.2454855, 0.2814819, 0.3234096, 
    0.2758275, 0.2725754, 0.2773463, 0.2347732, 0.2764001, 0.2096672, 
    0.1251529, 0.08422873, 0.1446562, 0.2012447, 0.1644485, 0.2150083, 
    0.1889528, 0.2272039, 0.282953, 0.1945074, 0.17384, 0.1060042, 0.1006016, 
    0.1787696, 0.2548906, 0.2991104,
  0.2637822, 0.1372495, 0.1009748, 0.1210822, 0.1687122, 0.1653102, 
    0.07365193, 0.1095629, 0.1472549, 0.1899289, 0.06458452, 0.02421219, 
    0.01074077, 0.04120598, 0.3028433, 0.07098827, 0.1512509, 0.09146006, 
    0.09453742, 0.1679731, 0.264423, 0.1611036, 0.08196545, 0.4045059, 
    0.01285969, 0.05484569, 0.1234387, 0.1321639, 0.2145549,
  0.02299799, 0.04885327, 0.006274341, 0.01178978, 0.01717398, 0.02984487, 
    0.009201836, 0.01236562, 0.03404583, 0.01981783, 0.001327217, 
    -6.720424e-07, 0.01905353, 0.01865702, 0.03690026, 0.02563169, 
    0.03827104, 0.03145593, 0.1305519, 0.05417624, 0.03743959, 0.004567141, 
    0.01288657, 0.01759082, 0.04142079, 0.02449081, 0.05420639, 0.01381253, 
    0.03600371,
  0.02416406, -4.004044e-05, -6.379951e-06, 0.002155761, -0.00353056, 
    0.01504189, 0.007723243, 0.001498022, 0.01566561, 5.483804e-05, 
    1.175576e-06, 2.011312e-05, 0.005526552, 0.0157066, 0.007020927, 
    0.002982221, 0.003759692, 0.01629795, 0.0002738945, 0.001227468, 
    0.000462098, 0.0009827266, 0.01154534, 0.08227782, 0.02401781, 
    0.03152895, 0.000177636, 0.0001495815, 0.004388282,
  0.05084064, 0.05150726, 0.03152477, 0.102522, 0.008021891, 0.002277836, 
    0.006093273, 0.002750402, 0.0070983, -0.0006698747, 0.01155602, 
    0.003115381, 0.05276037, 0.001837064, 0.0005909698, 0.0004692133, 
    0.001773534, 0.002333878, 0.0005152453, 0.001099144, 0.001253085, 
    0.00308672, 0.04287156, 0.01427979, 0.03709821, 9.965307e-05, 
    0.009716514, 0.002382598, 0.009453187,
  0.006589527, 0.01105426, 0.001177141, 0.001289729, 0.004250563, 
    0.002513502, 0.00225464, 0.0002961842, 0.04608154, 0.0519131, 0.01044162, 
    0.004252127, 0.006345551, 0.02419794, 0.001201773, 0.0034566, 
    0.007027911, 0.01054264, 0.0294745, 0.06309128, 0.02908237, 0.03212448, 
    0.1911422, 0.02085418, 0.01820319, 0.01782935, 0.002349741, 0.002998522, 
    0.01068904,
  8.893421e-08, 3.613886e-07, 1.972891e-08, 0.01501896, 0.01250143, 
    0.001935648, 0.001328453, 0.001813437, 0.0003153498, 0.003666512, 
    0.005615883, 0.002314118, 0.005666893, 0.001582013, 0.006771727, 
    0.01290188, 0.000817023, 0.002821486, 0.009531176, 0.01298, 0.01580739, 
    0.001374978, 0.1968626, 0.0612512, 0.0002150235, 0.004348485, 0.03039064, 
    0.03538192, 0.0001420899,
  2.967161e-07, 1.745435e-08, 7.734294e-10, 2.343237e-06, -1.003729e-05, 
    1.33432e-05, -3.338693e-05, 0.001456322, 3.663469e-05, 0.1370012, 
    0.01287812, 0.0153137, 0.005573125, 0.0002371082, 0.0002645839, 
    0.0006484708, 0.003630466, 0.007741098, 0.02500734, 0.0444883, 
    0.02457661, 0.04796299, 0.001004192, -0.0005871912, 0.002006412, 
    0.002696468, 0.05101822, 0.002250769, 2.293896e-07,
  1.090142e-07, 0.0001483885, 3.285973e-05, 0.001807389, 0.01520158, 
    0.002353164, -0.001158574, -6.994761e-05, 0.01550986, 0.09291118, 
    0.176311, 0.1326097, 0.2588018, 0.1517436, 0.08517325, 0.112373, 
    0.08917931, 0.06874638, 0.03294466, 0.02910182, 0.006262474, 0.179751, 
    0.05426432, 0.05886867, 0.05111911, 0.05684187, 0.01431557, 0.02294882, 
    0.01622226,
  -0.001195645, 0.0004904112, 0.01702531, 0.1174855, -0.0003829373, 
    6.831384e-05, 0.09059565, 0.005260339, 0.01152088, 0.06173415, 0.1258606, 
    0.07001197, 0.1174748, 0.1507266, 0.2279735, 0.2165306, 0.2138373, 
    0.1623903, 0.1452308, 0.1436152, 0.08584072, 0.2210809, 0.07873033, 
    0.09471354, 0.1794123, 0.1089786, 0.1210454, 0.1120296, 0.0414395,
  0.06791823, 0.1763872, 0.01728494, 0.008140627, 0.115524, 0.04443297, 
    0.08633525, 0.1263149, 0.03271198, 0.02044837, 0.07498821, 0.1875812, 
    0.148793, 0.2127566, 0.1059918, 0.1871305, 0.2038705, 0.2738632, 
    0.1715378, 0.2108965, 0.06531725, 0.1212577, 0.1001511, 0.3295078, 
    0.3504019, 0.4204882, 0.2814233, 0.1668555, 0.1649626,
  0.1508547, 0.3304296, 0.1329062, 0.09252501, 0.1669602, 0.1411673, 
    0.1350272, 0.05912202, 0.03799847, 0.01973384, 0.02553763, 0.0352163, 
    0.02287473, 0.1092047, 0.1355218, 0.2434488, 0.2471663, 0.2990405, 
    0.0663868, 0.02304663, 0.05594408, 0.09383909, 0.2386013, 0.2352029, 
    0.2568276, 0.106539, 0.06957085, 0.05964312, 0.1784276,
  0.1937125, 0.1329406, 0.277166, 0.1572724, 0.2479801, 0.2307609, 0.1318637, 
    0.07082571, 0.09896798, 0.1313477, 0.2342744, 0.2505862, 0.2007633, 
    0.3536866, 0.3708028, 0.4134361, 0.3025596, 0.1620956, 0.1505651, 
    0.3019714, 0.1208376, 0.08981454, 0.05118578, 0.1465637, 0.09635893, 
    0.3204425, 0.1974975, 0.002883022, 0.2090279,
  0.5213481, 0.423657, 0.4662616, 0.3260955, 0.3276922, 0.398087, 0.4497994, 
    0.3639887, 0.2734945, 0.2641392, 0.2222385, 0.2125053, 0.139403, 
    0.2009487, 0.2439911, 0.2752218, 0.202145, 0.1822088, 0.2298763, 0.2035, 
    0.2111183, 0.2256842, 0.2464908, 0.2305969, 0.1407242, 0.2463407, 
    0.2263988, 0.09671954, 0.2532643,
  0.2737293, 0.2692288, 0.2647282, 0.2602277, 0.2557271, 0.2512265, 0.246726, 
    0.2232644, 0.2343889, 0.2455133, 0.2566377, 0.2677621, 0.2788866, 
    0.290011, 0.3574201, 0.3588482, 0.3602763, 0.3617044, 0.3631325, 
    0.3645607, 0.3659888, 0.350253, 0.342201, 0.3341491, 0.3260971, 
    0.3180451, 0.3099931, 0.3019412, 0.2773298,
  0.312907, 0.3103174, 0.2125011, 0.186071, 0.2042402, 0.1717955, 0.1796052, 
    0.236274, 0.1494504, 0.1114648, 0.1152983, 0.2708628, 0.4656593, 
    0.009620432, 0.2950271, 0.3781086, 0.3784428, 0.3555036, 0.2949239, 
    0.3859185, 0.7759153, 0.7553384, 0.2845507, 0.2042081, 0.4304411, 
    0.5720146, 0.283426, 0.1565182, 0.2533362,
  0.1310255, 0.0691711, 0.1288457, 0.02242299, 0.08605018, 0.2239964, 
    0.01218145, 0.2745755, 0.3516477, 0.3008549, 0.2143963, 0.09553671, 
    0.09185771, 0.1002751, 0.2017103, 0.2925558, 0.2053356, 0.2522685, 
    0.3193706, 0.3894399, 0.4425113, 0.4845831, 0.3830329, 0.4576947, 
    0.3065204, 0.3409463, 0.3112645, 0.1607481, 0.324714,
  0.1923213, 0.1920913, 0.1285782, 0.1696409, 0.1924795, 0.2197495, 
    0.1993189, 0.1942755, 0.207437, 0.2193044, 0.2870338, 0.3475522, 
    0.3646598, 0.2593379, 0.2145056, 0.2575103, 0.3332792, 0.400277, 
    0.3617491, 0.3119899, 0.3557039, 0.3448085, 0.2842366, 0.1986793, 
    0.2440357, 0.3520767, 0.2864753, 0.204423, 0.1713651,
  0.2015919, 0.1947131, 0.2362854, 0.1629427, 0.2066676, 0.2358283, 
    0.2840171, 0.2175755, 0.2083872, 0.2275387, 0.1793585, 0.2137482, 
    0.1504537, 0.09933311, 0.05612187, 0.09286313, 0.1445557, 0.1169926, 
    0.1637208, 0.159022, 0.187945, 0.2195285, 0.1541701, 0.1453151, 
    0.08110581, 0.07503169, 0.1547691, 0.2162413, 0.2500157,
  0.1915429, 0.0774433, 0.068646, 0.08912271, 0.1281081, 0.1003354, 
    0.04467694, 0.07165273, 0.1002483, 0.1593076, 0.04938729, 0.01326618, 
    0.008354337, 0.02677056, 0.2623641, 0.05247926, 0.1173685, 0.07037378, 
    0.06771138, 0.1341216, 0.2179396, 0.1432521, 0.05596239, 0.3841088, 
    0.008042505, 0.04565988, 0.09267382, 0.08752928, 0.1712165,
  0.01016384, 0.02271698, 0.007871434, 0.004263564, 0.006422277, 0.01418326, 
    0.005660907, 0.007562366, 0.02048852, 0.01298107, 0.0007887911, 
    -5.296662e-07, 0.02155657, 0.01177047, 0.03553102, 0.01248013, 
    0.02208795, 0.01517298, 0.07344787, 0.02590866, 0.02447689, 0.00212735, 
    0.006822772, 0.01000178, 0.043236, 0.01556176, 0.0296527, 0.004633588, 
    0.01535755,
  0.01297314, -0.0001768862, -5.55039e-06, 0.001055716, -0.00274957, 
    0.006210314, 0.002192971, 0.0005276558, 0.004681225, 3.057202e-05, 
    4.615493e-07, 7.906514e-06, 0.00249393, 0.008976231, 0.004227002, 
    0.0003313808, 0.001222072, 0.007320154, 5.406463e-05, 0.0009178487, 
    0.0002307582, 0.0005369401, 0.006362132, 0.0378612, 0.01230211, 
    0.02906136, 6.731186e-05, 6.841825e-05, 0.002123208,
  0.02521694, 0.03507886, 0.04502499, 0.087868, 0.006172198, 0.0008053487, 
    0.00287672, 0.000950581, 0.002290105, -0.0002132475, 0.005819295, 
    0.001017994, 0.02995977, 0.0007420359, 0.0001176784, 0.0001895368, 
    0.0008230355, 0.0008853402, 0.0002643893, 0.0004590135, 0.0005824302, 
    0.001440498, 0.02190476, 0.01184448, 0.03985131, 6.497368e-05, 
    0.001973679, 0.001258217, 0.004951587,
  0.003195004, 0.01421599, 0.0006524131, 3.916967e-05, 0.002209034, 
    0.001398623, 0.001150809, 0.0001284752, 0.04380185, 0.04618508, 
    0.006858708, 0.001801917, 0.003153266, 0.01221361, 0.0005189788, 
    0.001631697, 0.003292463, 0.004695544, 0.01274525, 0.02487161, 
    0.007947584, 0.00771487, 0.07740615, 0.02207154, 0.01792447, 0.008124833, 
    0.0004802849, 0.001588312, 0.004863909,
  1.250666e-07, 3.598896e-07, 1.994724e-08, 0.01761248, 0.006997792, 
    0.001151207, -0.0005344168, 0.001075319, 0.0001693483, 0.002030116, 
    0.00101704, 0.0007753822, 0.0008382507, 0.0003756647, 0.00232085, 
    0.006373155, 0.0004706997, 0.001234842, 0.003214013, 0.004559204, 
    0.006785617, 0.0008250015, 0.1164003, 0.0491791, 0.0001173795, 
    0.002317626, 0.01515017, 0.01819436, 8.749803e-05,
  2.926432e-07, 1.647599e-08, 7.720876e-10, 2.322405e-05, -5.131531e-06, 
    6.036258e-06, -2.583074e-05, 0.0005595992, 1.826006e-05, 0.05779866, 
    0.004526511, 0.005672207, 0.00177871, 0.0001358333, 0.000144103, 
    0.0003664164, 0.001297727, 0.00279382, 0.01363358, 0.02835119, 
    0.02078087, 0.03421922, 0.0003856963, -0.0007584747, 0.0007982777, 
    0.00148022, 0.0287616, 0.001477047, 2.234551e-07,
  1.162293e-07, 0.0001250087, 9.17401e-06, 0.001068594, 0.00590863, 
    0.00172317, -0.001124206, -9.232664e-05, 0.01131025, 0.07063123, 
    0.139376, 0.1023886, 0.1893804, 0.1014695, 0.06450149, 0.07005399, 
    0.04636275, 0.03516893, 0.01831964, 0.02013925, 0.005112566, 0.1513412, 
    0.04547276, 0.0391329, 0.04103364, 0.035023, 0.005556738, 0.01278621, 
    0.01319073,
  -0.001098017, 0.0001137843, 0.00779586, 0.1055948, -0.000540046, 
    8.177648e-05, 0.07174923, 0.003572566, 0.008784354, 0.05912809, 
    0.1209652, 0.06941202, 0.09462068, 0.1295315, 0.1891601, 0.1762451, 
    0.1715506, 0.1266374, 0.1067513, 0.1331814, 0.07511158, 0.2049272, 
    0.0643349, 0.0905443, 0.1313761, 0.06563774, 0.06137148, 0.07157256, 
    0.02429881,
  0.04618753, 0.1481231, 0.01075764, 0.003506156, 0.1105619, 0.02845712, 
    0.07049579, 0.1020387, 0.02861421, 0.01473722, 0.06366803, 0.1652411, 
    0.1252883, 0.1457155, 0.07552879, 0.1624167, 0.1788957, 0.2145094, 
    0.125977, 0.1920216, 0.05249427, 0.09910633, 0.08072152, 0.3056799, 
    0.2993644, 0.4199956, 0.2432458, 0.1371727, 0.1220382,
  0.118096, 0.3091359, 0.117698, 0.08280008, 0.1545279, 0.1207088, 0.114043, 
    0.04584003, 0.03107319, 0.01695255, 0.01919768, 0.0240634, 0.02960469, 
    0.07176843, 0.1241299, 0.2386107, 0.2161207, 0.2582461, 0.04400064, 
    0.02234182, 0.0446768, 0.09448504, 0.2316413, 0.2189427, 0.2182488, 
    0.08395335, 0.05316358, 0.0449379, 0.1587183,
  0.1517109, 0.1023983, 0.2725467, 0.142379, 0.221951, 0.2057006, 0.09970304, 
    0.04966649, 0.07032634, 0.1071616, 0.2027659, 0.2119543, 0.172702, 
    0.3628951, 0.3251094, 0.442736, 0.2743809, 0.17455, 0.2068677, 0.309084, 
    0.1436602, 0.08820893, 0.03998941, 0.1452551, 0.1349773, 0.2948141, 
    0.2143747, -0.003287558, 0.1695862,
  0.5584288, 0.4271948, 0.4484685, 0.3506535, 0.3550723, 0.3934475, 
    0.4741659, 0.3936104, 0.2625802, 0.2622707, 0.2481448, 0.2303857, 
    0.1991179, 0.2495652, 0.2688216, 0.2896954, 0.2509086, 0.2436893, 
    0.2406825, 0.2275096, 0.2568051, 0.2124293, 0.2356063, 0.245655, 
    0.1400342, 0.2344929, 0.1923746, 0.09011603, 0.2321722,
  0.1920229, 0.1834596, 0.1748964, 0.1663331, 0.1577699, 0.1492066, 
    0.1406434, 0.1250083, 0.1321926, 0.139377, 0.1465613, 0.1537457, 0.16093, 
    0.1681143, 0.1932503, 0.2026094, 0.2119686, 0.2213278, 0.230687, 
    0.2400462, 0.2494054, 0.2765943, 0.268614, 0.2606337, 0.2526534, 
    0.2446731, 0.2366928, 0.2287125, 0.1988735,
  0.3483743, 0.2742096, 0.12767, 0.1967881, 0.1854157, 0.1244721, 0.145523, 
    0.1231048, 0.07985131, 0.1420134, 0.1294491, 0.2015968, 0.3481621, 
    0.004385056, 0.3405535, 0.5160519, 0.4356247, 0.3515514, 0.2483564, 
    0.3468225, 0.7899054, 0.8308687, 0.2569044, 0.1720911, 0.3743463, 
    0.5825449, 0.2430612, 0.131143, 0.2522301,
  0.1143888, 0.05176713, 0.1000103, 0.01132913, 0.06559508, 0.198483, 
    0.01337106, 0.198722, 0.2821295, 0.2325617, 0.1814652, 0.09208805, 
    0.05436747, 0.08615589, 0.1545053, 0.2296464, 0.14299, 0.1849877, 
    0.2427401, 0.3046646, 0.3683493, 0.4210585, 0.3439578, 0.4490648, 
    0.2663405, 0.3536954, 0.2713441, 0.1257714, 0.3382484,
  0.1392653, 0.1475434, 0.09648568, 0.1293372, 0.1427562, 0.1688924, 
    0.1514879, 0.1473792, 0.1657253, 0.1658789, 0.2282555, 0.2755797, 
    0.2957823, 0.2002113, 0.1462715, 0.1838815, 0.2407468, 0.3283724, 
    0.2940431, 0.2427905, 0.2914091, 0.2604476, 0.2250117, 0.1383121, 
    0.206206, 0.2923894, 0.2467722, 0.1659075, 0.1273262,
  0.1500024, 0.1503869, 0.1770955, 0.117388, 0.1668686, 0.191659, 0.2386003, 
    0.1583414, 0.1379541, 0.1677916, 0.1271066, 0.1500138, 0.09223796, 
    0.06605028, 0.03902799, 0.05580609, 0.09752999, 0.0850391, 0.1132563, 
    0.1095245, 0.1508486, 0.1505569, 0.121733, 0.1189992, 0.05486254, 
    0.05541551, 0.1235092, 0.179013, 0.1983939,
  0.1295383, 0.04388174, 0.0472649, 0.05747084, 0.08043501, 0.06443851, 
    0.02594549, 0.03944548, 0.05756063, 0.1138733, 0.03098559, 0.007604546, 
    0.005810279, 0.01549027, 0.2282352, 0.0333624, 0.07738815, 0.04574217, 
    0.04181117, 0.09363738, 0.1571235, 0.1157299, 0.03485454, 0.3470947, 
    0.00437141, 0.03237832, 0.06388354, 0.04802259, 0.1137148,
  0.006249215, 0.01333954, 0.01010858, 0.001721674, 0.002772027, 0.007099859, 
    0.002136573, 0.005341822, 0.01117742, 0.006862058, 0.0002561405, 
    -1.897125e-07, 0.02561783, 0.006854108, 0.0249816, 0.004674013, 
    0.01185701, 0.008759394, 0.04250262, 0.01304089, 0.01182178, 0.001325945, 
    0.004388583, 0.007208937, 0.04113743, 0.006544285, 0.01342284, 
    0.002473924, 0.007297244,
  0.008484619, -0.0001602814, -3.307352e-06, 0.0006252626, -0.001906338, 
    0.001207003, 0.0006394075, 0.0003505382, 0.001574548, 2.579188e-05, 
    -4.321434e-08, 2.788787e-06, 0.001423406, 0.005964288, 0.002964397, 
    0.0001270602, 0.0006311579, 0.003077709, 2.552474e-05, 0.0005373885, 
    0.000144517, 0.0003597355, 0.004251802, 0.02338756, 0.005800686, 
    0.02757646, 3.658259e-05, 4.113937e-05, 0.001305087,
  0.01545066, 0.02076871, 0.04184645, 0.07685068, 0.003441546, 0.0005011294, 
    0.001270938, 0.0004573736, 0.0007290582, 5.636485e-06, 0.003476945, 
    0.0002774871, 0.01217278, 0.0004409428, 6.049216e-05, 0.0001336847, 
    0.0005272716, 0.0002913885, 0.0001680916, 0.0002828945, 0.0003829181, 
    0.0008602896, 0.0138432, 0.01035115, 0.04458082, 3.880098e-05, 
    -0.0001733219, 0.0008057473, 0.003163077,
  0.001940298, 0.01722957, 0.0005211148, -0.0002431657, 0.001385182, 
    0.0009255387, 0.0007299807, 7.234758e-05, 0.03175055, 0.0493583, 
    0.004032576, 0.001069129, 0.001735173, 0.005583235, 0.0001736164, 
    0.0009706343, 0.001989088, 0.002785889, 0.00766551, 0.01445401, 
    0.003155641, 0.00407041, 0.03096244, 0.03068444, 0.01836425, 0.003562296, 
    0.0002320261, 0.001032027, 0.002775326,
  1.247957e-07, 3.603162e-07, 2.02971e-08, 0.02355558, 0.003292451, 
    0.0007945132, -0.0009137032, 0.000736522, 0.0001038394, 0.001315502, 
    0.0005109546, 0.0004922295, 0.0004647936, 0.0001256488, 0.0007491893, 
    0.003093084, 0.0002945618, 0.000730648, 0.001689513, 0.002404386, 
    0.002729034, 0.0005713871, 0.07478694, 0.03804665, 7.572147e-05, 
    0.001484898, 0.009397557, 0.01111222, 7.580532e-06,
  2.922474e-07, 1.575526e-08, 7.74844e-10, 7.894675e-08, -3.155506e-06, 
    3.303199e-06, -1.570576e-05, 0.0002093404, 2.956755e-05, 0.0162231, 
    0.002633897, 0.002812806, 0.0009671858, 8.683898e-05, 9.365408e-05, 
    0.0002456777, 0.0004731007, 0.001090492, 0.009181647, 0.02041711, 
    0.0100432, 0.02590539, 0.0002451795, -0.0007541429, 0.0004908839, 
    0.0009761909, 0.01831847, 0.001075205, 2.223949e-07,
  1.120637e-07, 0.0001246781, 3.360356e-06, 0.0005726444, 0.00192326, 
    0.0009556371, -0.001047734, -0.0001700342, 0.008963003, 0.05214312, 
    0.1076139, 0.06170682, 0.124981, 0.05880692, 0.04182517, 0.05201349, 
    0.02659328, 0.02150355, 0.01202366, 0.01478801, 0.004482661, 0.1233986, 
    0.03461531, 0.01853082, 0.02976231, 0.02155306, 0.003641906, 0.008744565, 
    0.01107664,
  -0.001007097, 4.065037e-05, 0.002844848, 0.09263162, -0.0005304785, 
    8.734391e-05, 0.05776612, 0.002567277, 0.006190981, 0.05241175, 
    0.1079194, 0.05639353, 0.07282521, 0.1104873, 0.1486294, 0.1335618, 
    0.1213052, 0.08452349, 0.06631298, 0.1162594, 0.06431782, 0.1801277, 
    0.05114566, 0.08601332, 0.09338041, 0.0335667, 0.03404754, 0.04446407, 
    0.01415038,
  0.02950928, 0.1189327, 0.006445058, 0.00185038, 0.1024528, 0.01924901, 
    0.05688504, 0.08375071, 0.02190566, 0.01098132, 0.05604542, 0.1379201, 
    0.1210319, 0.1050599, 0.05596339, 0.1207871, 0.1371692, 0.1566438, 
    0.08106142, 0.1770123, 0.04132464, 0.08411826, 0.06755979, 0.275136, 
    0.2708166, 0.4269944, 0.1927885, 0.09292206, 0.07763612,
  0.07894722, 0.2689928, 0.1011153, 0.07358611, 0.1483187, 0.1019563, 
    0.09396245, 0.03501296, 0.0247207, 0.0141891, 0.01492028, 0.02537301, 
    0.0459112, 0.04472263, 0.0924693, 0.2242841, 0.1933142, 0.2155057, 
    0.03526896, 0.02226919, 0.04274565, 0.1049704, 0.2122609, 0.221553, 
    0.1746336, 0.06783, 0.03676084, 0.03565108, 0.1341589,
  0.117568, 0.07675161, 0.2696607, 0.1130827, 0.1959561, 0.166103, 
    0.08163308, 0.04009282, 0.0649803, 0.1072635, 0.1706667, 0.1666792, 
    0.1689534, 0.3048189, 0.2535306, 0.3710463, 0.2299994, 0.1645443, 
    0.2544939, 0.2573244, 0.1650264, 0.07827138, 0.05149928, 0.1577019, 
    0.1585388, 0.2632218, 0.2207877, -0.005031075, 0.1404501,
  0.5427357, 0.4045099, 0.4071528, 0.3391902, 0.3370447, 0.4025644, 
    0.4201183, 0.3536188, 0.2686018, 0.2305944, 0.3033154, 0.2352774, 
    0.209385, 0.27721, 0.2728638, 0.3028996, 0.2668005, 0.2430557, 0.2571867, 
    0.2444869, 0.273482, 0.1654882, 0.2102817, 0.2382507, 0.1115, 0.2048089, 
    0.1527269, 0.06514722, 0.1930508,
  0.1678627, 0.1660403, 0.1642179, 0.1623954, 0.160573, 0.1587506, 0.1569282, 
    0.15797, 0.1609176, 0.1638652, 0.1668128, 0.1697605, 0.1727081, 
    0.1756557, 0.1625588, 0.1684068, 0.1742548, 0.1801028, 0.1859508, 
    0.1917988, 0.1976468, 0.2175238, 0.2105506, 0.2035774, 0.1966042, 
    0.189631, 0.1826578, 0.1756846, 0.1693206,
  0.3435206, 0.2074582, 0.0917547, 0.06199342, 0.07105962, 0.1039175, 
    0.0686342, 0.05942542, 0.04563085, 0.1319624, 0.1217412, 0.1628674, 
    0.304244, -0.001567457, 0.3479778, 0.5059018, 0.4505052, 0.3544988, 
    0.2128046, 0.3413729, 0.7951277, 0.8773548, 0.229872, 0.1443555, 
    0.3568338, 0.5847996, 0.1908228, 0.1207554, 0.3021091,
  0.103822, 0.04446605, 0.08994364, 0.00945493, 0.05482014, 0.1791048, 
    0.01257741, 0.1646539, 0.2315164, 0.1971597, 0.1518155, 0.08972267, 
    0.03946423, 0.07547637, 0.1244875, 0.1871556, 0.1117982, 0.1460635, 
    0.1916492, 0.2481968, 0.3208475, 0.3567204, 0.3266383, 0.4477088, 
    0.2162937, 0.3171633, 0.2462605, 0.1052416, 0.3380346,
  0.107502, 0.1182694, 0.0748356, 0.1023211, 0.110927, 0.1391003, 0.1212165, 
    0.1153291, 0.1335319, 0.1328287, 0.1895063, 0.2148287, 0.2497061, 
    0.1602738, 0.1095956, 0.1423602, 0.1838927, 0.2698822, 0.2470685, 
    0.1959047, 0.2288469, 0.1895707, 0.1671461, 0.1013044, 0.1653921, 
    0.2450406, 0.1997919, 0.1415772, 0.1023177,
  0.1225271, 0.1219684, 0.1414015, 0.09368846, 0.1421953, 0.1588157, 
    0.2039189, 0.1199424, 0.1031395, 0.1236511, 0.09195717, 0.1081837, 
    0.06084122, 0.04439248, 0.0289978, 0.03852602, 0.0667082, 0.0606746, 
    0.07733167, 0.07525272, 0.1228214, 0.1019421, 0.09153645, 0.1037493, 
    0.03649403, 0.04072563, 0.09993331, 0.1452436, 0.17266,
  0.09010429, 0.02894817, 0.03174508, 0.03545238, 0.04962733, 0.0399679, 
    0.01610226, 0.02111104, 0.03606867, 0.07444384, 0.01466756, 0.006118368, 
    0.004141215, 0.009737704, 0.2060711, 0.02284709, 0.04657947, 0.02306504, 
    0.02743522, 0.06121329, 0.1060832, 0.0827208, 0.02065295, 0.3139559, 
    0.002692349, 0.02249524, 0.04231757, 0.02992454, 0.07810356,
  0.004581345, 0.009613549, 0.01195952, 0.0009592879, 0.001952626, 
    0.003516493, 0.0009011102, 0.004165332, 0.006887239, 0.004028664, 
    -7.697414e-06, -1.224595e-07, 0.02220201, 0.00383573, 0.02201274, 
    0.002018547, 0.006714603, 0.005284714, 0.02407569, 0.007067855, 
    0.00579477, 0.0009705744, 0.003231305, 0.00519808, 0.03259974, 
    0.002981057, 0.006214749, 0.001509177, 0.004846434,
  0.006338533, -0.0001014033, -1.676016e-06, 0.0004403905, -0.00129196, 
    0.0005752319, 0.0003170551, 0.0002625813, 0.000905765, 2.043224e-05, 
    1.326478e-08, 1.02518e-06, 0.000982002, 0.003511137, 0.001291516, 
    8.696921e-05, 0.0004457547, 0.001647346, 1.741373e-05, 0.0003012219, 
    0.0001043209, 0.000271815, 0.003205291, 0.01698317, 0.006548092, 
    0.03355116, 2.469286e-05, 2.910744e-05, 0.0009312065,
  0.01096746, 0.01083707, 0.03999568, 0.06803688, 0.001771208, 0.0003654007, 
    0.0006811355, 0.0002125366, 0.0003722118, -1.14985e-05, 0.002382468, 
    0.0001380724, 0.006040428, 0.0003407551, 4.27263e-05, 0.0001005749, 
    0.0003909158, 0.0001631478, 0.0001224609, 0.0002047288, 0.0002823586, 
    0.0006109921, 0.0100194, 0.0106525, 0.03261203, 0.0001415243, 
    -0.0005524061, 0.0005896674, 0.002313577,
  0.001363614, 0.01354, 0.00116834, -0.0002980736, 0.0009903525, 
    0.0006740148, 0.0005219693, 4.847916e-05, 0.02466422, 0.05715571, 
    0.001913785, 0.0007464711, 0.000941967, 0.002441554, 0.0001122246, 
    0.0006748317, 0.00140102, 0.001950752, 0.005350604, 0.01008794, 
    0.001701897, 0.00276138, 0.01690759, 0.02333529, 0.01508995, 0.001656036, 
    0.0001535485, 0.0007592272, 0.001934896,
  8.905176e-08, 3.62705e-07, 2.066357e-08, 0.02081543, 0.001637506, 
    0.0006110403, -0.001325941, 0.0005606069, 7.279071e-06, 0.0009734576, 
    0.0003471612, 0.0003625602, 0.0003165292, 7.477755e-05, 0.0003391108, 
    0.001474951, 0.0002165454, 0.0005103495, 0.001182869, 0.001629952, 
    0.001236862, 0.0004265002, 0.04346568, 0.02398333, 5.54413e-05, 
    0.001086874, 0.006758695, 0.007858936, 0.0002682983,
  2.918814e-07, 1.527205e-08, 7.858705e-10, 9.335067e-09, -2.172876e-06, 
    2.035955e-06, -1.815259e-05, 0.000135432, 0.0002427987, 0.007983214, 
    0.001863775, 0.001712404, 0.0006788352, 6.247398e-05, 6.925123e-05, 
    0.0001866625, 0.0001783062, 0.0005077835, 0.00697304, 0.01608856, 
    0.00559564, 0.02212299, 0.0001927327, -0.0007033144, 0.0003667511, 
    0.0007095636, 0.01348479, 0.0008559243, 2.222917e-07,
  9.156859e-08, 0.0001095508, 2.448767e-06, 0.0003495216, 0.00149493, 
    0.0008711217, -0.0009949763, -0.0005791718, 0.00828182, 0.03903207, 
    0.08134096, 0.03666338, 0.07797511, 0.03639922, 0.02710656, 0.03861362, 
    0.01682429, 0.01504403, 0.008986483, 0.01010702, 0.004180639, 0.1041077, 
    0.02701799, 0.008417611, 0.01896261, 0.01413059, 0.002792645, 
    0.006717524, 0.009638354,
  -0.0008291274, 0.0001150169, 0.001260443, 0.08737888, -0.0005201099, 
    9.543158e-05, 0.05059579, 0.002067763, 0.004328341, 0.04380441, 
    0.09083111, 0.03864837, 0.05630416, 0.08959886, 0.1178192, 0.1031498, 
    0.09232301, 0.05297667, 0.04155125, 0.1002007, 0.0568369, 0.158376, 
    0.03954619, 0.08316509, 0.07056855, 0.01864927, 0.0219278, 0.02771469, 
    0.01068631,
  0.0184871, 0.0995848, 0.003859367, 0.001237008, 0.09454516, 0.01544709, 
    0.04686432, 0.07172406, 0.01813644, 0.009190039, 0.05192384, 0.1191181, 
    0.102972, 0.07970212, 0.04662593, 0.09128135, 0.1004616, 0.1158497, 
    0.05304311, 0.1647401, 0.03586354, 0.07366917, 0.05952552, 0.2457928, 
    0.2626299, 0.4180408, 0.1476594, 0.06695928, 0.05137031,
  0.04793958, 0.2402202, 0.09286395, 0.07053337, 0.1530127, 0.09357525, 
    0.08635429, 0.03174292, 0.02056086, 0.01300882, 0.01182415, 0.04802656, 
    0.09755663, 0.0357656, 0.07841456, 0.1913223, 0.1848802, 0.1851569, 
    0.05207885, 0.02229771, 0.04268883, 0.1117381, 0.1751992, 0.2308199, 
    0.1468992, 0.05403604, 0.0271065, 0.0290582, 0.11487,
  0.09140618, 0.05851994, 0.268837, 0.08501583, 0.1831492, 0.156732, 
    0.0954042, 0.06646553, 0.08410475, 0.1313666, 0.1580993, 0.1450653, 
    0.2000827, 0.235141, 0.2210033, 0.2919485, 0.2028514, 0.1590374, 
    0.2793851, 0.2250177, 0.1684077, 0.08072317, 0.09450864, 0.1706524, 
    0.1610114, 0.2234946, 0.1985309, -0.001302142, 0.1158927,
  0.5209078, 0.3627789, 0.3178606, 0.3018006, 0.3181464, 0.3643401, 
    0.3523062, 0.296649, 0.2112464, 0.1568455, 0.2363762, 0.1874349, 
    0.1464462, 0.2202907, 0.2217072, 0.2394158, 0.2145829, 0.2094111, 
    0.2051971, 0.1815758, 0.2260998, 0.1369192, 0.1900057, 0.248222, 
    0.0944295, 0.1643284, 0.1250823, 0.04396088, 0.1504457,
  0.1657239, 0.1641073, 0.1624908, 0.1608743, 0.1592578, 0.1576412, 
    0.1560247, 0.1340892, 0.1367352, 0.1393812, 0.1420271, 0.1446731, 
    0.147319, 0.149965, 0.1570007, 0.162656, 0.1683112, 0.1739664, 0.1796216, 
    0.1852769, 0.1909321, 0.1950191, 0.1883345, 0.1816498, 0.1749652, 
    0.1682805, 0.1615959, 0.1549112, 0.1670171,
  0.2655927, 0.1419661, 0.0472956, 0.04723784, 0.02118974, 0.07737876, 
    0.02321621, 0.01201347, 0.02923124, 0.12222, 0.1072495, 0.1413529, 
    0.2914527, 0.0002364878, 0.3493153, 0.4615062, 0.4284021, 0.3527676, 
    0.1940027, 0.3432102, 0.8122711, 0.8694745, 0.2294445, 0.136015, 
    0.309002, 0.5559449, 0.1816408, 0.1155123, 0.2840378,
  0.1146098, 0.04069798, 0.08365001, 0.00917997, 0.04711748, 0.1659977, 
    0.0114861, 0.1502832, 0.2102277, 0.1857262, 0.1455943, 0.08684495, 
    0.03582209, 0.06813385, 0.1079487, 0.1628519, 0.093842, 0.124837, 
    0.1642551, 0.2187794, 0.2936334, 0.3236276, 0.3019377, 0.4237727, 
    0.1884715, 0.28892, 0.2289313, 0.09402122, 0.3068028,
  0.09108328, 0.1028285, 0.06374848, 0.08813462, 0.09443101, 0.1226762, 
    0.1043493, 0.09815966, 0.1152879, 0.113673, 0.1653798, 0.1796469, 
    0.2145526, 0.1352056, 0.09128401, 0.1218021, 0.1518903, 0.231422, 
    0.2067606, 0.1672282, 0.1917334, 0.1487295, 0.1322788, 0.08510529, 
    0.1395728, 0.2116351, 0.1685405, 0.1274622, 0.08993059,
  0.1077293, 0.102336, 0.1227538, 0.0832436, 0.1231959, 0.1286954, 0.1703071, 
    0.1000312, 0.0868428, 0.1028939, 0.0722085, 0.08635347, 0.04635758, 
    0.03476837, 0.02457434, 0.02991103, 0.0506173, 0.04381468, 0.05650987, 
    0.05929957, 0.105109, 0.07888657, 0.07061088, 0.1143686, 0.02847535, 
    0.03143284, 0.08383007, 0.1218657, 0.149367,
  0.06659991, 0.02231593, 0.02253146, 0.02284436, 0.03356376, 0.02846866, 
    0.01143351, 0.01363747, 0.02496517, 0.05159045, 0.009511461, 0.005147548, 
    0.002864032, 0.006132026, 0.2137659, 0.01678493, 0.03059226, 0.01474095, 
    0.01997634, 0.03996379, 0.07485702, 0.05830275, 0.01379813, 0.3135023, 
    0.001825748, 0.01545919, 0.02785465, 0.02186472, 0.05933117,
  0.003766846, 0.007828371, 0.02134947, 0.00072783, 0.001616583, 0.002500356, 
    0.0005353332, 0.00355917, 0.005019139, 0.00306035, -9.84027e-05, 
    -4.267001e-08, 0.02555527, 0.002627441, 0.01292065, 0.001397166, 
    0.004418245, 0.002792773, 0.01532309, 0.004280091, 0.003295352, 
    0.0008062906, 0.00265957, 0.00332702, 0.05154064, 0.00186232, 
    0.003850132, 0.001170445, 0.003897636,
  0.005315128, -5.483258e-05, -1.341328e-06, 0.0003526749, -0.001119896, 
    0.0004002772, 0.0002201003, 0.0002246431, 0.0007043471, 1.747371e-05, 
    1.357438e-08, 5.663637e-07, 0.0007753636, 0.00212348, 0.0006815835, 
    7.208055e-05, 0.0003650996, 0.001123614, 1.417424e-05, 0.0001852398, 
    8.493941e-05, 0.000226726, 0.002649121, 0.01361357, 0.02962534, 
    0.08169499, 1.942022e-05, 2.353425e-05, 0.0007566491,
  0.008866382, 0.007179236, 0.03464789, 0.09601568, 0.001103107, 
    0.0002984702, 0.00049512, 0.000141354, 0.0002657833, -0.0001885628, 
    0.001915951, 0.0001057379, 0.004017734, 0.0002827629, 2.769139e-05, 
    8.042154e-05, 0.0003192495, 0.0001162676, 0.0001013244, 0.000168714, 
    0.000230953, 0.0005004588, 0.00817239, 0.0303533, 0.05108838, 0.01097572, 
    -0.0004624985, 0.0004619575, 0.001913203,
  0.00108082, 0.01650913, 0.007146611, -0.0003089467, 0.0007913506, 
    0.0005491271, 0.0003894708, 3.939892e-05, 0.03243872, 0.07709572, 
    0.00130896, 0.0005927617, 0.0006586648, 0.001503903, 9.077131e-05, 
    0.000533317, 0.001118047, 0.001512765, 0.004261233, 0.007917577, 
    0.001211859, 0.002093638, 0.01188848, 0.02173442, 0.0706065, 
    0.0009756897, 0.0001204008, 0.000619375, 0.001538976,
  -8.812211e-06, 3.667951e-07, 2.086428e-08, 0.02877958, 0.001139191, 
    0.0005100568, 0.0005745956, 0.0003920342, -0.0002489675, 0.0007822288, 
    0.0002775085, 0.0002994307, 0.0002593228, 5.850943e-05, 0.0002345001, 
    0.0009352989, 0.0001827743, 0.0004165689, 0.0009712712, 0.001329708, 
    0.0008029321, 0.0003577349, 0.04448036, 0.02063322, 4.700482e-05, 
    0.0009038029, 0.005530082, 0.006304026, 0.008588193,
  2.934153e-07, 1.495631e-08, 7.939767e-10, 3.256252e-09, -1.623436e-06, 
    1.555473e-06, -1.363556e-05, 0.0001053374, 0.003126265, 0.004094502, 
    0.001480985, 0.001258961, 0.0005489876, 5.174215e-05, 5.918726e-05, 
    0.0001617052, 0.0001178094, 0.0002960731, 0.005869078, 0.013728, 
    0.003540926, 0.0220178, 0.0001664651, -0.0007500213, 0.0003109438, 
    0.0005953694, 0.01107309, 0.000746905, 2.25332e-07,
  9.036052e-08, 9.49327e-05, 9.525485e-06, 0.0002681714, 0.002280091, 
    0.0007327611, -0.001039618, -0.0009550444, 0.01291229, 0.03293463, 
    0.05402587, 0.02508782, 0.05153742, 0.02397069, 0.01858758, 0.02898566, 
    0.01148443, 0.01117553, 0.007451914, 0.007260366, 0.003439098, 0.1007961, 
    0.05349527, 0.004834002, 0.01277175, 0.009493232, 0.00236645, 
    0.005679023, 0.00759538,
  -0.0007457756, -4.881135e-05, 0.0004266853, 0.08384898, -0.0005295031, 
    8.308084e-05, 0.04770049, 0.001744789, 0.003409563, 0.03731623, 
    0.08830255, 0.02999488, 0.04739359, 0.07249358, 0.09573618, 0.08090512, 
    0.07504214, 0.03771344, 0.02834052, 0.09076412, 0.05145302, 0.1451784, 
    0.03732551, 0.07505014, 0.05899105, 0.01301132, 0.01637469, 0.02097428, 
    0.008278679,
  0.0140326, 0.09173896, 0.004520294, 0.001009775, 0.0889052, 0.01285301, 
    0.04312492, 0.09155571, 0.01991045, 0.01198089, 0.05536841, 0.1166397, 
    0.09407059, 0.06545312, 0.03936752, 0.07478043, 0.08020759, 0.09312557, 
    0.03980359, 0.1831474, 0.03314996, 0.06598189, 0.06013179, 0.238731, 
    0.2681215, 0.3734335, 0.1182395, 0.05111707, 0.03822898,
  0.02792633, 0.2579423, 0.1048427, 0.09434541, 0.2272681, 0.1105208, 
    0.08776563, 0.04040602, 0.02273827, 0.01807566, 0.01495829, 0.1638655, 
    0.2146869, 0.04015842, 0.07113821, 0.1831763, 0.213026, 0.1716065, 
    0.09880469, 0.028415, 0.05177865, 0.1335087, 0.1540692, 0.2508107, 
    0.1278801, 0.04526878, 0.02190161, 0.02558338, 0.1019339,
  0.0719562, 0.04955501, 0.2990637, 0.07143477, 0.1730822, 0.1519298, 
    0.1860454, 0.1871696, 0.1643564, 0.1836545, 0.215812, 0.1644193, 
    0.2917378, 0.2125709, 0.2231059, 0.2697894, 0.2126099, 0.1727122, 
    0.3138448, 0.2041121, 0.1839269, 0.1209079, 0.2020791, 0.1883244, 
    0.1563142, 0.188998, 0.2170206, 0.008855572, 0.0976756,
  0.4808082, 0.3397096, 0.2700957, 0.2774399, 0.2987178, 0.3331275, 
    0.3160846, 0.2541464, 0.1959996, 0.1105281, 0.1772856, 0.1552702, 
    0.1066127, 0.1749219, 0.1754382, 0.1945411, 0.1658424, 0.1733814, 
    0.1758757, 0.1676619, 0.1859876, 0.1305615, 0.1820834, 0.2605473, 
    0.09087302, 0.1415679, 0.112979, 0.0306756, 0.1333182,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0008435438, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -2.001011e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, -1.444806e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, -7.590593e-06, 6.592929e-06, 0, 0, 0.001982404, 0, 
    9.254623e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001298433, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, -2.785742e-05, 0, 9.776893e-05, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0.00145893, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, -0.0001037924, 4.895674e-05, 0, 0, 0.00508892, 0, 
    0.0009712941, 0, 0, 0, -1.728199e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0.000270351, 0, 0, 0, 0, 0, 0, 2.121699e-06, 0.001367004, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 3.030511e-06, -4.022265e-05, 0.002191254, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001467489, -2.994806e-05, 0, 
    0.0008767795, 0, 0, 0, 0, 0, -3.581956e-06, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, -0.0001395632, 0, 0.001114922, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3.157373e-06, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0.006540603, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0.001303692, -2.103255e-05, 0.0003070124, 0, -0.0003258779, 
    9.757477e-05, 0, 0, 0.01287108, 0.0003822081, 0.003161121, 0, 0, 
    0.0003605193, 0.000863859, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0.001949943, -5.085192e-06, 0, 0, 0, 0, 0, 2.762897e-06, 0.005215535, 
    3.526378e-07, -2.763783e-11, 0, 0, 0, -1.504594e-06, 0, 0, 0, 0, 0, 0, 0, 
    0.001217007, 0.0002292728, 0.005210803, 1.212979e-05, 0, -5.232054e-06,
  0, 0, 0, -2.694786e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0.001846019, 0.00273591, 
    -0.0001796372, -2.314633e-05, 0.002046022, 0, -6.421433e-05, 
    9.876226e-05, -5.174038e-06, 0, -6.947998e-05, 1.774412e-05, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, -0.0002765437, 0, 0.00286778, 0, 0, -1.856731e-06, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -1.780925e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001935652, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0006020511, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0.008522071, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0.001496691, 0.003616791, -3.365209e-05, 0.0008835337, 0, 
    -0.000678012, 0.0003630378, -2.53147e-05, 0.001718738, 0.02889357, 
    0.0009145281, 0.005831772, 6.325018e-05, -2.351183e-05, 0.003033654, 
    0.005084222, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0.002836386, 0.002521597, 0, 0, 0, 0, 0, -2.220276e-06, 0.01207084, 
    9.911791e-06, 6.812733e-06, 0, 0, 0, -8.104234e-06, 0, 0, 0, 0, 0, 0, 
    -6.55112e-09, 0.003438476, 0.0005153949, 0.01347112, 0.002724425, 0, 
    3.092617e-06,
  0.0004400007, 0, 0, -6.249767e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0.005789789, 
    0.005949078, -0.0001460586, -0.0001676795, 0.003558055, 5.560725e-05, 
    0.0003805835, 0.001308392, -5.695454e-05, 6.159233e-05, -5.075903e-05, 
    3.548823e-05, 0, 0, 0, -2.543307e-06, 0,
  0, 0, 0, 0, 0, 0, 0, 0.001166349, 0, 0.01117252, 0, 1.952283e-05, 
    0.0008395193, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, -2.900502e-05, -6.532268e-07, 0.0004575585, 0, 0, 
    3.821308e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0004370351, 0, 
    0.000168907, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.788681e-05, 0, 0, 
    0.005532278, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0.01301569, 0, 0, 0, 0, -9.787175e-06, 
    -8.524112e-06, 0, -5.662062e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0.003694195, 0.006238575, -7.527825e-05, 0.003759803, 0, 
    -9.862805e-05, 0.001188986, -4.700377e-05, 0.003076246, 0.04604317, 
    0.0041733, 0.007997663, 0.0005557666, 0.001210061, 0.008698504, 
    0.01504207, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0.004684248, 0.004805697, 0, 0, 0, 0, 0, 0.0004701046, 0.01603415, 
    1.818509e-05, 8.311988e-06, 0, 0, 0, -1.379802e-05, 0, 0, 0, 0, 0, 0, 
    -8.460155e-06, 0.005356101, 0.001221392, 0.03241169, 0.006246582, 0, 
    -2.849498e-07,
  0.001277295, 0, 0, -8.080542e-05, 0, -1.127493e-05, 0.0001442523, 
    4.073382e-05, 0, 0, 0, 0, 0.007664628, 0.01889618, 0.002227926, 
    -0.0002703289, 0.0053073, 0.001102102, 0.001648463, 0.004651151, 
    -0.0001303078, 0.0006945718, -0.0002565693, 4.520237e-05, 0, 0, 0, 
    -1.255116e-05, -1.565343e-05,
  0, 0, 0, 0, 0, 0, 0, 0.001765647, -4.613849e-05, 0.02925001, 0, 
    1.801898e-05, 0.004119424, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -2.533782e-06, 0, 0, 0, 0, -4.683336e-05, 0.00120357, 0.001265531, 
    0.0001002396, 4.026946e-06, 0.000145218, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -1.723833e-05, 0.0002447916, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0005768602, 0.0002179491, 0, 0.0009524387, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.0005612781, 0, -2.610617e-06, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6.210371e-06, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001075468, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, -1.348966e-06, 0, -9.423438e-06, 0, 0, 0, 0, 0, 0, 0, 0, 
    -8.855031e-06, -4.651165e-05, -3.054367e-05, 0.002846459, 0.001405079, 
    0.005094715, 0.0003181653, 0, 0, 0, -1.958369e-05, -5.817689e-10, 0, 
    0.000372041, 0,
  0, 0, 0, 0, 0, 5.867727e-05, 0, 0, 0.0001279287, -6.485749e-06, 0, 0, 0, 0, 
    0, 0.0005961849, 0, -5.212975e-05, 0.01013592, -5.719885e-06, 0, 0, 0, 0, 
    0, 0.0003200835, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -5.771632e-05, 0, 0.02151337, 0, 0, 0, -1.385242e-07, 
    0.0002472378, 0.0004229835, 0, -9.790222e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0.006008263, 0.009534256, -0.0001407975, 0.006347116, 0, 
    0.00118189, 0.002191508, 0.0001215166, 0.003740117, 0.06477649, 
    0.00856834, 0.01222413, 0.0006500771, 0.005119934, 0.01454386, 
    0.02047109, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0.008201114, 0.008818529, 0, 0, 0, 0, 0, 0.0005034181, 0.02217181, 
    0.0003296761, 0.001224398, -7.991061e-06, 0, 2.731535e-06, -2.510422e-05, 
    0, 0, 0, -6.459797e-06, 0, 0, -6.593174e-05, 0.01062076, 0.006912716, 
    0.04330582, 0.007294037, -1.961352e-05, 5.646644e-06,
  0.002786364, 0, 0, -3.194189e-05, 0, -1.415878e-05, 6.278835e-05, 
    -1.832989e-05, -1.227919e-05, 0, 0, -3.663169e-05, 0.01059381, 
    0.03113719, 0.01628347, 0.004504145, 0.008516057, 0.007304003, 
    0.003629498, 0.01187708, -0.0003073437, 0.006013901, 2.25961e-05, 
    0.0001831657, 0, 0, 0, -2.839563e-05, -7.626382e-05,
  0, 0, 0, 0, 0, 0, 0, 0.006410779, 6.629464e-05, 0.05980246, 0, 
    4.498586e-05, 0.008942598, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.122743e-05, 
    0, 0, 0, 0, 0,
  0, 0, 0.001177962, -3.103169e-07, 0, 0, 0, -0.0001225511, 0.003524208, 
    0.002802066, 0.002982395, 5.074692e-05, 0.0007203048, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, -6.382292e-05, 0.003843767, 0, 0, 0, 0,
  0, 0, 0, 0, 0.000422892, 0.0001202762, 0, 0, 0, -2.411982e-05, 0.002478995, 
    0.0006171159, -7.875378e-05, 0.001980276, 0, 0, 0, 0, 0, 0, 0, 
    7.435808e-05, 0.004019798, 0.004062449, 1.206067e-06, 0.00219477, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.095224e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.001974163, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0.001588002, 0, -7.296675e-06, -2.55001e-05, -1.573951e-05, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.003974232, 0.001858223, 0.0004934801, 0, 0, 
    0, 0, 0, 0, 0,
  0, 0, 0, -2.430704e-05, 9.377178e-05, 0.0001429798, 0, 0, 0, 0, 0, 0, 0, 0, 
    -3.932654e-05, -0.000286057, 0.001964875, 0.00822238, 0.00467738, 
    0.01830866, 0.006925981, 0, 0.0007439548, 0, 0.003881555, -3.769415e-05, 
    0.000169417, 0.005089737, 0.004209477,
  0, 0, 0, 6.459094e-06, -2.728043e-05, 0.0008318876, -2.587338e-05, 0, 
    0.002184505, 0.0001564752, 0, 0, 0, -2.814762e-06, 0.002791567, 
    0.002492324, -4.509372e-05, 0.004718069, 0.01314084, -4.04594e-06, 0, 0, 
    0, 0, -2.581647e-08, 0.00574611, -2.34887e-05, -9.417404e-08, 0,
  0, 0, 0, 0.0006784907, 0.0002009048, -2.751149e-05, -0.0001283074, 0, 
    0.03508357, 0, 0, 0, -8.683813e-06, 0.002271348, 0.001340494, 0, 
    0.0001946373, 9.153078e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -2.730543e-05, 0.007832233, 0.01586004, -0.0001560149, 0.01303495, 
    0.0002776744, 0.00753968, 0.005939492, 0.000139891, 0.006159948, 
    0.1014604, 0.01814079, 0.02279996, 0.003473581, 0.006062543, 0.02089174, 
    0.03046695, -4.34253e-05, 0, 0, 0, -1.005494e-05, -1.407277e-05, 0, 
    -1.625481e-06, 0, 0,
  0.0009934941, 0.01909017, 0.01336561, -9.061141e-06, 0, -2.437114e-06, 
    -1.3396e-05, -7.268581e-06, 0.002193452, 0.02990128, 0.005637256, 
    0.004145563, 0.0002648954, -1.994712e-06, 9.704057e-05, -4.584328e-05, 0, 
    -3.290486e-09, 0, -6.918219e-05, 0, -3.226129e-05, 0.0004665073, 
    0.02100987, 0.01474127, 0.0597381, 0.0128477, 3.324792e-05, 0.005754595,
  0.004855108, -6.069427e-05, 0.0004414243, -0.000207748, 9.08006e-05, 
    -3.154311e-05, 0.0008181523, 0.0006402395, 0.00225586, 0, -7.108636e-05, 
    -0.0001958506, 0.02415795, 0.04310983, 0.05926545, 0.0208594, 0.01533645, 
    0.01144536, 0.01198727, 0.0238053, 0.0001991821, 0.009593213, 
    0.006156178, 0.004772654, -1.470697e-05, 0, -4.842555e-06, -0.0001156525, 
    -0.0001284122,
  0, 0, 0, 0, 0, 0, 0, 0.01906594, 0.002808877, 0.09808741, 1.077471e-05, 
    0.002034115, 0.01500047, 0, 0, -2.879786e-05, 0, 0, -8.923794e-05, 
    -6.675278e-06, 0, 0.0002316796, 0, -9.113779e-05, 0, 0, 0, 0, 0,
  0, -3.32792e-05, 0.002994912, 6.691064e-05, -2.416373e-05, 0, 0, 
    -0.0002091226, 0.005226575, 0.004523539, 0.008908737, 0.00549597, 
    0.01197713, 0, 0, 0, 0, 0, 0, 0, 0, -9.286769e-06, -5.204286e-06, 
    -0.0002560601, 0.01082792, 0, 0, 0, 0,
  0, 0, 0, 0, 0.00358485, 0.003995913, 0.0006911465, 0, 0, 5.4908e-05, 
    0.007935409, 0.003018325, 0.005536237, 0.005022572, 2.580768e-07, 
    0.000620444, -1.918033e-05, 0, 0, 0, 0, 0.008382888, 0.01260184, 
    0.006573016, 0.0005378321, 0.0053666, 0, 0, 0,
  0, 0, 0, 0, 0, -1.576516e-05, 0, 0, 0, 0, -2.771948e-06, 0.001271383, 
    -0.0001005365, 0, -7.719148e-07, 0, 0, 0, 0, 0, 0, 0.003172147, 
    -3.923869e-05, 0, 0, -9.481671e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, -1.051537e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0.0007920325, -9.052118e-07, 0, 0.0006421793, 0.003682868, 0, 
    -2.430705e-05, 0.0004324147, -4.719633e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -5.061424e-06, 0.004913496, 0.004817642, 0.004053692, 0.0002161455, 0, 0, 
    -1.799228e-05, -2.124654e-06, 0.0001420991, 0.001230328,
  0.001237265, 0, -7.518534e-06, -4.643337e-05, 0.003524243, 0.0006404227, 
    0.0004326888, 0, 0, 0, 0, 0, 0, 0, -0.0002559589, 0.002521352, 0.0140961, 
    0.01237499, 0.01713366, 0.03009421, 0.02980798, 0.0006031835, 0.00502754, 
    0, 0.008002508, -3.550404e-05, 0.002997084, 0.008522555, 0.007607213,
  0, 0, 0, 0.001555703, 0.004037387, 0.002123947, 0.0004939623, 0, 
    0.00938158, 0.003276532, 0, 0.0003035473, -1.921734e-05, 0.001916413, 
    0.02955923, 0.01370479, 0.00474137, 0.0204991, 0.02774597, 0.002056108, 
    0.0009414319, -6.239547e-05, 0, 0, -2.137434e-05, 0.01730848, 
    6.206345e-05, -0.0001214332, 0.0001691795,
  1.002595e-09, 0, 0, 0.01083201, 0.002115031, -5.014617e-05, -0.0002035619, 
    -2.206479e-10, 0.0490889, 4.191573e-05, 5.380381e-09, 0, -3.312181e-05, 
    0.00989694, 0.00921376, -6.266294e-06, 0.0004435382, 0.0001546625, 
    0.0001487566, -3.131861e-07, 0, 0, 0, 0, 0, -4.511813e-08, 0, 0, 0,
  0, 0, 0.0003858451, 0.008290704, 0.02767733, 0.0004060964, 0.0183977, 
    0.002402921, 0.0403429, 0.01883677, 0.005812387, 0.01015313, 0.1290225, 
    0.03811304, 0.03672654, 0.02042152, 0.01279109, 0.02558993, 0.03965452, 
    -8.512149e-05, 0, 0, 0, 0.001429002, 0.0009409648, 0, 0.000210896, 
    0.0003896926, 0,
  0.008358386, 0.0434338, 0.0236457, 5.203615e-05, -2.249831e-06, 
    0.001013899, 0.003076472, 0.0006388245, 0.03203106, 0.05982117, 
    0.01154582, 0.01080707, 0.007467825, 0.01119618, 0.003360366, 
    -0.0001417948, -4.763041e-06, 0.0001724913, 0, -0.0001467448, 0, 
    -7.954297e-05, 0.007879901, 0.06428048, 0.02925479, 0.07801359, 
    0.01853566, 0.005522738, 0.01399794,
  0.02134056, -0.0001340102, 0.003776275, 0.004588521, 8.714528e-05, 
    0.0006241638, 0.004747313, 0.008117883, 0.005959873, -1.765571e-05, 
    -0.0001359863, 7.917858e-05, 0.07879113, 0.08100503, 0.1118043, 
    0.05044308, 0.02060483, 0.02053484, 0.02039088, 0.04826133, 0.01301667, 
    0.01621031, 0.02797087, 0.0286644, 0.000256488, 0, -3.849066e-05, 
    -0.0002268447, 0.006053491,
  -9.635293e-10, 1.19971e-08, 0, -2.09514e-06, 0, 0, 0, 0.04270577, 
    0.01716579, 0.1470471, 4.846174e-05, 0.006025424, 0.03683487, 
    -1.440788e-05, 0.0001456205, 0.001807, 7.687649e-06, -7.118013e-05, 
    0.001045953, -3.67705e-05, 3.092585e-08, 0.001338469, 0, 0.001756359, 
    0.0002499999, -1.712916e-10, 0, 0, 0,
  0, -8.628864e-05, 0.00541651, 0.00155262, 0.0005148094, 0, 0, 0.0001667841, 
    0.0122905, 0.01270711, 0.02004018, 0.0161245, 0.02237709, -0.0001120043, 
    -2.91866e-08, 0, 0, -1.858133e-05, 0, 0, 0, 0.001240491, 0.0001965587, 
    -0.000351513, 0.02452689, 0, 0, 0, 0,
  0, 0, 0.00136691, -1.110435e-05, 0.009564799, 0.008757615, 0.004927643, 0, 
    -1.035843e-05, 0.002327809, 0.01611856, 0.01206518, 0.02190142, 
    0.02049533, 0.002585091, 0.004131653, 0.000583382, 0, 0, 0, 
    -2.036467e-05, 0.02020967, 0.02578717, 0.01124259, 0.005236345, 
    0.00724966, -1.893435e-05, 0, 0,
  0, 0, -1.411527e-08, 0, 0, -0.0001140241, 0, 0, 0, 0, 1.264611e-05, 
    0.002122991, 0.004933392, -8.166523e-07, 0.001179489, -3.392432e-05, 
    0.0001951702, 0, 0, 0, -4.216807e-05, 0.006038473, 0.0002646449, 
    -5.166661e-05, 0, 0.0008734883, -1.965521e-05, 0, 6.626819e-05,
  0, 0, 0.001803833, 0, 0.003937283, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0.0001308004, 0, -9.513731e-06, 0.001230021, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.003943308, 0.0007539084, -3.993326e-05, 0.002443929, 0.01136073, 
    -0.000135875, -0.0001084721, 0.00116787, -0.0001335494, 0, 0, 
    0.002758504, 0, 3.558867e-05, 0, 0.001907713, 0, 6.851097e-05, 
    0.001131737, 0.006221392, 0.01234336, 0.009247988, 0.0007468873, 
    -1.078151e-05, 0, 0.0002347823, 0.00342007, 0.002515017, 0.009472914,
  0.01504056, 0.00197174, 0.000428791, -4.109428e-05, 0.01103132, 0.00254137, 
    0.003198919, 0, 0, -2.231892e-06, -1.752866e-05, 0, -5.454265e-06, 
    0.001831422, 0.0006592167, 0.01661895, 0.02452275, 0.02187148, 
    0.03258331, 0.06757554, 0.05075476, 0.006816341, 0.01079935, 
    -8.496261e-06, 0.01552876, 0.002349822, 0.006100295, 0.02448243, 
    0.01210555,
  7.715498e-06, -1.171009e-10, 0, 0.01124507, 0.02486716, 0.009231417, 
    0.001202197, 0.0009703205, 0.04179471, 0.02583166, 0.002508036, 
    0.001767252, -0.0001649111, 0.00945221, 0.06477445, 0.03861239, 
    0.01918309, 0.04326322, 0.05763979, 0.01326669, 0.02462847, 0.004491925, 
    0.004358579, 0.0003943116, -5.505417e-05, 0.02725083, 0.001114155, 
    0.0003658013, 0.0006217443,
  2.912183e-06, 0, 0, 0.02961565, 0.01247605, 4.408491e-05, -0.0003307966, 
    0.002283286, 0.05442157, 0.03085829, 0.0003344529, 6.814633e-06, 
    0.0006335719, 0.02822547, 0.04981066, 0.007806363, 0.002416778, 
    0.00291906, 0.002322916, 0.001457856, -1.197707e-05, 0, -1.203266e-06, 
    8.265009e-06, 3.807797e-05, -1.131316e-05, -4.036602e-06, 0.001210721, 
    -1.876375e-08,
  5.211541e-07, 0.001720386, 0.0005954383, 0.009697094, 0.06916784, 
    0.02458874, 0.03234909, 0.05861213, 0.145759, 0.1294782, 0.02217033, 
    0.01439407, 0.1928238, 0.1358089, 0.1257984, 0.1261467, 0.02936834, 
    0.03161494, 0.04909264, 0.0006907737, 1.875223e-08, 4.101848e-07, 
    -3.138567e-07, 0.008999054, 0.01565718, -1.152348e-07, 0.0001266661, 
    0.001148171, 3.850444e-06,
  0.1011103, 0.08777632, 0.101929, -0.0001254619, 0.008807051, 0.001833814, 
    0.0546245, 0.02348033, 0.1509359, 0.1636408, 0.1052351, 0.0712256, 
    0.08593753, 0.02397348, 0.07542034, 0.02023567, 0.008797633, 0.01823331, 
    -1.795196e-05, 0.01471351, 1.506369e-05, 0.004103914, 0.03276119, 
    0.1866117, 0.1225342, 0.1119988, 0.05334684, 0.0447367, 0.03917241,
  0.1302597, 0.02500865, 0.0102862, 0.00484126, -3.409624e-05, 0.0437056, 
    0.09133518, 0.1215205, 0.1079734, 0.001276186, 0.001395614, 0.02030566, 
    0.2656976, 0.2263752, 0.2544712, 0.1682374, 0.0464344, 0.03038073, 
    0.03856134, 0.09280287, 0.06659056, 0.05181409, 0.05543597, 0.1411341, 
    0.00697902, -3.08483e-06, -5.70042e-05, 0.0004535461, 0.0515147,
  0.0001361253, -2.800947e-05, -1.358026e-07, -1.393081e-05, -5.154991e-05, 
    -9.995931e-06, 5.106375e-05, 0.06637701, 0.0797088, 0.3010242, 
    0.02659977, 0.04283214, 0.09501267, 0.001491204, 0.006935111, 0.00894355, 
    0.0001269626, 0.001961858, 0.01260248, 0.006407439, 0.0001765883, 
    0.004086768, -7.438193e-06, 0.01387371, 0.00129027, 5.047341e-05, 
    4.014553e-05, -4.819684e-07, 5.018029e-05,
  0, 0.00355829, 0.006591185, 0.007708103, 0.0003443218, 3.472499e-05, 
    0.0001162944, 0.0004121196, 0.02861292, 0.03575466, 0.06317107, 
    0.03488629, 0.04414171, 0.001832628, -4.640558e-06, 0.001017539, 
    0.0001474581, -8.402165e-05, 0, 0, 0, 0.005044438, 0.003536534, 
    0.001616624, 0.03323071, 1.650518e-05, 0, -2.244826e-06, 0,
  0, -2.769175e-05, 0.004671228, 0.0008012746, 0.01855345, 0.01604439, 
    0.005879204, 0, -2.367281e-05, 0.005961284, 0.0222869, 0.02454948, 
    0.04609703, 0.03779357, 0.0179056, 0.02086285, 0.003443234, 
    -5.886615e-06, 0, 0, -0.0001168433, 0.04076837, 0.05305118, 0.02276423, 
    0.02441303, 0.01361672, 0.0003138312, 0, 0,
  0.0006601498, 0.001482667, 0.0003742932, -9.484377e-06, -4.033804e-06, 
    0.0007305719, 0.0002832904, -2.972835e-06, 0, 0, 0.001295908, 
    0.006139582, 0.01048214, -3.182957e-05, 0.007548373, 0.003684157, 
    0.0002952855, 0.0003443196, 0, 0, -0.0001865496, 0.007291077, 
    0.0007620105, -9.443827e-05, 0, 0.005995431, 0.008448829, 0.001655437, 
    0.005702548,
  0.0004206307, 0, 0.003756146, -3.652234e-06, 0.00736874, -2.877407e-05, 
    -7.22082e-05, 0, -1.797918e-05, 0, 0, 0, 0, 0, 0, 0, 0, -6.418403e-05, 0, 
    0, 0, -1.466847e-05, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  -4.30372e-06, -4.56835e-06, -5.408407e-06, 0.003232097, 0, 1.120737e-05, 
    0.00413775, 0, 0, 0, 0, 0, 0, 0, 7.825597e-06, 0, 0, 0, 0, 0, 
    0.0001530236, 0, -1.812997e-05, -9.049274e-07, 0, 0.0003056377, 0, 0, 0,
  0.01862401, 0.004776263, -0.0001644459, 0.008845696, 0.01662272, 
    -0.0003962476, 0.002551646, 0.00335468, 0.001518557, 0.001057893, 0, 
    0.006390765, 0, 0.001090701, -4.715312e-05, 0.001879124, 0.003402328, 
    0.002197774, 0.003491604, 0.009448539, 0.01785463, 0.02218246, 
    0.008617689, 0.001767136, 0.0005369981, 0.002362968, 0.0122686, 
    0.01309852, 0.01937572,
  0.02361862, 0.004777186, 0.001774645, 0.0007603476, 0.01811567, 
    0.004717567, 0.008370222, 0.002003264, 0.001348256, -0.0001458426, 
    0.002988444, -6.054016e-05, 0.001116115, 0.003706408, 0.005956463, 
    0.03120063, 0.04233935, 0.03828433, 0.05677946, 0.1240561, 0.08477116, 
    0.02352053, 0.01755651, 0.004709078, 0.02403564, 0.01118954, 0.0128292, 
    0.04281505, 0.02158566,
  0.001587609, 0.0004228721, -1.654868e-09, 0.02019363, 0.05652503, 
    0.02591689, 0.004710606, 0.001660441, 0.06098573, 0.03930027, 0.01699035, 
    0.01450633, 0.001694826, 0.02427367, 0.1239334, 0.1254515, 0.0765598, 
    0.08697278, 0.1331928, 0.08957397, 0.05561985, 0.05176578, 0.016134, 
    0.00640127, 0.001942937, 0.03952376, 0.01069769, 0.003645213, 0.00250952,
  8.117926e-05, 5.894836e-06, 2.789202e-06, 0.1012498, 0.1152097, 0.07858949, 
    0.04158244, 0.02842141, 0.0633781, 0.08256029, 0.01326834, 0.00138721, 
    0.002197284, 0.08265317, 0.1376887, 0.04675123, 0.03251217, 0.07748754, 
    0.133783, 0.03169583, 0.002085281, 0.006265899, 0.0003184878, 
    0.004743835, 0.01154815, 0.000520956, 0.003973361, 0.03615593, 0.002770887,
  1.899839e-05, 0.0325122, 0.003381829, 0.01410337, 0.1220189, 0.07576384, 
    0.04698183, 0.07481112, 0.1272107, 0.09570815, 0.03318651, 0.01599363, 
    0.1804536, 0.1163466, 0.1281082, 0.1400525, 0.05219084, 0.04337279, 
    0.07533287, 0.002883046, 3.720128e-07, 1.243409e-05, 0.008660612, 
    0.1338442, 0.09655017, 0.0009830989, 0.003498956, 0.0003749614, 
    0.0005135423,
  0.1805414, 0.3834306, 0.2892654, 0.002110828, 0.01726526, 0.0269544, 
    0.06983897, 0.06398264, 0.3410903, 0.3567291, 0.07519779, 0.06274719, 
    0.08516073, 0.01845262, 0.08151373, 0.0167487, 0.003571082, 0.009773645, 
    0.0001496027, 0.0146023, -8.874826e-05, 0.001977132, 0.1426113, 
    0.3949066, 0.2179141, 0.1328175, 0.06001104, 0.07861065, 0.03179315,
  0.248963, 0.1512488, 0.0847931, 0.007021572, 0.002572011, 0.05996932, 
    0.07801598, 0.1036227, 0.08254472, 0.0008772893, 0.002967853, 0.01311284, 
    0.2105209, 0.2075463, 0.2547926, 0.2157255, 0.1211381, 0.06123814, 
    0.07285358, 0.1334652, 0.1179776, 0.04085372, 0.153846, 0.3066095, 
    0.01760153, 0.0101395, 0.002720647, 0.006798595, 0.4052756,
  0.02654097, 0.001682547, 2.811542e-05, 0.0302464, 0.05260284, 3.012158e-06, 
    0.01682975, 0.05624728, 0.2098901, 0.2843025, 0.1195113, 0.08773912, 
    0.1135919, 0.034638, 0.01299096, 0.09043562, 0.05637239, 0.1212425, 
    0.1261064, 0.1303869, 0.05362591, 0.009850185, 0.02063195, 0.1646753, 
    0.2442187, 0.04780721, 0.03357274, 0.02043041, 0.07403201,
  -3.677079e-05, 0.009804343, 0.01191485, 0.02335578, 0.001731745, 
    0.001369449, 0.004507517, 0.002444474, 0.07485253, 0.2629447, 0.2313523, 
    0.1529801, 0.1088586, 0.08015359, 0.04761204, 0.01369802, 0.01447591, 
    0.002081226, 0, -9.503259e-06, -8.163657e-07, 0.0193945, 0.02314742, 
    0.01521448, 0.09022103, 0.0144776, -8.637806e-05, 2.652956e-05, 
    -4.140746e-06,
  3.53857e-05, 0.0002076838, 0.005256198, 0.003015874, 0.03238023, 
    0.02396796, 0.01038409, 0.0008575984, 4.085221e-05, 0.01355296, 
    0.0403089, 0.0453329, 0.1380614, 0.1416277, 0.05975276, 0.03595531, 
    0.01476272, 0.009581969, 0.003990573, 0.001608573, -0.0001247999, 
    0.05991792, 0.08253413, 0.03837823, 0.04492595, 0.02715989, 0.002701053, 
    -1.652045e-09, 0,
  0.003729359, 0.001507387, 0.002360814, -0.0002592327, 0.0007923829, 
    0.009230505, 0.005105645, 8.367473e-05, 0, -5.593109e-05, 0.003887543, 
    0.0109446, 0.01797283, -0.0001256635, 0.01217148, 0.006698436, 
    0.005201454, 0.006343124, 4.104209e-07, 0, 0.001603584, 0.01329511, 
    0.001840632, -0.0001852276, -2.455793e-05, 0.009355704, 0.01391295, 
    0.002199959, 0.01188478,
  0.001834362, 0.0005235684, 0.004715757, 0.005505602, 0.01521299, 
    0.00127368, 0.0003636025, 0, -7.71367e-05, 0, 9.962424e-07, 
    -3.969627e-06, -2.809856e-05, 0, 0, 2.652377e-06, -1.51477e-09, 
    -6.418541e-05, 0, 0, -8.342485e-05, -0.0003701307, 0, 0, 0, 
    -5.768066e-05, 0, 0, 0,
  0, 0, 0, 3.909432e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.704968e-05, 
    0, 0, 0, 0, 0, 0, 0, 0,
  -6.215712e-05, 0.001499712, -2.909181e-05, 0.01087096, -0.0001026557, 
    0.004458282, 0.008911831, -2.930287e-07, 0, -5.892711e-05, 0, 0, 
    8.299665e-05, -5.608098e-06, 0.001094377, 0, 0, 0, -0.0001505774, 
    -4.36454e-05, 0.0009034283, 0.001956812, 0.004237803, -1.678475e-05, 0, 
    0.001663111, -0.000339237, 0, 0,
  0.0418538, 0.01888737, 0.0006715463, 0.01841103, 0.02422435, 0.004706485, 
    0.007906446, 0.01072316, 0.009339978, 0.005822842, 0.0008738823, 
    0.01159364, -4.503167e-05, 0.004199545, 0.003511364, 0.001896781, 
    0.01139439, 0.01202265, 0.006416208, 0.01516449, 0.03507366, 0.04410539, 
    0.0390199, 0.02033998, 0.02408611, 0.007380153, 0.02009036, 0.02201501, 
    0.0319507,
  0.03644618, 0.01085778, 0.007684646, 0.003670875, 0.06210542, 0.01977552, 
    0.01814441, 0.003433441, 0.00751982, -0.0002547731, 0.01153236, 
    0.003825194, 0.005480387, 0.008225718, 0.01641717, 0.05174666, 0.0581951, 
    0.05510803, 0.09448641, 0.2189323, 0.1757169, 0.08280542, 0.03491207, 
    0.02273963, 0.0490294, 0.03916759, 0.04860064, 0.07203641, 0.05149677,
  0.03745533, 0.01483689, 0.0005171581, 0.0407424, 0.1316921, 0.07729007, 
    0.04577137, 0.0297111, 0.1297184, 0.1238486, 0.0727997, 0.05725698, 
    0.009765974, 0.06234298, 0.1645258, 0.1834479, 0.111967, 0.1679082, 
    0.2674425, 0.2152512, 0.1066215, 0.08589166, 0.02122505, 0.03037727, 
    0.02758166, 0.08449346, 0.0840481, 0.05474764, 0.02516064,
  6.50987e-08, 8.756494e-07, 8.996863e-05, 0.1260285, 0.1201134, 0.07045999, 
    0.03268864, 0.02752351, 0.06787967, 0.08248049, 0.01102081, 0.001009907, 
    0.006971046, 0.09219441, 0.1139549, 0.03222403, 0.03392656, 0.06122708, 
    0.08722308, 0.02430438, 0.0001281328, 0.003040557, 5.522613e-05, 
    0.001136482, 0.001663727, 0.009649187, 0.00325587, 0.03275318, 
    -0.0002938178,
  8.43328e-06, 0.03314577, 0.002863374, 0.01588481, 0.09625786, 0.03721317, 
    0.03859133, 0.04247729, 0.1136065, 0.08432756, 0.02867633, 0.0122771, 
    0.1558238, 0.09820829, 0.1041513, 0.1055761, 0.03795283, 0.04099642, 
    0.06651571, -4.069389e-05, 1.26976e-08, 5.226259e-06, 0.02291049, 
    0.06886232, 0.06897744, 0.0001041032, 0.001847189, 2.405088e-05, 
    2.956308e-05,
  0.1283988, 0.3638692, 0.2089197, 0.0009393782, 0.01013693, 0.01749909, 
    0.06030108, 0.0239791, 0.2399564, 0.3027828, 0.04488514, 0.04359288, 
    0.05989435, 0.01865581, 0.05865848, 0.01122997, 0.002306666, 0.003459369, 
    0.0001075969, 0.009770254, 2.453217e-06, 7.651645e-05, 0.08230302, 
    0.3491469, 0.1547917, 0.1222976, 0.05583498, 0.04638572, 0.01126917,
  0.2295668, 0.1173226, 0.07553115, 0.1127874, 0.00223006, 0.03395331, 
    0.04517128, 0.08410587, 0.05926505, 0.001447056, 0.004033721, 
    0.007443869, 0.1683879, 0.1744439, 0.2149743, 0.1598789, 0.09201969, 
    0.06688207, 0.04725149, 0.1129903, 0.08877172, 0.02749453, 0.1273391, 
    0.2707722, 0.01315305, 0.00486964, 0.002115792, 0.002214308, 0.3564757,
  0.02045912, 0.01834071, 0.0238007, 0.03681982, 0.1019197, 0.03904048, 
    0.009406361, 0.04195248, 0.1544421, 0.2494233, 0.1060691, 0.06413461, 
    0.08799456, 0.03272069, 0.001314291, 0.06970803, 0.06774965, 0.09788384, 
    0.1533646, 0.1004013, 0.03680728, 0.01197614, 0.009526904, 0.1218008, 
    0.2419144, 0.03188302, 0.05522252, 0.06396683, 0.094653,
  0.0210709, 0.02566588, 0.01982175, 0.0784208, 0.03823185, 0.05201206, 
    0.05624462, 0.006000862, 0.1226604, 0.2336524, 0.2203045, 0.1642339, 
    0.1198724, 0.09986196, 0.07340924, 0.06576422, 0.1100324, 0.03141422, 
    0.03272158, 0.01214262, 0.003263008, 0.07500686, 0.09550542, 0.1264987, 
    0.1558593, 0.1281515, 0.09618384, 0.04134053, -0.000773216,
  0.001984027, 0.002017976, 0.01160019, 0.008441082, 0.06301245, 0.1049607, 
    0.01826675, 0.0632255, 0.033018, 0.051524, 0.0775168, 0.08225985, 
    0.2096007, 0.2503883, 0.1654952, 0.1312724, 0.1298176, 0.08241516, 
    0.0325237, 0.005942704, 1.974698e-05, 0.07671845, 0.1355153, 0.09599047, 
    0.1390974, 0.1044405, 0.05427619, 0.01217419, 0.004981146,
  0.008854148, 0.001410244, 0.006405801, 0.002122483, 0.006359065, 
    0.02037497, 0.01976559, 0.002190505, 7.893405e-05, 0.0007549336, 
    0.01561965, 0.02095595, 0.03465687, 0.01537208, 0.02072989, 0.02696069, 
    0.0353156, 0.0404917, 0.0007393713, 0, 0.004598617, 0.02339156, 
    0.006292083, 6.183871e-05, 0.0002594387, 0.02186566, 0.04832523, 
    0.01527636, 0.02096386,
  0.008919569, 0.002550677, 0.008531469, 0.007610702, 0.0180878, 0.007251919, 
    0.0007966688, 0, 0.0002557789, 0.0001651212, 0.0002297128, 0.004157257, 
    0.003358552, -4.382171e-05, 0, -1.394175e-05, 0.0001076924, 0.0009885905, 
    0, -2.682464e-06, -9.918554e-05, 0.001413917, 0, -1.750118e-05, 0, 
    0.007287077, -2.351397e-05, 0, -3.80844e-05,
  0, 0, 0, -0.0001483699, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001311723, 0, 
    0, 0, 0, 0, 0, -0.0003667788, 0.0004377735, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.587294e-05, 0, 0, 0, 0, 0, 0, 0, 
    -5.225478e-05, 0.001035172, 0, 0, 1.840193e-05, 0, 0, 0, 0,
  0.002142405, 0.01465419, 0.006878418, 0.0201918, 0.001945122, 0.004603112, 
    0.01129744, 0.003273274, -2.332718e-11, -0.0001297826, 2.9733e-05, 
    2.83761e-05, 0.001214748, -1.99842e-05, 0.002620884, 0.00063448, 
    0.0008369559, 0.0001548619, -0.0004330438, 0.0002753368, 0.005758597, 
    0.003506985, 0.01432706, 0.003671353, 0.001667691, 0.006291527, 
    0.003111708, -1.951659e-05, 0.001003659,
  0.0755319, 0.09639406, 0.04713617, 0.05464653, 0.07592478, 0.06337512, 
    0.04190349, 0.0274113, 0.02366704, 0.01848, 0.004868689, 0.03216538, 
    0.001458182, 0.01349903, 0.018101, 0.01210769, 0.02171056, 0.03280677, 
    0.02475846, 0.02749847, 0.06594574, 0.09001022, 0.1417068, 0.05990169, 
    0.05702295, 0.05018701, 0.06861733, 0.05038919, 0.0683909,
  0.1037458, 0.1172947, 0.1013308, 0.1075261, 0.1618028, 0.05853869, 
    0.07666152, 0.05543341, 0.03070425, 0.05382542, 0.06072588, 0.05893859, 
    0.02888123, 0.02429621, 0.04883641, 0.09142739, 0.08980016, 0.0845984, 
    0.13714, 0.2848781, 0.2092932, 0.1326645, 0.1260028, 0.07184578, 
    0.1171836, 0.0977855, 0.08740726, 0.1386599, 0.1757234,
  0.02250515, 0.01364046, 0.0206378, 0.08664843, 0.1379973, 0.08811385, 
    0.07730216, 0.06651896, 0.1596892, 0.1324776, 0.1080492, 0.07468833, 
    0.04346212, 0.07461138, 0.1911287, 0.1277584, 0.1071177, 0.1459627, 
    0.2461452, 0.1638813, 0.1013443, 0.08227019, 0.01591455, 0.03402202, 
    0.0245358, 0.09192459, 0.07474453, 0.06980375, 0.02311169,
  4.266354e-06, 5.200968e-07, 0.0005738869, 0.129728, 0.1390449, 0.05035182, 
    0.0299089, 0.03749636, 0.06465202, 0.06481201, 0.01491557, 0.00263008, 
    0.01002027, 0.08519769, 0.09972282, 0.02609514, 0.0417921, 0.04703545, 
    0.04821715, 0.009654612, 0.0001158046, 1.600602e-05, 2.970143e-06, 
    4.344287e-05, 0.002121991, 0.004886121, 0.002038479, 0.007753292, 
    0.001665867,
  1.227711e-05, 0.02459329, 0.00105118, 0.02638296, 0.0853611, 0.02524078, 
    0.04502491, 0.03179168, 0.112589, 0.07788254, 0.02546905, 0.0174769, 
    0.1486143, 0.09127007, 0.09160227, 0.08710277, 0.04052741, 0.04674056, 
    0.06216817, -0.0001974058, 3.306655e-08, 2.742542e-06, 0.01941254, 
    0.04099698, 0.05389579, 0.0001416189, 0.001502683, 9.987263e-06, 
    5.576328e-06,
  0.09960101, 0.3889594, 0.181948, 0.001891098, 0.006071324, 0.01274861, 
    0.0536112, 0.02240872, 0.1942828, 0.2804302, 0.03347535, 0.03915793, 
    0.0537268, 0.01900661, 0.05160894, 0.01185992, 0.001904843, 0.001022762, 
    1.324142e-05, 0.004388743, 3.406525e-05, -1.077839e-05, 0.0477644, 
    0.3096165, 0.1509784, 0.1217639, 0.05335079, 0.03889278, 0.01207789,
  0.2293007, 0.1052435, 0.06809449, 0.08871091, 0.00245337, 0.0263513, 
    0.0424322, 0.06607512, 0.04877469, 0.003110617, 0.004822639, 0.007887457, 
    0.1443444, 0.1695657, 0.1958995, 0.162136, 0.07744265, 0.06391341, 
    0.04514351, 0.09297012, 0.06561383, 0.02747591, 0.1080822, 0.2467207, 
    0.01318991, 0.005191876, 0.00231635, 0.0026464, 0.3219433,
  0.02595188, 0.01435519, 0.02225823, 0.03622876, 0.1052336, 0.01011092, 
    0.02482593, 0.02736438, 0.1128488, 0.2337428, 0.100329, 0.05316103, 
    0.08449603, 0.01607332, -0.0005594598, 0.04985343, 0.05678648, 
    0.07570034, 0.1667874, 0.08007352, 0.03119004, 0.01396681, 0.003070372, 
    0.09257036, 0.1947457, 0.01858834, 0.04846674, 0.04729881, 0.08290562,
  0.0718786, 0.0858587, 0.09750625, 0.1694039, 0.08119843, 0.0985594, 
    0.05441683, 0.01060473, 0.1934581, 0.1757347, 0.1869447, 0.1684714, 
    0.1204468, 0.08624656, 0.05720014, 0.07373464, 0.08188803, 0.06186916, 
    0.02637236, 0.01029389, 0.03946001, 0.05805362, 0.08039556, 0.1043895, 
    0.1355612, 0.1012311, 0.1029111, 0.04011943, 0.04725269,
  0.06423144, 0.06482687, 0.0564161, 0.02153417, 0.1594244, 0.1691542, 
    0.03882658, 0.1270075, 0.1694245, 0.1183759, 0.1353164, 0.1299729, 
    0.2074749, 0.2621417, 0.2294724, 0.2579268, 0.1844822, 0.1389336, 
    0.08029465, 0.02361623, 0.007746023, 0.1452372, 0.1774259, 0.1782701, 
    0.2074206, 0.1550535, 0.1169418, 0.09840946, 0.08483451,
  0.03458212, 0.007271616, 0.04457606, 0.02758012, 0.02099676, 0.09735231, 
    0.09104921, 0.008082526, 0.0005151524, 0.006960676, 0.04362785, 
    0.03417217, 0.04902659, 0.03153661, 0.05045635, 0.07897302, 0.1173358, 
    0.1137467, 0.09116028, -0.0001015841, 0.03217443, 0.07424398, 
    0.006292622, 0.001942432, 0.02092673, 0.05902158, 0.06536317, 0.07625188, 
    0.0607361,
  0.02692898, 0.005500237, 0.01384275, 0.02288892, 0.03047939, 0.01066556, 
    0.0008890733, 0.002845628, 0.0003121658, 0.002833686, 0.012526, 
    0.01890895, 0.03037737, 0.006195644, -1.361469e-09, 0.009982717, 
    0.004979268, 0.01136293, -7.219712e-11, 6.92286e-05, -0.0005674818, 
    0.01580945, 0.004642976, 0.008328716, 0.0003327129, 0.01966047, 
    0.01094081, 0.005780457, 0.03958714,
  0, -1.480145e-08, 0, 0.003382555, 0, 0, 0, 0, 0, 0, 0.009416554, 
    0.01200401, 0.03538601, 0.02697592, 0.02275941, 0.0002224264, 
    0.001082067, -2.895001e-08, -3.263198e-05, 0, 1.673306e-06, 2.917567e-05, 
    0.0006292635, 0.00131116, -3.411209e-06, 0, 0, 0.001050232, -0.0004647899,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.437761e-08, 
    -1.440762e-06, -2.272353e-08, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0001182145, 
    0.0006346832, 0, 0, 0, 0.0001677235, -8.094923e-05, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0003497714, 0, 0, -5.192052e-05, 
    -0.0001378832, 0.0006576773, -9.321905e-05, 0, 0, 0, -0.0002171736, 
    0.0167049, 0.003681475, -6.905026e-05, 0.00151692, 0.001844357, 0, 0, 0, 0,
  0.02449065, 0.04338085, 0.03814333, 0.07334083, 0.0582676, 0.0420657, 
    0.0281286, 0.008636983, 9.370313e-05, 0.003293579, 0.005307619, 
    0.008351292, 0.01744148, 0.03970196, 0.03557269, 0.0240919, 0.014855, 
    0.01533828, 0.005136178, 0.007112693, 0.04182806, 0.0120454, 0.04116476, 
    0.02332578, 0.0105152, 0.01745461, 0.02616729, 0.0078705, 0.01238337,
  0.1631443, 0.1945999, 0.1647147, 0.1139611, 0.1126279, 0.1602094, 
    0.1350179, 0.1142024, 0.1092982, 0.1019034, 0.06392392, 0.1499375, 
    0.06953673, 0.08168712, 0.07477511, 0.0285348, 0.08885469, 0.1167126, 
    0.06990219, 0.07218952, 0.1261403, 0.1201662, 0.2206161, 0.1298621, 
    0.1438514, 0.1182964, 0.1123904, 0.08283069, 0.1123922,
  0.1684072, 0.1568318, 0.1512562, 0.1759789, 0.1764877, 0.07849163, 
    0.08741665, 0.08203059, 0.1172416, 0.1307267, 0.1618665, 0.1716693, 
    0.1240911, 0.07235716, 0.06065647, 0.1204132, 0.09963029, 0.1131328, 
    0.1762569, 0.2849548, 0.187574, 0.1176845, 0.1183374, 0.1118959, 
    0.1157375, 0.09624063, 0.1275467, 0.1637211, 0.2020296,
  0.02356099, 0.0245796, 0.0239036, 0.05990236, 0.1093845, 0.08143609, 
    0.0671754, 0.04657975, 0.1947767, 0.1160652, 0.1145376, 0.06225299, 
    0.04436525, 0.06259183, 0.1555596, 0.1123694, 0.09005262, 0.1302652, 
    0.2099451, 0.1403733, 0.09114963, 0.07120505, 0.02308112, 0.0391307, 
    0.01955388, 0.07943703, 0.06181591, 0.05777856, 0.02469075,
  1.350593e-05, 1.444742e-06, 0.0002106343, 0.1012079, 0.1222754, 0.02919295, 
    0.02344903, 0.05126456, 0.07488193, 0.05851513, 0.01847758, 0.004368467, 
    0.01695042, 0.0900278, 0.1035655, 0.01708935, 0.03877369, 0.03210065, 
    0.03021266, 0.01581188, 2.521252e-05, 2.318024e-06, 1.690809e-07, 
    8.204503e-05, 0.002416693, 0.001451162, 0.0004969093, 0.001779076, 
    0.000102787,
  1.83269e-05, 0.01037416, 0.0009883135, 0.04039055, 0.08307324, 0.0157187, 
    0.04936443, 0.02114321, 0.1070654, 0.05729404, 0.02194047, 0.02176451, 
    0.1503056, 0.07179505, 0.07295079, 0.05859815, 0.03959321, 0.04150494, 
    0.05964593, -0.0002424827, -4.40967e-09, 2.27075e-06, 0.0007396815, 
    0.02789829, 0.0424678, 0.0003739269, 0.00307681, 2.13323e-06, 3.731139e-06,
  0.06718554, 0.3314025, 0.1601875, 0.003517116, 0.00403795, 0.01269321, 
    0.04125947, 0.01843603, 0.1518521, 0.2173367, 0.02236959, 0.03838145, 
    0.0382179, 0.01971583, 0.03611244, 0.01290304, 0.002007611, 0.0002078721, 
    -1.095125e-06, 0.006073423, -0.0001172428, 2.597349e-06, 0.02743062, 
    0.2802593, 0.1484225, 0.1415097, 0.05976427, 0.02909147, 0.01486734,
  0.2244712, 0.0644239, 0.04989837, 0.06168878, 0.001868075, 0.0196871, 
    0.0336963, 0.04231128, 0.02757825, 0.003532092, 0.004002934, 0.006786677, 
    0.1185971, 0.1808717, 0.2003857, 0.1569382, 0.06551082, 0.0659751, 
    0.06258289, 0.07255991, 0.04175128, 0.02780622, 0.08314273, 0.1831231, 
    0.01371629, 0.002638008, 0.00130386, 0.005165956, 0.2557782,
  0.02929084, 0.01078255, 0.03196349, 0.02208834, 0.07207334, 4.844116e-05, 
    0.027345, 0.02366082, 0.07249846, 0.2348132, 0.08557262, 0.03887006, 
    0.08135894, 0.005700632, 0.001069744, 0.03134984, 0.03231407, 0.03223914, 
    0.1522273, 0.04837652, 0.03309973, 0.01425952, 0.00243777, 0.07104763, 
    0.1579643, 0.01414623, 0.05762366, 0.02175756, 0.06357771,
  0.06397015, 0.07906745, 0.09022073, 0.1428792, 0.0560181, 0.0686996, 
    0.04387002, 0.02036977, 0.3078146, 0.1297825, 0.1498505, 0.1891789, 
    0.121885, 0.05174895, 0.04590241, 0.06551843, 0.04958907, 0.04562331, 
    0.0187815, 0.007163337, 0.03401245, 0.06178284, 0.07279958, 0.09271346, 
    0.1254388, 0.07593745, 0.07509647, 0.03030507, 0.04613945,
  0.1040768, 0.09054518, 0.1056382, 0.05436474, 0.1400485, 0.1521482, 
    0.0903863, 0.126085, 0.1640393, 0.1516235, 0.1585823, 0.1454504, 
    0.1986108, 0.2577172, 0.2429984, 0.2360712, 0.1873559, 0.1498461, 
    0.07880798, 0.09457577, 0.02828912, 0.1598017, 0.168992, 0.2100498, 
    0.2060869, 0.1582038, 0.09252806, 0.08050209, 0.08277693,
  0.1656109, 0.0564889, 0.1264373, 0.1076738, 0.07892597, 0.1173099, 
    0.1554633, 0.03640373, 0.02039797, 0.0664655, 0.1111281, 0.06549942, 
    0.1486963, 0.08683352, 0.09052897, 0.1144847, 0.1938656, 0.1687794, 
    0.1501905, 0.02873053, 0.1546772, 0.1409012, 0.01605078, 0.0264667, 
    0.07047923, 0.1124826, 0.1000566, 0.1647374, 0.1564491,
  0.1706931, 0.09637321, 0.1280212, 0.04807913, 0.03269547, 0.02093716, 
    0.006290999, 0.02481141, 0.01304909, 0.007769153, 0.0336856, 0.0248668, 
    0.04529891, 0.03194864, 0.0004795214, 0.01474157, 0.0180201, 0.05542217, 
    0.00545834, 0.05794075, 0.04062178, 0.0297203, 0.02064634, 0.02350572, 
    0.01372721, 0.09019045, 0.04984321, 0.09251413, 0.1361689,
  0.0372131, 0.02767716, 4.768549e-05, 0.0126264, 0.006970289, 0, 0, 
    -4.087559e-07, 0, -9.113275e-05, 0.02325665, 0.02061969, 0.02853911, 
    0.02453097, 0.02168588, 0.006554455, 0.0113478, 0.04204722, 0.05012693, 
    0.08683282, 0.03796531, 0.01621107, 0.0230933, 0.02588404, 0.01548557, 
    -1.237446e-05, -1.811295e-06, 0.01462199, 0.03997575,
  -1.98839e-05, 0, 0, 0, -1.794999e-10, 3.188138e-10, 0, 0, 0, 0, 0, 
    0.0002509782, 0.00798863, 0.01296248, 0.02016297, 0.02121039, 0.01590701, 
    0.001199434, -2.857617e-08, 6.839722e-06, 2.246331e-06, -2.497999e-05, 
    -5.894575e-07, 0, -4.250295e-07, 0, 0, -0.0001703923, 9.015411e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0002775179, 
    0.006437604, -9.23616e-05, -1.897936e-05, 0, 0.002401208, 0.003422722, 
    -5.07258e-05, 0, 0, 0, 0,
  0, 0.0002584468, -9.165994e-06, 0.00016791, 0, 0, 0, 0, 0, 0.001370391, 0, 
    0, 0.0003138207, 0.00577522, 0.001180842, 0.00235383, -7.856131e-05, 
    -8.989078e-05, -5.029991e-05, 0.01008169, 0.06335805, 0.04837646, 
    0.007359813, 0.002601441, 0.006308641, -0.0001625308, 0.001985594, 
    1.857746e-05, 6.775482e-05,
  0.05769893, 0.0810067, 0.1019855, 0.1634279, 0.1567877, 0.1327486, 
    0.08450617, 0.05586649, 0.04361417, 0.03881603, 0.05564607, 0.09712002, 
    0.2047881, 0.1781292, 0.1218077, 0.1013451, 0.07565433, 0.03778183, 
    0.03424137, 0.1083241, 0.08071841, 0.06511086, 0.1067761, 0.09070963, 
    0.08285838, 0.05718762, 0.06689002, 0.07189195, 0.04388232,
  0.2179336, 0.2538643, 0.2156243, 0.1943167, 0.1475358, 0.2070043, 
    0.1579586, 0.1742801, 0.1492652, 0.1740874, 0.1659853, 0.2177865, 
    0.1698946, 0.1276294, 0.1229653, 0.1100332, 0.1436916, 0.1353022, 
    0.1199505, 0.1130049, 0.1444516, 0.1523857, 0.2564803, 0.1923805, 
    0.1908006, 0.2216108, 0.1817169, 0.1548037, 0.1799182,
  0.1728194, 0.1316076, 0.1551652, 0.1493451, 0.1473244, 0.06532517, 
    0.08904167, 0.08679925, 0.1132974, 0.1123549, 0.1560346, 0.1818316, 
    0.1641249, 0.08236822, 0.08455728, 0.1887956, 0.1207832, 0.1071723, 
    0.1721776, 0.252606, 0.1829577, 0.1220313, 0.1372435, 0.1316904, 
    0.09712587, 0.08002301, 0.1205703, 0.160002, 0.2029731,
  0.01503179, 0.009861374, 0.01457121, 0.04006801, 0.08691742, 0.06052288, 
    0.06402185, 0.02596462, 0.1686027, 0.09646817, 0.0898385, 0.05199236, 
    0.04035505, 0.04808126, 0.1080278, 0.1025773, 0.08892395, 0.1106145, 
    0.2008307, 0.1161955, 0.1017866, 0.08500122, 0.0220783, 0.05528346, 
    0.01675518, 0.06771783, 0.05022496, 0.04997164, 0.02488958,
  4.439465e-06, 8.949585e-07, 0.0001517622, 0.06962112, 0.09564848, 
    0.02378882, 0.01648085, 0.03777822, 0.08315133, 0.07076858, 0.008293374, 
    0.003632973, 0.02398946, 0.09684399, 0.1019561, 0.009737272, 0.03717651, 
    0.03167334, 0.02284188, 0.02038009, 1.904224e-06, 7.875926e-07, 
    1.270886e-08, 0.0001890652, 0.001940227, 0.0004373341, 9.860082e-05, 
    0.0007621545, 6.331627e-06,
  2.032854e-05, 0.002699015, 0.002321599, 0.0604829, 0.08036449, 0.0121427, 
    0.04872355, 0.01457231, 0.09896854, 0.03777769, 0.01553893, 0.02765932, 
    0.1500472, 0.04774263, 0.05594962, 0.03584033, 0.03946857, 0.03942413, 
    0.05758494, -0.0001038749, 1.315738e-08, 7.53394e-07, -6.678547e-05, 
    0.02357007, 0.02711304, 0.001201046, 0.002522187, 5.266571e-05, 
    1.63124e-06,
  0.04645478, 0.2762443, 0.1440375, 0.007473727, 0.004096085, 0.006277502, 
    0.02430931, 0.01712444, 0.1137699, 0.163928, 0.01784898, 0.03382936, 
    0.0233777, 0.01420272, 0.02436233, 0.01024077, 0.002364151, 0.00043435, 
    0.0002218135, 0.0117404, 2.270746e-05, 0.001323778, 0.02226766, 
    0.2353921, 0.1414367, 0.1536891, 0.06475889, 0.02916128, 0.01450923,
  0.1455694, 0.03494254, 0.03888163, 0.05272538, 0.003573617, 0.01371668, 
    0.0259941, 0.02171666, 0.01192712, 0.002793207, 0.003256738, 0.006511641, 
    0.09101064, 0.182464, 0.2135375, 0.1187838, 0.06389419, 0.06159401, 
    0.08793975, 0.05745851, 0.02472382, 0.02664149, 0.071416, 0.1309131, 
    0.01624086, 0.002304019, 0.0009254331, 0.00378621, 0.1995604,
  0.02028712, 0.005787453, 0.03160535, 0.01060466, 0.04725897, 9.663107e-06, 
    0.03123696, 0.0282694, 0.04876374, 0.2428224, 0.05906092, 0.03342921, 
    0.07716695, 0.002528015, 0.0007952247, 0.02381159, 0.01005336, 
    0.03844176, 0.09973998, 0.01762523, 0.02221072, 0.01487469, 0.002691531, 
    0.06526649, 0.1229872, 0.02129134, 0.02059316, 0.004020887, 0.06337494,
  0.05533438, 0.06174839, 0.08452877, 0.1143181, 0.04020434, 0.05649887, 
    0.04421506, 0.05622907, 0.3516096, 0.1063999, 0.1244285, 0.1995987, 
    0.135421, 0.04503162, 0.04249937, 0.04372106, 0.02987474, 0.02534239, 
    0.01730227, 0.003628128, 0.02797172, 0.05344927, 0.06866196, 0.07477055, 
    0.09538136, 0.06248533, 0.05206138, 0.01998324, 0.03982656,
  0.08879691, 0.07632133, 0.1052047, 0.1165518, 0.1328614, 0.1362565, 
    0.1374435, 0.09684824, 0.146934, 0.1431639, 0.1620357, 0.1220348, 
    0.1889527, 0.2516507, 0.2462101, 0.2287028, 0.1462932, 0.1353735, 
    0.07162411, 0.1332621, 0.09631862, 0.1430683, 0.1459177, 0.2028052, 
    0.2058342, 0.1608122, 0.0813236, 0.06828732, 0.07158393,
  0.1739822, 0.1046327, 0.1321468, 0.1373583, 0.09330744, 0.1191394, 
    0.1455671, 0.09773873, 0.06681056, 0.1551829, 0.2060583, 0.1536582, 
    0.1901783, 0.1091897, 0.109172, 0.1402897, 0.2203992, 0.2010406, 
    0.1860473, 0.1043174, 0.2423217, 0.1259815, 0.02123054, 0.05680733, 
    0.1288585, 0.1322767, 0.1368492, 0.1684186, 0.1729859,
  0.2759547, 0.1883366, 0.1865567, 0.1427213, 0.0978311, 0.07585417, 
    0.1054075, 0.07705104, 0.06028059, 0.07677013, 0.09840251, 0.0660143, 
    0.08623687, 0.05577976, 0.04154307, 0.0765698, 0.0445487, 0.1168799, 
    0.06905372, 0.09065569, 0.06409835, 0.09220652, 0.0251814, 0.07289227, 
    0.1424905, 0.1715424, 0.1446052, 0.2019261, 0.1789888,
  0.1846614, 0.1405677, 0.07152187, 0.03944952, 0.006093662, 0, 
    -8.816487e-07, 0.0009603439, 0.01586927, 0.0280086, 0.03305823, 
    0.0271839, 0.04655863, 0.07290822, 0.04795872, 0.03199246, 0.1044575, 
    0.1078657, 0.1389307, 0.1467588, 0.06843682, 0.09386484, 0.06687573, 
    0.02477966, 0.02804852, -0.0001398527, 3.887996e-05, 0.1378482, 0.2239634,
  -0.0003678371, 7.832998e-05, 0.002291162, 0.0007449272, -0.0002081106, 
    0.001540557, 0.02442846, 0.03503199, 0.03083915, 0.02116645, 0.02035471, 
    0.01648151, 0.03756419, 0.03965763, 0.04894991, 0.05834197, 0.08066525, 
    0.1121351, 0.0823435, 0.08695683, 0.09728623, 0.07501165, 0.01336873, 
    -0.001606027, 0.001508606, 1.272564e-05, 0, -0.0002514055, 0.001155233,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0009713783, 
    0.008742504, -7.234743e-05, -0.0003008647, -0.0001365967, 0.004074199, 
    0.04957789, 0.03114064, -0.0008042764, -6.987351e-08, 0, 0,
  0.006936261, 0.02774658, 0.03023747, 0.008201281, -8.63297e-05, 0, 
    -0.0001243174, 0, -0.0001150729, 0.002435428, -4.163269e-05, 
    -0.0002601424, 0.002570459, 0.03823582, 0.05369695, 0.05800037, 
    0.02573021, 0.003998356, 0.01271995, 0.05936287, 0.1497885, 0.1841859, 
    0.1436684, 0.06749772, 0.06311619, 0.02198954, 0.03165125, 0.01142867, 
    0.005991456,
  0.09640791, 0.1562241, 0.1622608, 0.1849505, 0.1949056, 0.1806976, 
    0.114613, 0.1304348, 0.141698, 0.1114738, 0.1587396, 0.25987, 0.2916202, 
    0.2280549, 0.1780914, 0.1778296, 0.1755138, 0.1544993, 0.1283183, 
    0.1965025, 0.1553558, 0.1414368, 0.157977, 0.1885183, 0.2179898, 
    0.180267, 0.1260184, 0.1223985, 0.05628711,
  0.2492351, 0.2814319, 0.2264195, 0.2000599, 0.1638561, 0.1857896, 
    0.1679671, 0.1845431, 0.1673583, 0.1704114, 0.1844632, 0.2618061, 
    0.1713385, 0.1546418, 0.1204786, 0.1065788, 0.1530462, 0.1389975, 
    0.1391819, 0.1530496, 0.1742241, 0.215261, 0.2833418, 0.2645878, 
    0.2191076, 0.2257638, 0.1999983, 0.1894716, 0.2243262,
  0.1664733, 0.1190591, 0.1295611, 0.1215535, 0.1261677, 0.06352081, 
    0.07409472, 0.09037098, 0.08472072, 0.1049614, 0.1374408, 0.1700186, 
    0.1582976, 0.07819468, 0.1013244, 0.212847, 0.1128722, 0.09685659, 
    0.1575936, 0.2261107, 0.1823894, 0.1299692, 0.1374512, 0.1238215, 
    0.0743609, 0.08004908, 0.1156076, 0.1536891, 0.1986784,
  0.008890727, 0.0003054241, 0.0050348, 0.02340187, 0.0740257, 0.04864126, 
    0.05488301, 0.01657185, 0.1529132, 0.07592877, 0.05964082, 0.05167153, 
    0.04513768, 0.03827893, 0.07834886, 0.1015774, 0.0938173, 0.1100068, 
    0.1901432, 0.08335344, 0.08180671, 0.0710975, 0.02043964, 0.07040903, 
    0.01668569, 0.05509604, 0.04954457, 0.05564791, 0.0258493,
  9.326003e-07, 2.274433e-07, 0.000351851, 0.04626751, 0.07968993, 
    0.02065937, 0.002917633, 0.01984835, 0.07952872, 0.05306228, 0.004280929, 
    0.00737708, 0.02875865, 0.09960736, 0.1020036, 0.009369698, 0.03935354, 
    0.02601384, 0.01537485, 0.01187393, -7.744911e-08, 5.216567e-07, 
    6.035393e-08, 0.0003943652, 0.002019949, 2.80788e-05, 0.0001251618, 
    2.144347e-05, 1.107979e-06,
  1.39723e-05, 0.002081973, 0.008110165, 0.07991891, 0.08976253, 0.009189713, 
    0.04715509, 0.01126567, 0.09917779, 0.03201757, 0.01401243, 0.01414322, 
    0.1593076, 0.03850186, 0.04678087, 0.0212086, 0.03982821, 0.03698449, 
    0.05905869, 0.008127553, -6.553221e-07, 3.789929e-07, 0.002085819, 
    0.0252564, 0.01073719, 0.0004914249, 0.007898345, 0.002135564, 5.6332e-07,
  0.03529455, 0.2208937, 0.1373054, 0.01234211, 0.004602502, 0.00529848, 
    0.01300355, 0.01318732, 0.08582336, 0.1491975, 0.01842315, 0.03130048, 
    0.01446557, 0.01138365, 0.0161508, 0.008785388, 0.0028931, 0.0005337805, 
    0.0006623078, 0.01327365, 0.000368659, 0.001301226, 0.02377862, 
    0.2128934, 0.1281642, 0.1733066, 0.07140268, 0.03776937, 0.02297194,
  0.09031221, 0.02493709, 0.03731402, 0.03565756, 0.003415237, 0.01002827, 
    0.01774339, 0.01162089, 0.005947301, 0.002613035, 0.003998759, 
    0.006441291, 0.08566539, 0.1781483, 0.2132782, 0.0992021, 0.06567054, 
    0.04292584, 0.08871962, 0.04200203, 0.01741885, 0.02484496, 0.05720731, 
    0.1022624, 0.02194613, 0.001097946, 0.0006272395, 0.002354929, 0.1529884,
  0.006871779, 0.01029829, 0.03392737, 0.006172976, 0.01907537, 7.737147e-06, 
    0.01798525, 0.03113719, 0.03990362, 0.2483868, 0.03715495, 0.0280279, 
    0.07786272, 0.0001102726, 0.0006857335, 0.02035227, 0.002037658, 
    0.02997834, 0.05383189, 0.000698221, 0.01230024, 0.01866762, 0.002517489, 
    0.05564705, 0.08489103, 0.01760257, 0.009276404, 0.0004648275, 0.04827477,
  0.0349888, 0.05208889, 0.08758441, 0.1013389, 0.03687493, 0.04801065, 
    0.04310874, 0.08434684, 0.3325291, 0.08520489, 0.1081968, 0.1791763, 
    0.1228586, 0.01906579, 0.01918806, 0.02269964, 0.01436996, 0.01319289, 
    0.012224, -1.698435e-05, 0.02381847, 0.04216769, 0.05481676, 0.06576236, 
    0.08835726, 0.02562173, 0.02733542, 0.002297443, 0.02778787,
  0.06658498, 0.05861123, 0.09841014, 0.1113163, 0.1186366, 0.1234722, 
    0.1397861, 0.08305676, 0.1269008, 0.1147816, 0.1580439, 0.1021731, 
    0.1801859, 0.2305343, 0.2235314, 0.2227288, 0.1307507, 0.1239624, 
    0.06753215, 0.1204231, 0.160761, 0.1445006, 0.1173056, 0.1875401, 
    0.199551, 0.1694843, 0.08159695, 0.07377526, 0.04863781,
  0.1341167, 0.1034378, 0.1154724, 0.1125012, 0.08353215, 0.1090785, 
    0.1600977, 0.1364436, 0.1579466, 0.1706168, 0.2527997, 0.1897651, 
    0.1978073, 0.1287498, 0.1102357, 0.1525827, 0.2220847, 0.1843963, 
    0.1592417, 0.1091373, 0.2208043, 0.1163356, 0.05253356, 0.1063415, 
    0.1723885, 0.1453481, 0.162198, 0.1531334, 0.1520882,
  0.2185496, 0.1689212, 0.1661312, 0.1533939, 0.125993, 0.1256955, 0.1671994, 
    0.1645212, 0.1459582, 0.1673303, 0.1232444, 0.09213759, 0.104648, 
    0.1550124, 0.1237233, 0.1053323, 0.1168555, 0.1927, 0.1794576, 0.1616909, 
    0.07842315, 0.0858966, 0.05347904, 0.1455413, 0.2208728, 0.2262222, 
    0.1437448, 0.2052003, 0.1717729,
  0.25475, 0.178461, 0.1101192, 0.09001095, 0.04147343, 0.0238414, 
    0.04350593, 0.08250347, 0.0742118, 0.1045879, 0.1060459, 0.09627917, 
    0.08585234, 0.09674014, 0.1076354, 0.1344955, 0.1767006, 0.1947986, 
    0.1433, 0.1314526, 0.0684799, 0.07852077, 0.07741866, 0.03742087, 
    0.0599185, 0.0006505795, -0.0001175811, 0.287863, 0.2723178,
  0.07314336, 0.09981824, 0.08579124, 0.0694987, 0.06427545, 0.06811557, 
    0.08350024, 0.1171948, 0.07905539, 0.07203677, 0.06714471, 0.1210737, 
    0.1983512, 0.216076, 0.2199881, 0.2114599, 0.1903253, 0.1647449, 
    0.1338344, 0.1079406, 0.1009029, 0.09796257, 0.04768187, 0.0247422, 
    0.006563324, 0.000275396, -0.001847196, 0.008759896, 0.08302807,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002368521, 0.0003683763, 
    0.004091725, 0.003255693, 0.01637995, 0.0001818558, -0.0007000362, 
    -0.0006771439, 0.02865341, 0.1163156, 0.07059322, 0.004841869, 
    0.001924089, -0.0006619827, 0,
  0.1146769, 0.1179924, 0.1288479, 0.05992271, -0.0009962739, -2.51956e-05, 
    0.0294563, -7.651523e-05, -0.0003326167, 0.002005254, 0.003329374, 
    0.006324784, 0.03107954, 0.1120923, 0.1312456, 0.1125926, 0.06125804, 
    0.04584854, 0.02755217, 0.09242181, 0.3194093, 0.2697802, 0.2557583, 
    0.1592828, 0.1309635, 0.1034087, 0.0901645, 0.07388386, 0.1193921,
  0.1052002, 0.1586328, 0.2119767, 0.2074196, 0.2194118, 0.2014793, 
    0.1704975, 0.154959, 0.1878291, 0.1584978, 0.2208889, 0.2698736, 
    0.2877123, 0.2517393, 0.1985563, 0.1979648, 0.1900735, 0.1874609, 
    0.1772682, 0.2546605, 0.2393472, 0.2109933, 0.2436813, 0.2342582, 
    0.2954712, 0.2708577, 0.1860958, 0.1329647, 0.1302437,
  0.239361, 0.2783909, 0.1915486, 0.1880818, 0.1502723, 0.1882109, 0.1701751, 
    0.1632871, 0.1568276, 0.166751, 0.2125499, 0.2476351, 0.1497417, 
    0.1382779, 0.1141599, 0.1012323, 0.1630889, 0.1474351, 0.1231998, 
    0.1473074, 0.186537, 0.2281584, 0.2471614, 0.2810296, 0.2176507, 
    0.2166957, 0.1954739, 0.2171583, 0.2142415,
  0.1526093, 0.1096262, 0.1150042, 0.09055049, 0.1153537, 0.05655604, 
    0.08559258, 0.06767871, 0.06462123, 0.08616693, 0.1147347, 0.1428691, 
    0.1393692, 0.07484014, 0.1063166, 0.1997748, 0.09536576, 0.09179463, 
    0.1583, 0.1906053, 0.1690388, 0.1195349, 0.1254737, 0.1187502, 
    0.06058659, 0.07186446, 0.100834, 0.1404945, 0.1796206,
  0.01227663, 0.003612823, 0.009289641, 0.01837034, 0.07252665, 0.05220162, 
    0.03782586, 0.01003164, 0.1146431, 0.05686094, 0.04861816, 0.04947321, 
    0.04599943, 0.03370734, 0.06630409, 0.109619, 0.1120535, 0.09870037, 
    0.1696959, 0.06111356, 0.06514155, 0.05819181, 0.02382424, 0.09488887, 
    0.01980808, 0.05317355, 0.04739364, 0.0609924, 0.03648676,
  1.973376e-07, 4.601736e-08, 0.000408812, 0.02625207, 0.06982762, 0.015842, 
    -0.0004394812, 0.02087614, 0.07083122, 0.0320025, 0.0004817093, 
    0.0007879431, 0.03223133, 0.09119781, 0.0812935, 0.001945749, 0.04461723, 
    0.01846316, 0.01269908, 0.002054583, 2.526408e-07, 1.33276e-07, 
    1.697575e-08, 0.0005594415, 0.002074387, 0.0001301706, 0.000483351, 
    -9.501537e-06, 4.577588e-07,
  8.634504e-06, 0.02017804, 0.003985283, 0.08922853, 0.09334704, 0.009488049, 
    0.04691847, 0.009988637, 0.09751213, 0.03871124, 0.004591984, 
    0.008124046, 0.1634597, 0.03232611, 0.03821959, 0.01762403, 0.03880928, 
    0.03811083, 0.06206475, 0.01911756, -0.0001732092, 1.929033e-06, 
    0.000259929, 0.02384947, 0.006298033, 0.0004080077, 0.008158539, 
    0.0005356006, 1.216372e-07,
  0.02790921, 0.1994119, 0.146406, 0.009015718, 0.004660015, 0.007820104, 
    0.01411562, 0.01103558, 0.07469491, 0.1262456, 0.01806622, 0.02525447, 
    0.01139134, 0.008853004, 0.01283843, 0.009041618, 0.004070027, 
    0.005860223, 0.001951348, 0.007231069, 3.329053e-05, 0.00494017, 
    0.03511447, 0.1970614, 0.1278091, 0.1862568, 0.08574913, 0.03460125, 
    0.03132419,
  0.04928784, 0.02570052, 0.05234919, 0.03116341, 0.003360668, 0.007262857, 
    0.01147946, 0.007407327, 0.00406035, 0.002997523, 0.006834712, 
    0.005582196, 0.07282429, 0.1520788, 0.2169743, 0.09835389, 0.07746828, 
    0.02842775, 0.1053536, 0.03481397, 0.01292779, 0.02529197, 0.04214389, 
    0.08937044, 0.02389915, 0.001410945, 0.0004624623, 0.01295691, 0.111176,
  0.002384933, 0.02902271, 0.03316175, 0.01109943, 0.003401082, 3.295675e-06, 
    0.004183853, 0.03231014, 0.04154279, 0.2312775, 0.01966261, 0.02674366, 
    0.0728144, 0.0001009105, 0.009095006, 0.01915222, 0.000637325, 
    0.006102141, 0.02767914, 0.0004253289, 0.01707485, 0.02536384, 
    0.00185074, 0.04938313, 0.0589727, 0.01618004, 0.0009447345, 0.007181202, 
    0.03228986,
  0.03149231, 0.05983416, 0.08329175, 0.08855678, 0.03744523, 0.04292559, 
    0.07661565, 0.1330006, 0.3228662, 0.07236954, 0.09803382, 0.1743003, 
    0.1173797, 0.01806504, 0.01241543, 0.006431073, 0.008493715, 0.01072665, 
    0.009134026, 7.476179e-06, 0.01508881, 0.0378034, 0.05574828, 0.05934104, 
    0.08325717, 0.02907223, 0.008242167, 0.0001379605, 0.0161659,
  0.05957512, 0.04271664, 0.09540402, 0.09323129, 0.1049961, 0.111356, 
    0.1477379, 0.0787256, 0.1174492, 0.09372049, 0.1554696, 0.08537181, 
    0.1574242, 0.220266, 0.1976309, 0.2180733, 0.1275321, 0.1130378, 
    0.05644529, 0.1255574, 0.1534667, 0.1498221, 0.09618147, 0.1880044, 
    0.1956974, 0.1571823, 0.05897992, 0.06812239, 0.04545973,
  0.1072064, 0.09445885, 0.1089169, 0.1006364, 0.07875165, 0.1093044, 
    0.1522908, 0.1557989, 0.1844409, 0.166286, 0.2765903, 0.2059996, 
    0.1961457, 0.1167029, 0.09872475, 0.1667937, 0.2239992, 0.1647144, 
    0.138815, 0.09812337, 0.1916392, 0.1173368, 0.06836429, 0.1257068, 
    0.1793698, 0.1363117, 0.1550474, 0.1429107, 0.1434954,
  0.1805879, 0.1437845, 0.1406675, 0.1620838, 0.13952, 0.1578415, 0.2271371, 
    0.2193735, 0.193424, 0.2276039, 0.1985878, 0.1288293, 0.1333618, 
    0.1879213, 0.135975, 0.1418668, 0.1555325, 0.2560275, 0.1756756, 
    0.1440349, 0.07759208, 0.07536105, 0.05014864, 0.2057371, 0.2135628, 
    0.2299568, 0.1216995, 0.178583, 0.1378643,
  0.2269312, 0.1558769, 0.1211276, 0.1179327, 0.08236526, 0.2016703, 
    0.1058729, 0.1907137, 0.1424943, 0.1906702, 0.1304814, 0.1532554, 
    0.1470502, 0.1535468, 0.1246537, 0.1431068, 0.1702751, 0.1770205, 
    0.1432357, 0.1089597, 0.06721056, 0.06041093, 0.08356441, 0.06126341, 
    0.08748955, 0.01684792, -0.001403711, 0.2500425, 0.225325,
  0.1008848, 0.1479491, 0.1641841, 0.1976067, 0.1971233, 0.1986454, 
    0.1065635, 0.1421417, 0.1026742, 0.08953957, 0.07493819, 0.1728337, 
    0.2493241, 0.2079485, 0.2200085, 0.217324, 0.183585, 0.1670466, 
    0.1276423, 0.1005484, 0.08328689, 0.0858269, 0.06862419, 0.06354795, 
    0.02607802, 0.00404356, -0.005235537, 0.06055393, 0.09868871,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.713419e-05, -1.713419e-05, 
    -1.713419e-05, -1.713419e-05, -1.713419e-05, -1.713419e-05, 
    -1.713419e-05, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.704719e-05, 0.01835143, 0.04374435, 
    0.09455585, 0.09837599, 0.03931641, 0.03981231, 0.00524681, 0.002722418, 
    -0.001740858, 0.1030576, 0.2302865, 0.1732069, 0.04708578, 0.01229202, 
    0.0003242886, 0,
  0.1782957, 0.2405498, 0.2037584, 0.1225946, -0.002516051, -0.001176387, 
    0.06984939, -0.0004106409, 0.0001942032, 0.007147259, 0.008995079, 
    0.009432752, 0.09197792, 0.1637071, 0.1582555, 0.1407306, 0.09132707, 
    0.09490141, 0.1144502, 0.2285594, 0.4617833, 0.3421134, 0.312672, 
    0.24157, 0.2653107, 0.1616722, 0.1273697, 0.1704415, 0.1951085,
  0.1395097, 0.1560363, 0.2456988, 0.209529, 0.235936, 0.2168956, 0.2078012, 
    0.1936994, 0.192454, 0.2288986, 0.3101062, 0.3120443, 0.3278793, 
    0.2529153, 0.2015996, 0.2097407, 0.2085708, 0.2201907, 0.2391746, 
    0.2995371, 0.2955612, 0.2705014, 0.2638955, 0.2638615, 0.2901231, 
    0.3062075, 0.2062513, 0.1285715, 0.1585253,
  0.253758, 0.2907147, 0.2011458, 0.1928063, 0.1433538, 0.1893171, 0.1737254, 
    0.1435586, 0.172609, 0.1785897, 0.2184153, 0.2347135, 0.1472859, 
    0.1209495, 0.1039874, 0.07829489, 0.1618343, 0.1480183, 0.1349871, 
    0.1483338, 0.1838164, 0.2303997, 0.2466068, 0.2648362, 0.2254478, 
    0.2196146, 0.1810738, 0.2345189, 0.2183906,
  0.1433868, 0.0926298, 0.1004421, 0.082849, 0.1024786, 0.04985543, 
    0.08498564, 0.06976458, 0.05801418, 0.0768717, 0.1020932, 0.128414, 
    0.1323166, 0.06955511, 0.09473774, 0.185799, 0.08827902, 0.08360511, 
    0.148908, 0.2005974, 0.1486921, 0.1093233, 0.119205, 0.120074, 
    0.04567944, 0.07996639, 0.08060689, 0.1363057, 0.2077924,
  0.008275694, 0.004432788, 0.01142226, 0.02281531, 0.07197494, 0.04494044, 
    0.02549599, 0.005945705, 0.09829645, 0.04166124, 0.03450931, 0.04690698, 
    0.04354855, 0.02953578, 0.06168658, 0.1154667, 0.1517237, 0.08748793, 
    0.1468567, 0.05434811, 0.05538215, 0.04625705, 0.01269778, 0.1036562, 
    0.01833957, 0.04446661, 0.03757701, 0.05245702, 0.03003944,
  7.57154e-08, 1.237648e-08, 0.0003529408, 0.0146728, 0.0525037, 0.02137724, 
    -0.0008111947, 0.0203052, 0.07514715, 0.007593046, 1.378943e-05, 
    1.878889e-05, 0.03420547, 0.0960232, 0.05458251, 0.001707331, 0.05048193, 
    0.01326345, 0.01140693, 0.0008373653, 3.371598e-07, 3.610263e-08, 
    1.217947e-08, 0.0003118917, 0.001569534, 2.277886e-05, 0.0003059067, 
    1.901789e-05, 3.267665e-07,
  2.670168e-06, 0.0262964, 0.00443985, 0.09492535, 0.0880525, 0.01006869, 
    0.05674361, 0.00879748, 0.09204732, 0.04173706, 0.002714806, 0.004685087, 
    0.156855, 0.03594488, 0.03223773, 0.01711682, 0.03484785, 0.04002442, 
    0.06375042, 0.0276012, 0.001867763, 3.978724e-07, 2.734002e-07, 
    0.02273002, 0.00416223, 0.0002015486, 0.006985913, -9.901178e-05, 
    3.883945e-07,
  0.01584998, 0.1900633, 0.1413628, 0.006989155, 0.00443501, 0.010194, 
    0.009281172, 0.008486147, 0.07153697, 0.1211764, 0.01442651, 0.02172748, 
    0.009137206, 0.00715528, 0.01235813, 0.01062801, 0.005016468, 
    0.004219847, 0.002514389, 0.007614481, 0.002556437, 0.02601964, 
    0.03665924, 0.1978348, 0.1232734, 0.1856259, 0.1055149, 0.02347082, 
    0.02158172,
  0.04254818, 0.02443863, 0.05296866, 0.02970554, 0.002916576, 0.005993314, 
    0.01088071, 0.00636715, 0.003364662, 0.003043088, 0.007910588, 
    0.005504678, 0.07125383, 0.1445789, 0.2181413, 0.1274382, 0.05732953, 
    0.02147156, 0.109911, 0.06044243, 0.01510697, 0.02416093, 0.04091951, 
    0.07987846, 0.01802885, 0.00172054, 0.0002699408, 0.01534178, 0.09116601,
  0.0008874404, 0.04448713, 0.03146952, 0.01524349, 0.0001570903, 
    1.335816e-06, 0.0008314712, 0.03921252, 0.03634011, 0.2400208, 0.0101504, 
    0.02928801, 0.07346867, 0.0003780043, 0.001459044, 0.01207953, 
    0.0005320763, 0.001559743, 0.01851255, 0.0004277266, 0.001181681, 
    0.03053224, 0.001531897, 0.04755995, 0.03670719, 0.0130974, 2.305871e-05, 
    0.03468356, 0.0180802,
  0.04914802, 0.0632743, 0.06584686, 0.08020793, 0.03597836, 0.03754443, 
    0.05686617, 0.151304, 0.3062634, 0.06367411, 0.08991766, 0.173886, 
    0.113337, 0.01853229, 0.001878314, 0.007690615, 0.01021406, 0.009404712, 
    0.0006656802, 2.181783e-05, 0.009466884, 0.02675653, 0.04939079, 
    0.05330911, 0.07898936, 0.01887586, 0.0008296865, 1.149686e-05, 
    0.006158231,
  0.06322151, 0.03287251, 0.0911274, 0.08444498, 0.09589842, 0.1124092, 
    0.1436547, 0.07653224, 0.110197, 0.09252927, 0.1462667, 0.07847113, 
    0.1373414, 0.2073642, 0.1688987, 0.1927687, 0.1042555, 0.100503, 
    0.0451402, 0.1259938, 0.1487469, 0.1469547, 0.08568059, 0.1845388, 
    0.1845579, 0.1566752, 0.0665318, 0.06733376, 0.03400452,
  0.09285993, 0.1011006, 0.1045853, 0.0972713, 0.08963039, 0.1111684, 
    0.1454357, 0.1620929, 0.186329, 0.1555476, 0.2724701, 0.2068012, 
    0.1910432, 0.09964047, 0.1003396, 0.1704593, 0.2409792, 0.1595518, 
    0.1192364, 0.08793819, 0.1697158, 0.1214275, 0.06871819, 0.1292374, 
    0.177508, 0.1212174, 0.1304064, 0.1530723, 0.136848,
  0.180785, 0.1339123, 0.123201, 0.1652271, 0.1391727, 0.1617569, 0.2774836, 
    0.2514153, 0.1984392, 0.2374573, 0.1887915, 0.1617965, 0.1620066, 
    0.1877244, 0.1499047, 0.1500698, 0.1714393, 0.2824266, 0.1718964, 
    0.1432602, 0.07602269, 0.07676955, 0.04485229, 0.1856601, 0.2023955, 
    0.2460648, 0.1167309, 0.1743413, 0.1298361,
  0.2039615, 0.1530507, 0.1105252, 0.1153909, 0.09070779, 0.2393692, 
    0.1265679, 0.2002815, 0.1686934, 0.203746, 0.144969, 0.1397047, 
    0.1432211, 0.142993, 0.1214454, 0.1514601, 0.1504091, 0.1517923, 
    0.1339211, 0.1010806, 0.07436533, 0.04914792, 0.1028587, 0.07836429, 
    0.08959904, 0.03911794, -3.857312e-05, 0.2301844, 0.2175399,
  0.08704207, 0.1382954, 0.1683529, 0.208499, 0.1940459, 0.2028231, 
    0.08706716, 0.1362023, 0.1266239, 0.07473247, 0.06340312, 0.1286109, 
    0.2311284, 0.2013573, 0.2172561, 0.2370263, 0.1818013, 0.1675931, 
    0.1259245, 0.09310087, 0.07336303, 0.07560787, 0.06506167, 0.09201358, 
    0.05657246, 0.0380909, 0.02299978, 0.05429249, 0.07459331,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0002458093, -0.0002365476, 
    -0.0002272859, -0.0002180242, -0.0002087625, -0.0001995008, 
    -0.0001902391, -1.573879e-05, -2.50005e-05, -3.42622e-05, -4.352391e-05, 
    -5.278561e-05, -6.204731e-05, -7.130901e-05, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001385303, 0.1340293, 0.1772728, 
    0.1607335, 0.1843821, 0.1242902, 0.1247705, 0.03203015, 0.02381104, 
    0.02478341, 0.1920608, 0.2436404, 0.2294853, 0.1350814, 0.06123955, 
    0.009301276, 6.530838e-05,
  0.3000757, 0.3319438, 0.3171317, 0.1924275, -0.002867692, -8.261007e-05, 
    0.1310864, 0.002673379, 0.004653442, 0.0366171, 0.05364944, 0.06155575, 
    0.1456896, 0.1650873, 0.2071723, 0.1956522, 0.1360961, 0.2098945, 
    0.2660109, 0.2977964, 0.5200376, 0.3288713, 0.3105363, 0.3062572, 
    0.3736052, 0.185836, 0.1233144, 0.2090007, 0.2994992,
  0.1557633, 0.1955384, 0.2703214, 0.2531469, 0.2797185, 0.2725781, 
    0.2504404, 0.2440801, 0.2138841, 0.2688943, 0.3119731, 0.3064955, 
    0.3392227, 0.247592, 0.2017394, 0.2220665, 0.2311437, 0.241452, 
    0.2882538, 0.3201833, 0.3186872, 0.2750023, 0.3125269, 0.260912, 
    0.2791619, 0.3288402, 0.2233227, 0.1649803, 0.1381772,
  0.2509318, 0.2760779, 0.1794284, 0.18559, 0.1286139, 0.1671612, 0.1637037, 
    0.1360017, 0.1930807, 0.1919296, 0.2087859, 0.2445687, 0.1388667, 
    0.1288012, 0.1133657, 0.08325872, 0.1447816, 0.1348359, 0.1198414, 
    0.1454582, 0.182414, 0.1951084, 0.2110861, 0.2455664, 0.1878644, 
    0.1996304, 0.1706591, 0.2086463, 0.2235744,
  0.1313394, 0.06626981, 0.08160415, 0.07163955, 0.09007212, 0.03218811, 
    0.08782528, 0.05792248, 0.06047798, 0.07682076, 0.09700068, 0.1143213, 
    0.1077294, 0.06683878, 0.09436092, 0.1587067, 0.08304922, 0.08850155, 
    0.137612, 0.2055194, 0.1426353, 0.1170587, 0.1094824, 0.1233444, 
    0.03553703, 0.07794993, 0.08790575, 0.1367019, 0.1990786,
  0.01062273, 0.001467207, 0.01103091, 0.03579488, 0.07820106, 0.04364058, 
    0.01578836, 0.004286055, 0.07851091, 0.03688589, 0.01718523, 0.03015593, 
    0.04790846, 0.02699217, 0.07449279, 0.1162124, 0.1331002, 0.07834455, 
    0.1340254, 0.04207534, 0.04830485, 0.04617143, 0.01122356, 0.09683333, 
    0.0135572, 0.04240821, 0.03542085, 0.0402844, 0.03295621,
  9.748481e-08, 3.67555e-08, 0.0002373487, 0.004112756, 0.05393158, 
    0.02849832, -0.0005869658, 0.01257168, 0.0880182, 0.005819898, 
    1.084059e-05, 1.247321e-06, 0.03959958, 0.09409931, 0.04936418, 
    0.001494191, 0.04844656, 0.01097015, 0.01147731, 0.0007921213, 
    8.498567e-08, 8.81317e-09, 1.458269e-09, 8.997612e-05, 0.001993839, 
    0.0001174743, 0.0004113546, 0.0003470838, 2.907957e-07,
  4.129447e-06, 0.005748174, 0.006639168, 0.09634055, 0.09563505, 0.02082811, 
    0.06282783, 0.008499677, 0.08698528, 0.046141, 0.00510605, 0.003967425, 
    0.1812669, 0.04401528, 0.03593192, 0.01721313, 0.02979106, 0.04266393, 
    0.05948989, 0.02720269, 0.001982889, 4.155361e-06, 9.095536e-05, 
    0.02004789, 0.003402023, 0.0003024099, 0.01887735, -5.427423e-06, 
    7.709962e-07,
  0.01310286, 0.1825054, 0.1513879, 0.01040832, 0.004895024, 0.009019668, 
    0.006362834, 0.006600736, 0.08873869, 0.1316459, 0.01129246, 0.01772057, 
    0.008219787, 0.006319597, 0.01131122, 0.01218977, 0.005172388, 
    0.002308301, 0.002827838, 0.008841438, 0.02142961, 0.02680094, 
    0.04833196, 0.221513, 0.1185348, 0.1869388, 0.1084834, 0.04538333, 
    0.0320501,
  0.05444395, 0.02852966, 0.04910228, 0.02740603, 0.004142083, 0.005516214, 
    0.01205046, 0.005242745, 0.003741684, 0.003699078, 0.006334883, 
    0.007946065, 0.07933372, 0.148174, 0.2410599, 0.15509, 0.05726985, 
    0.01687165, 0.1142638, 0.08140329, 0.01640491, 0.02522221, 0.04492971, 
    0.07584214, 0.01469872, 0.001704928, 0.0004652381, 0.01503922, 0.09943556,
  0.0004946368, 0.03534615, 0.03621854, 0.02007803, 0.002652246, 
    8.131998e-07, 0.004927714, 0.03480563, 0.0466003, 0.2416803, 0.006835082, 
    0.03009073, 0.07694127, 0.0007781707, 0.001119545, 0.0144596, 
    0.0006532724, 0.0007570094, 0.007663677, 0.0004702989, 0.000400668, 
    0.0282739, 0.002588589, 0.04726183, 0.02391745, 0.007742542, 
    7.927846e-05, 0.02610437, 0.01836016,
  0.04615464, 0.05138415, 0.04071362, 0.06028312, 0.03869263, 0.03951075, 
    0.03074635, 0.1686417, 0.3065883, 0.06329719, 0.0856576, 0.1745441, 
    0.1071503, 0.01680503, 0.0004290631, 0.003129299, 0.01163352, 
    0.004366799, 1.149106e-05, 4.908995e-06, 0.002633011, 0.022723, 
    0.03105284, 0.0436698, 0.07161822, 0.0137423, 8.685679e-05, 2.880927e-06, 
    0.002637245,
  0.06308203, 0.02163754, 0.09213029, 0.08302599, 0.09316915, 0.1163004, 
    0.1352522, 0.06714978, 0.09915723, 0.09453939, 0.1313988, 0.07169948, 
    0.1366003, 0.2016459, 0.158987, 0.1908619, 0.09702583, 0.08340356, 
    0.04701216, 0.1212361, 0.1658695, 0.1296132, 0.08172537, 0.1831962, 
    0.183497, 0.1339632, 0.06478351, 0.0601521, 0.03080878,
  0.07833434, 0.103085, 0.09872413, 0.0936565, 0.09644157, 0.1297059, 
    0.1393905, 0.1577307, 0.1840576, 0.1437249, 0.2749477, 0.2096606, 
    0.1777988, 0.08848179, 0.117054, 0.1788335, 0.2574044, 0.1655996, 
    0.1088823, 0.06902642, 0.1590038, 0.1207661, 0.06661128, 0.1462496, 
    0.1815133, 0.1274188, 0.1274139, 0.1374049, 0.1220351,
  0.1900503, 0.1281294, 0.09047835, 0.1702572, 0.1370448, 0.1739946, 
    0.263837, 0.2525335, 0.1958149, 0.2181, 0.1849386, 0.174073, 0.1907134, 
    0.1866407, 0.1639006, 0.1483456, 0.1962035, 0.2828249, 0.1698199, 
    0.1517533, 0.0765924, 0.07827396, 0.04342541, 0.1645295, 0.198953, 
    0.2685047, 0.1401088, 0.185858, 0.1244239,
  0.1907442, 0.1682449, 0.1059579, 0.1116705, 0.1032264, 0.2382942, 
    0.1268181, 0.2323868, 0.1718805, 0.1912962, 0.1316825, 0.1329377, 
    0.1346025, 0.127186, 0.1057083, 0.1600874, 0.148709, 0.1521129, 
    0.1319041, 0.1067429, 0.07758647, 0.04763361, 0.1136593, 0.09200988, 
    0.0824606, 0.1334682, 0.0589511, 0.2102183, 0.2047541,
  0.06038702, 0.09872598, 0.1560039, 0.2042156, 0.197467, 0.1800712, 
    0.07627758, 0.130801, 0.1327786, 0.07171881, 0.05874548, 0.09679459, 
    0.1974639, 0.2085557, 0.2075078, 0.2363869, 0.1612543, 0.1722127, 
    0.1199326, 0.08558309, 0.07172981, 0.07139851, 0.06052048, 0.08384997, 
    0.0452961, 0.04380991, 0.06530418, 0.04424867, 0.05585584,
  4.244298e-05, 4.244298e-05, 4.244298e-05, 4.244298e-05, 4.244298e-05, 
    4.244298e-05, 4.244298e-05, -0.001625399, -0.001060029, -0.0004946587, 
    7.071149e-05, 0.0006360817, 0.001201452, 0.001766822, 0.0004148119, 
    0.0001234467, -0.0001679184, -0.0004592835, -0.0007506486, -0.001042014, 
    -0.001333379, 0.0003927255, 0.0001187205, -0.0001552846, -0.0004292896, 
    -0.0007032947, -0.0009772998, -0.001251305, 4.244298e-05,
  -2.760227e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.338263e-05, 0.01408784, 
    0.1896468, 0.2092115, 0.2262547, 0.2330938, 0.211429, 0.1880931, 
    0.1033239, 0.09232318, 0.08779376, 0.2786008, 0.2642112, 0.249815, 
    0.149325, 0.0811051, 0.0471093, 0.001241599,
  0.3339376, 0.3927763, 0.3923641, 0.273877, 0.003776934, 0.01877858, 
    0.1874755, 0.03954792, 0.03162298, 0.08016925, 0.103562, 0.1234974, 
    0.1703917, 0.176497, 0.2200139, 0.2053956, 0.1990358, 0.235132, 
    0.3145317, 0.2945613, 0.5068222, 0.3375382, 0.3079704, 0.312973, 
    0.3741878, 0.2090182, 0.1277779, 0.2053463, 0.325656,
  0.1482305, 0.2000882, 0.2773523, 0.2567739, 0.30183, 0.2898909, 0.2817396, 
    0.2600985, 0.254786, 0.2598539, 0.3317916, 0.3359778, 0.3469728, 
    0.2440728, 0.1947262, 0.2303193, 0.2411457, 0.2411127, 0.2949627, 
    0.3120857, 0.3070735, 0.2559509, 0.2979483, 0.2258665, 0.2547035, 
    0.3277006, 0.2000602, 0.1606335, 0.1416844,
  0.2480512, 0.2588328, 0.186763, 0.1821588, 0.1086073, 0.1680755, 0.1559168, 
    0.1255715, 0.1809022, 0.1947071, 0.197889, 0.2397398, 0.1434473, 
    0.1190185, 0.1202745, 0.08237088, 0.1377628, 0.1165362, 0.1239439, 
    0.1435808, 0.1731039, 0.1918192, 0.2227415, 0.2310744, 0.1803597, 
    0.1861991, 0.1674842, 0.2342195, 0.2256389,
  0.1267699, 0.05204171, 0.07972187, 0.07275292, 0.07812565, 0.04384659, 
    0.07198311, 0.0598183, 0.05734876, 0.07302841, 0.1001627, 0.1043261, 
    0.1077686, 0.06960272, 0.09827477, 0.1468423, 0.09127358, 0.0922438, 
    0.141462, 0.1700501, 0.1285583, 0.11106, 0.1059216, 0.1321708, 
    0.03065025, 0.06934365, 0.08561211, 0.1347198, 0.1965405,
  0.005427745, 0.001295799, 0.00613264, 0.04215519, 0.07301529, 0.04930184, 
    0.0131248, 0.007330908, 0.08621179, 0.04418375, 0.01717186, 0.02093958, 
    0.04181992, 0.03498287, 0.08778488, 0.1226432, 0.1256943, 0.07794797, 
    0.1316632, 0.04829573, 0.04427607, 0.04911527, 0.01821495, 0.07436062, 
    0.01814857, 0.03828581, 0.03105301, 0.04437698, 0.03044081,
  4.254342e-07, 1.450401e-07, 0.0002120606, 0.001331795, 0.06031262, 
    0.02740758, 0.002700321, 0.002220073, 0.1107236, 0.004341198, 
    1.195611e-05, 1.184485e-07, 0.04334229, 0.09460213, 0.04992408, 
    0.002083803, 0.05173235, 0.01233224, 0.01638411, 0.0009452818, 
    2.617633e-07, 1.710028e-08, 1.109968e-07, 1.750401e-05, 0.003246535, 
    0.0001214102, 0.0003874114, 0.002007649, 1.938375e-07,
  1.560473e-05, 0.004043372, 0.008942555, 0.1130656, 0.1079194, 0.03728152, 
    0.09287596, 0.01120859, 0.08949404, 0.06164194, 0.01110418, 0.003313681, 
    0.2138607, 0.06369331, 0.0474243, 0.02675188, 0.03413845, 0.04540473, 
    0.05057567, 0.03295137, 0.001484474, 2.705278e-07, 0.001081903, 
    0.02200821, 0.004439979, 0.0004160515, 0.03431139, 6.759173e-06, 
    2.800305e-06,
  0.02344204, 0.2100787, 0.1872818, 0.01414699, 0.003670501, 0.008991918, 
    0.007526182, 0.009495068, 0.1185293, 0.1585388, 0.01579465, 0.0196058, 
    0.01190576, 0.00748551, 0.01149487, 0.01237057, 0.006343686, 0.003837814, 
    0.002383641, 0.003649999, 0.02520762, 0.0151142, 0.04989727, 0.2559193, 
    0.1271625, 0.1966304, 0.1130737, 0.04033421, 0.04004808,
  0.0565601, 0.04577287, 0.03726389, 0.04889582, 0.005949821, 0.007522764, 
    0.01302275, 0.006769408, 0.006560924, 0.003558309, 0.005461313, 
    0.00910711, 0.09317017, 0.177048, 0.2816738, 0.181193, 0.07954118, 
    0.02378123, 0.1186703, 0.08014783, 0.02639426, 0.02803105, 0.06457759, 
    0.08718757, 0.01250984, 0.002240079, 0.0004926224, 0.01543655, 0.1241824,
  0.003416469, 0.01390693, 0.01942291, 0.01455011, 0.02240539, 3.695754e-06, 
    0.005414411, 0.03545894, 0.08042108, 0.2732873, 0.008777159, 0.03199878, 
    0.08318505, 0.001047706, 0.00170372, 0.02744917, 0.002522739, 
    0.007668467, 0.001077608, 0.0008491254, 0.004260464, 0.02648505, 
    0.003625166, 0.05500079, 0.02229806, 0.007450433, 4.986926e-05, 
    0.02479474, 0.0100901,
  0.03160294, 0.04325146, 0.02082628, 0.03781918, 0.04140729, 0.02312415, 
    0.02047741, 0.1762813, 0.2980046, 0.05734588, 0.09484925, 0.1800714, 
    0.09835084, 0.01687218, 0.0003180261, 0.003474368, 0.01583491, 
    0.003155752, 3.723302e-06, 1.13417e-06, 0.002463578, 0.01673725, 
    0.02829765, 0.036545, 0.06900106, 0.009404593, 0.0002197261, 
    1.004036e-05, 0.001304161,
  0.0489157, 0.01620811, 0.08668257, 0.08170079, 0.09619456, 0.08746636, 
    0.1287573, 0.06459286, 0.07981228, 0.1083069, 0.1191949, 0.06886648, 
    0.1383943, 0.1873542, 0.1476378, 0.1882045, 0.08111467, 0.07602674, 
    0.05876821, 0.1214607, 0.1942589, 0.1116097, 0.08042854, 0.1737951, 
    0.1851883, 0.1253928, 0.06989902, 0.04463657, 0.03770347,
  0.0798425, 0.09783559, 0.09021804, 0.1065251, 0.09784532, 0.1442958, 
    0.1465501, 0.1598401, 0.188642, 0.1252076, 0.2545694, 0.2049218, 
    0.1787609, 0.08151565, 0.1268113, 0.1886047, 0.2727906, 0.165927, 
    0.09545016, 0.08840782, 0.1416356, 0.1201839, 0.07690591, 0.1672908, 
    0.2015008, 0.1318528, 0.1185206, 0.1581962, 0.1275179,
  0.1817832, 0.1324552, 0.07272877, 0.1764914, 0.1680035, 0.1819441, 
    0.2424919, 0.2817127, 0.2158315, 0.1912027, 0.1820796, 0.1841094, 
    0.2021095, 0.1862038, 0.1615525, 0.1640429, 0.2130704, 0.3099346, 
    0.1706531, 0.1494182, 0.1011852, 0.09175913, 0.05033338, 0.1823094, 
    0.1506097, 0.2945994, 0.1809856, 0.1791108, 0.1278319,
  0.207022, 0.1726856, 0.1239704, 0.1141334, 0.09561407, 0.2319491, 
    0.1281932, 0.2526871, 0.1727992, 0.1925524, 0.1238875, 0.120141, 
    0.1349871, 0.1137152, 0.09094612, 0.1635767, 0.1434021, 0.1611265, 
    0.1168244, 0.1089348, 0.07774804, 0.04074654, 0.1134628, 0.09537033, 
    0.07409216, 0.1345404, 0.1320213, 0.2233509, 0.1951059,
  0.04043823, 0.06315205, 0.1472161, 0.1987455, 0.1850321, 0.1668143, 
    0.06644505, 0.1168558, 0.1378539, 0.08226775, 0.06330042, 0.08129404, 
    0.1530238, 0.208129, 0.2068326, 0.2259799, 0.1499382, 0.1779078, 
    0.1109294, 0.07656649, 0.05746893, 0.0623369, 0.05174905, 0.06370626, 
    0.03726265, 0.04451386, 0.08635088, 0.02385218, 0.03698935,
  0.002817712, 0.002147224, 0.001476735, 0.0008062464, 0.0001357578, 
    -0.0005347308, -0.00120522, -0.001690623, -0.0008375441, 1.553527e-05, 
    0.0008686146, 0.001721694, 0.002574773, 0.003427853, 0.00226682, 
    0.003542034, 0.004817248, 0.006092462, 0.007367677, 0.00864289, 
    0.009918105, 0.005992463, 0.004534659, 0.003076854, 0.001619049, 
    0.000161244, -0.001296561, -0.002754366, 0.003354103,
  -9.475026e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002517459, 0.02964985, 
    0.2342189, 0.2324339, 0.2387823, 0.2730051, 0.2222172, 0.2395076, 
    0.1763038, 0.2148771, 0.1997463, 0.3111653, 0.289538, 0.2452029, 
    0.1473939, 0.08224393, 0.06411993, 0.004493339,
  0.3279002, 0.4464103, 0.3819084, 0.2815592, 0.0588054, 0.04017946, 
    0.2238981, 0.07595399, 0.09697117, 0.2152526, 0.1871629, 0.1794358, 
    0.1683992, 0.1606846, 0.2143199, 0.2111404, 0.2233193, 0.246401, 
    0.3384876, 0.2953424, 0.547192, 0.3497069, 0.3292518, 0.2998922, 
    0.3536234, 0.204077, 0.1271262, 0.225435, 0.3429832,
  0.1742628, 0.2294003, 0.2821914, 0.2617841, 0.3259224, 0.2981414, 0.281316, 
    0.2727966, 0.2536277, 0.3063114, 0.3457467, 0.2984897, 0.3243892, 
    0.2647663, 0.2081873, 0.2398127, 0.232489, 0.2394861, 0.2922508, 
    0.3161514, 0.3089243, 0.2192128, 0.2989056, 0.2640955, 0.2497123, 
    0.308005, 0.2109196, 0.1423887, 0.1577807,
  0.2446015, 0.257765, 0.1736306, 0.1781875, 0.1042053, 0.1618898, 0.1472613, 
    0.1303777, 0.1850297, 0.1879444, 0.2292616, 0.2364302, 0.1429678, 
    0.1225516, 0.1192884, 0.09713579, 0.1271078, 0.1113598, 0.1362772, 
    0.1372025, 0.1895403, 0.1870183, 0.2034659, 0.2180345, 0.1630019, 
    0.1813042, 0.1707455, 0.2317722, 0.2265149,
  0.132742, 0.05091786, 0.08155753, 0.07427564, 0.08211614, 0.04976537, 
    0.09464137, 0.06589352, 0.05878749, 0.1001777, 0.1042948, 0.081821, 
    0.1095371, 0.07836186, 0.1210834, 0.1443694, 0.09285749, 0.08013925, 
    0.1412623, 0.1670513, 0.1347049, 0.1171893, 0.1030461, 0.1319489, 
    0.02691242, 0.06734864, 0.0928374, 0.1302533, 0.1931328,
  0.01091677, 0.001112063, 0.004038778, 0.03930496, 0.06670144, 0.04946052, 
    0.0128795, 0.007618681, 0.09649298, 0.04838926, 0.03002791, 0.0205631, 
    0.04427951, 0.04053776, 0.0835728, 0.1404086, 0.1158534, 0.09000545, 
    0.1400508, 0.05570834, 0.04286584, 0.05057367, 0.02745668, 0.04912956, 
    0.02741079, 0.03140902, 0.02822501, 0.04893602, 0.03294899,
  3.0182e-07, 1.668872e-07, 0.00191966, 0.001369033, 0.07717024, 0.03791254, 
    0.01256891, -2.311279e-05, 0.1165303, 0.002220306, 6.035951e-06, 
    1.786118e-07, 0.04302239, 0.09572717, 0.05288013, 0.002024621, 
    0.06300394, 0.01529543, 0.02740172, 0.003104313, 1.98055e-06, 
    -4.909227e-07, -6.653232e-07, 3.015598e-05, 0.006914867, 0.0002210698, 
    0.0005635711, 0.003676244, 2.260897e-07,
  2.249437e-05, 0.002475378, 0.006611631, 0.1202325, 0.1192566, 0.05071681, 
    0.1127925, 0.01267162, 0.09784613, 0.06700427, 0.02934017, 0.005063201, 
    0.2422209, 0.07109062, 0.04043696, 0.03081573, 0.0341283, 0.04431558, 
    0.05337009, 0.0293821, 0.0008415586, 3.391423e-07, 0.003077651, 
    0.03551362, 0.005719179, 0.000618187, 0.03759368, 0.0002026917, 
    3.989238e-06,
  0.03717611, 0.2608929, 0.2366619, 0.01615441, 0.002734561, 0.007116412, 
    0.008824529, 0.009220032, 0.1410129, 0.2108634, 0.01854947, 0.02437116, 
    0.01267197, 0.008399776, 0.01126935, 0.01107049, 0.009684529, 
    0.003066964, 0.002934688, 0.01399781, 0.03553729, 0.01544776, 0.07419267, 
    0.3009977, 0.1578673, 0.208359, 0.1239069, 0.04334053, 0.04861085,
  0.07498579, 0.0677562, 0.03672042, 0.09421962, 0.005074973, 0.007131502, 
    0.01195364, 0.005650886, 0.009243781, 0.003005149, 0.004635986, 
    0.01255106, 0.1036271, 0.191348, 0.3012118, 0.2033425, 0.09176915, 
    0.0319644, 0.1136168, 0.0762689, 0.02900364, 0.0271189, 0.07989427, 
    0.1170418, 0.01151788, 0.002385952, 0.002079167, 0.02029114, 0.1555038,
  0.00303624, 0.01396731, 0.004002424, 0.009063631, 0.04945091, 5.04326e-06, 
    0.0008797679, 0.02743439, 0.1168356, 0.299641, 0.01356492, 0.03235418, 
    0.08268613, 0.0009267997, 0.002583249, 0.02174965, 0.01095707, 
    0.02394397, 0.000235339, 0.001447584, 0.001217309, 0.02907027, 
    0.003656899, 0.06678189, 0.03061293, 0.0087464, -0.0001260263, 
    0.008598396, 0.003356752,
  0.01838621, 0.02484955, 0.008772263, 0.01923478, 0.04825116, 0.01131028, 
    0.00439281, 0.1551924, 0.2761207, 0.06657422, 0.1003226, 0.1969755, 
    0.1079135, 0.02386752, 0.004126313, 0.007011267, 0.01928934, 0.001500759, 
    3.903697e-06, 1.035193e-06, 0.0006230463, 0.01419243, 0.03177301, 
    0.03612331, 0.0693552, 0.01429382, 0.0001463573, 1.939437e-05, 0.001132461,
  0.04248221, 0.02530639, 0.08698429, 0.07474364, 0.09767815, 0.06033101, 
    0.1329719, 0.04969285, 0.04731828, 0.09632023, 0.1070793, 0.07088136, 
    0.1506888, 0.1816352, 0.1515823, 0.1682588, 0.08661461, 0.08634464, 
    0.04406813, 0.1233541, 0.187089, 0.0927014, 0.07522262, 0.1625149, 
    0.1777723, 0.1269909, 0.08167374, 0.04672276, 0.04305716,
  0.09174829, 0.1106156, 0.09178606, 0.1023888, 0.09893129, 0.1639683, 
    0.1707768, 0.1657983, 0.1998689, 0.1142617, 0.2291301, 0.1979167, 
    0.1835961, 0.06704246, 0.1323773, 0.1743534, 0.2731267, 0.1870933, 
    0.08671877, 0.117813, 0.1444183, 0.1103931, 0.09785882, 0.1752762, 
    0.2252063, 0.1543779, 0.1422588, 0.1679529, 0.1228293,
  0.1835081, 0.127924, 0.0825131, 0.1820045, 0.2041095, 0.1732464, 0.2285311, 
    0.2775036, 0.2190533, 0.1771884, 0.1703332, 0.2019488, 0.2041804, 
    0.1837708, 0.1476351, 0.1966916, 0.2453225, 0.3412633, 0.1773352, 
    0.1535454, 0.1116068, 0.1091925, 0.0657748, 0.2058765, 0.1595029, 
    0.3187654, 0.2065175, 0.1510264, 0.1160047,
  0.2077516, 0.1662148, 0.168154, 0.1167319, 0.1060001, 0.2126148, 0.12641, 
    0.2706648, 0.176744, 0.2056056, 0.1258739, 0.1099446, 0.1211164, 
    0.09049823, 0.0695511, 0.1539577, 0.1487976, 0.1692674, 0.1199753, 
    0.1188828, 0.07704835, 0.04254595, 0.08718879, 0.1046465, 0.06906464, 
    0.1619118, 0.1708373, 0.2221889, 0.2120747,
  0.03465759, 0.07344317, 0.146607, 0.2090847, 0.173833, 0.156396, 
    0.05711321, 0.1051289, 0.136852, 0.08964793, 0.09301186, 0.08751491, 
    0.1491864, 0.2183884, 0.2239372, 0.2345518, 0.1670849, 0.1671572, 
    0.09968553, 0.06201436, 0.04877194, 0.05967559, 0.05440452, 0.05027642, 
    0.03042186, 0.04018144, 0.07408155, 0.02330639, 0.03575904,
  0.06244681, 0.05529452, 0.04814222, 0.04098993, 0.03383764, 0.02668534, 
    0.01953304, 0.02194041, 0.02386414, 0.02578787, 0.02771159, 0.02963532, 
    0.03155904, 0.03348277, 0.02512238, 0.03292669, 0.040731, 0.04853531, 
    0.05633961, 0.06414393, 0.07194823, 0.1204228, 0.1178471, 0.1152714, 
    0.1126956, 0.1101199, 0.1075441, 0.1049684, 0.06816866,
  -0.001292572, -2.575446e-05, -4.372894e-06, 0, 0, 0, 0, 0, 0, 0, 
    -9.880385e-05, 0.006571823, 0.05943272, 0.2902931, 0.2815976, 0.297393, 
    0.3151378, 0.2479314, 0.2659013, 0.289013, 0.3361475, 0.3273998, 
    0.3171487, 0.290815, 0.2355829, 0.1410414, 0.08132929, 0.0605279, 
    0.0219937,
  0.3128211, 0.4426846, 0.3852667, 0.2554449, 0.1118007, 0.05771233, 
    0.2566963, 0.1483693, 0.2120767, 0.3146433, 0.2939515, 0.2568783, 
    0.1649993, 0.1724191, 0.2247946, 0.2120074, 0.2375495, 0.2729803, 
    0.3937641, 0.2892458, 0.5063644, 0.3452729, 0.3004504, 0.2988444, 
    0.3745517, 0.2186311, 0.109349, 0.2038099, 0.3676976,
  0.2268004, 0.2697951, 0.2488354, 0.2752369, 0.3238424, 0.297033, 0.3208252, 
    0.2832863, 0.2759308, 0.2472976, 0.3185514, 0.2995677, 0.3191164, 
    0.3060141, 0.2042126, 0.2219572, 0.239287, 0.2374091, 0.2724574, 
    0.2956128, 0.3028583, 0.247824, 0.3120284, 0.2535583, 0.2500468, 
    0.3017672, 0.2549549, 0.1728058, 0.2105762,
  0.264394, 0.2388096, 0.176952, 0.1719606, 0.1092423, 0.1567656, 0.1424088, 
    0.1751191, 0.2125377, 0.2111809, 0.2294544, 0.2325068, 0.1341918, 
    0.1186167, 0.1119999, 0.08994179, 0.1356896, 0.1306453, 0.1431139, 
    0.1592489, 0.1936992, 0.1720193, 0.1937335, 0.212494, 0.1497902, 
    0.1690057, 0.1574207, 0.2455454, 0.233462,
  0.1423589, 0.05897927, 0.07040384, 0.07978445, 0.09690809, 0.05342636, 
    0.09679545, 0.07570878, 0.06007488, 0.07873035, 0.09859782, 0.08966433, 
    0.1310699, 0.07149033, 0.1160272, 0.1587401, 0.1047882, 0.08794347, 
    0.1356936, 0.1585436, 0.1468977, 0.1220576, 0.1090594, 0.1342439, 
    0.03007713, 0.07184924, 0.09806696, 0.1332054, 0.2224585,
  0.01504956, 0.0008517621, 0.00692737, 0.03909788, 0.05601873, 0.04743471, 
    0.01398587, 0.01432835, 0.1027812, 0.06203701, 0.02060995, 0.0202359, 
    0.04869133, 0.04547959, 0.09549001, 0.142446, 0.1230808, 0.1011934, 
    0.1547929, 0.07405145, 0.03832522, 0.04623295, 0.03041327, 0.02892632, 
    0.03354516, 0.02526952, 0.03026621, 0.05207373, 0.03907607,
  2.234352e-07, -4.905175e-06, 0.01431322, 0.00629692, 0.09383575, 0.0378566, 
    0.01693352, 0.001360716, 0.1098778, 0.000882717, 3.092825e-06, 
    1.601313e-07, 0.04711169, 0.08482517, 0.03727289, 0.00424562, 0.07096618, 
    0.01862432, 0.03949082, 0.009765378, 6.547434e-06, -2.04631e-06, 
    1.835095e-07, 3.699749e-05, 0.01497751, 0.0003356093, 0.001362972, 
    0.009260481, 2.64826e-07,
  2.214059e-05, 0.002111526, 0.009807449, 0.1204023, 0.1153665, 0.05473258, 
    0.1093359, 0.01408827, 0.07926939, 0.04642138, 0.03180205, 0.007623764, 
    0.2458287, 0.05770524, 0.03512448, 0.02659543, 0.03023059, 0.04544543, 
    0.0523274, 0.02135059, 0.0030617, 3.72591e-07, 0.0003395976, 0.05482474, 
    0.007580123, 0.001954291, 0.04652752, 4.560277e-05, 2.816221e-06,
  0.02148033, 0.2821787, 0.2601066, 0.0178835, 0.003253551, 0.005084283, 
    0.008039151, 0.006617886, 0.1483419, 0.2367138, 0.02072412, 0.01823712, 
    0.01271914, 0.007725906, 0.01159123, 0.01280447, 0.01379437, 0.004931048, 
    0.002836127, 0.00620469, 0.0190593, 0.01395763, 0.05001615, 0.29136, 
    0.2083254, 0.1982827, 0.1348038, 0.02979084, 0.02282281,
  0.06446923, 0.04774649, 0.03003946, 0.1315755, 0.00735651, 0.005978405, 
    0.008024362, 0.004595142, 0.007266865, 0.002931412, 0.004975254, 
    0.01261697, 0.08791102, 0.1546614, 0.2587708, 0.1693764, 0.09981431, 
    0.02983537, 0.08089933, 0.06297307, 0.02432887, 0.02546158, 0.08769411, 
    0.1272115, 0.01016928, 0.002366313, 0.004721576, 0.01415734, 0.1647064,
  1.340982e-05, 0.005599292, 0.0003459272, 0.002136455, 0.01723082, 
    9.294589e-06, 0.000332767, 0.01228199, 0.1412507, 0.2290785, 0.00937569, 
    0.01797209, 0.06631725, 0.001836365, 0.005064816, 0.008718832, 
    0.008962108, 0.02467946, 0.0005075392, 0.001427335, 3.819794e-05, 
    0.03500322, 0.003254205, 0.07157164, 0.04023699, 0.00708448, 
    -8.193067e-05, 8.002705e-05, 0.0005669444,
  0.006546606, 0.00722924, 0.005797737, 0.008872881, 0.04224248, 0.004401492, 
    0.0007155612, 0.1263864, 0.287378, 0.07003252, 0.1182041, 0.1886419, 
    0.1036914, 0.01655594, 0.01504434, 0.01064946, 0.02056545, 0.002357464, 
    1.21416e-05, 2.529863e-06, -0.0001353699, 0.01009664, 0.03237284, 
    0.03556564, 0.07363631, 0.01797999, 0.0002370102, 2.596043e-05, 
    0.0002414921,
  0.04670836, 0.03435083, 0.08567768, 0.07720029, 0.09153835, 0.0377584, 
    0.1349033, 0.04017249, 0.03245512, 0.07982986, 0.1005891, 0.07141273, 
    0.1583106, 0.1841801, 0.1619607, 0.172173, 0.0929571, 0.1068091, 
    0.05420615, 0.1277483, 0.172545, 0.0868111, 0.08184312, 0.1604716, 
    0.1830585, 0.1261846, 0.08669954, 0.05078117, 0.04193033,
  0.09752432, 0.1043238, 0.08658274, 0.09160641, 0.1004703, 0.1647119, 
    0.1584447, 0.1779099, 0.1887505, 0.1041772, 0.2192414, 0.1897031, 
    0.1753695, 0.06664252, 0.1360837, 0.1922583, 0.2605726, 0.2028243, 
    0.0891249, 0.1430759, 0.1379401, 0.1287095, 0.1273167, 0.1778127, 
    0.2201969, 0.1822049, 0.1350857, 0.1687474, 0.1169787,
  0.1837737, 0.1340772, 0.07248839, 0.197706, 0.2027901, 0.179045, 0.2352428, 
    0.2795428, 0.2332643, 0.1875436, 0.1498679, 0.2015157, 0.207745, 
    0.1871765, 0.151172, 0.284878, 0.2412664, 0.3733458, 0.1931804, 
    0.1590226, 0.1326651, 0.1502435, 0.08102177, 0.2199936, 0.1559956, 
    0.3321965, 0.2102238, 0.1864898, 0.1470299,
  0.217771, 0.1505335, 0.1878899, 0.0923447, 0.1239501, 0.1906042, 0.1235506, 
    0.289624, 0.1808392, 0.2152241, 0.1209385, 0.1029027, 0.1079435, 
    0.06445115, 0.05369573, 0.1330764, 0.1399608, 0.1686068, 0.1036321, 
    0.122686, 0.06872915, 0.0516794, 0.08858857, 0.08741347, 0.0859488, 
    0.1752306, 0.1788184, 0.2219322, 0.2087416,
  0.03755607, 0.07199845, 0.1494063, 0.2499879, 0.1895557, 0.1539736, 
    0.06411456, 0.1196583, 0.134863, 0.1069794, 0.1048221, 0.130958, 
    0.1758411, 0.2321884, 0.2422781, 0.3108756, 0.2271681, 0.2022296, 
    0.1049734, 0.05544406, 0.04821385, 0.0669729, 0.04882672, 0.04850378, 
    0.0244533, 0.04624428, 0.07308443, 0.05099357, 0.05413499,
  0.1596455, 0.1557184, 0.1517914, 0.1478644, 0.1439374, 0.1400104, 
    0.1360834, 0.1230768, 0.124515, 0.1259532, 0.1273914, 0.1288296, 
    0.1302679, 0.1317061, 0.1229782, 0.1299295, 0.1368809, 0.1438322, 
    0.1507836, 0.1577349, 0.1646863, 0.1918314, 0.1873689, 0.1829063, 
    0.1784438, 0.1739812, 0.1695187, 0.1650561, 0.1627871,
  0.01434967, -0.0008734533, -1.743503e-05, 0, 0, 0, 0, 0, 0, 0, 
    -0.0005938916, 0.06128438, 0.1525715, 0.3050476, 0.2868837, 0.2987906, 
    0.3029579, 0.2259104, 0.2710673, 0.3190928, 0.3858949, 0.4142735, 
    0.3380404, 0.2962872, 0.2291767, 0.1487956, 0.08977766, 0.06245167, 
    0.05228568,
  0.3327585, 0.4492857, 0.3845511, 0.3003829, 0.1605052, 0.06636014, 
    0.2534381, 0.2376005, 0.3054515, 0.3500866, 0.3231104, 0.287281, 
    0.1666398, 0.1992855, 0.2717174, 0.2208806, 0.2662074, 0.308976, 
    0.4036997, 0.3657753, 0.4886365, 0.3625996, 0.2774448, 0.3346053, 
    0.3790117, 0.1882182, 0.127324, 0.2083317, 0.3717273,
  0.2274711, 0.2842176, 0.2440483, 0.2765964, 0.2934735, 0.3094516, 
    0.3204312, 0.2961187, 0.265575, 0.3383828, 0.3352322, 0.2787, 0.2718542, 
    0.2603347, 0.1909614, 0.2304393, 0.2324556, 0.2463243, 0.280388, 
    0.3442447, 0.3329795, 0.2537729, 0.2936649, 0.2317596, 0.2675567, 
    0.292044, 0.196159, 0.1795854, 0.2106598,
  0.2675213, 0.2332435, 0.1766118, 0.1579202, 0.1171755, 0.15571, 0.1405012, 
    0.1698821, 0.2052241, 0.2260196, 0.2145869, 0.2336809, 0.1346715, 
    0.1430046, 0.1071392, 0.08816563, 0.1481858, 0.1139488, 0.1433234, 
    0.1878184, 0.2032752, 0.1570638, 0.1788244, 0.2095053, 0.1384289, 
    0.161283, 0.1552507, 0.2465799, 0.239865,
  0.1562921, 0.06592651, 0.06750432, 0.08486912, 0.112382, 0.06927028, 
    0.1126838, 0.07323696, 0.06140994, 0.09197076, 0.1197001, 0.1042339, 
    0.1368301, 0.07714421, 0.1574025, 0.1604122, 0.1077459, 0.09703109, 
    0.1372499, 0.159903, 0.1649344, 0.1165906, 0.1140577, 0.1382931, 
    0.03892342, 0.08200457, 0.1138455, 0.1356346, 0.2106591,
  0.01873222, 0.0009181503, 0.01743912, 0.03445822, 0.06255157, 0.04563542, 
    0.0179407, 0.02223048, 0.1009647, 0.0659705, 0.0189027, 0.02362271, 
    0.05145539, 0.0511496, 0.1040369, 0.1469502, 0.1311553, 0.1186684, 
    0.1485928, 0.08776305, 0.03711896, 0.04997792, 0.03589503, 0.01465916, 
    0.04681008, 0.02375078, 0.03280738, 0.05377126, 0.04501477,
  8.55666e-08, 6.968335e-05, 0.02189646, 0.01651387, 0.1221784, 0.04412472, 
    0.02373022, 0.003878527, 0.08539408, 0.0006755455, 6.91967e-07, 
    1.135131e-07, 0.04421623, 0.06376083, 0.03177391, 0.003504022, 
    0.07398736, 0.02312325, 0.05054915, 0.01551924, 0.001226598, 
    -4.427254e-06, -1.631867e-06, 3.764971e-05, 0.01883131, 0.0004908711, 
    0.006146614, 0.01288202, 2.484138e-07,
  1.41615e-05, 0.00248761, 0.02092018, 0.1093697, 0.1050923, 0.05458316, 
    0.1081309, 0.0180977, 0.0677861, 0.03623321, 0.02907948, 0.01153324, 
    0.2422268, 0.04420671, 0.03416098, 0.02918604, 0.02913268, 0.04637356, 
    0.04827123, 0.01737859, 0.003757095, 1.425796e-07, 3.581576e-05, 
    0.04562937, 0.007703762, 0.006423494, 0.06631018, 6.84881e-05, 
    8.619746e-07,
  0.0127205, 0.1893025, 0.2038671, 0.02835439, 0.003938058, 0.005980402, 
    0.00767639, 0.005797269, 0.1357508, 0.2175918, 0.02509197, 0.01677018, 
    0.01270004, 0.00802361, 0.01446831, 0.01405065, 0.01632968, 0.006455388, 
    0.002574909, 0.002999775, 0.01976117, 0.002648719, 0.0472449, 0.2588704, 
    0.1984634, 0.1768833, 0.1419369, 0.02197228, 0.01092617,
  0.04181618, 0.02126165, 0.01846892, 0.1566927, 0.006968374, 0.004903776, 
    0.002937885, 0.003867701, 0.005667666, 0.003180647, 0.005887331, 
    0.0105984, 0.07951363, 0.1398431, 0.2308138, 0.1364387, 0.1041213, 
    0.02957978, 0.06259903, 0.05288792, 0.0121158, 0.02333542, 0.08236673, 
    0.08781474, 0.01032781, 0.002726355, 0.006016226, 0.004105486, 0.0897081,
  -3.05825e-06, 0.00155184, 1.828338e-05, 3.150135e-05, 0.001429991, 
    1.206847e-05, 0.0001876407, 0.007941707, 0.1247303, 0.1796802, 
    0.00663304, 0.01281347, 0.05758889, 0.005335638, 0.009925632, 
    0.008511058, 0.02467685, 0.02102263, 0.0001985643, 0.0001360025, 
    1.007844e-05, 0.0351397, 0.003614577, 0.04105337, 0.02950198, 
    0.006711828, 3.410273e-07, 7.217614e-06, 6.836225e-05,
  0.001435288, 0.003631503, 0.004049812, 0.003415229, 0.03169171, 
    0.001492105, -0.0009275224, 0.08231048, 0.3093773, 0.05758221, 0.1133011, 
    0.1855621, 0.09417668, 0.02059171, 0.03016754, 0.01426246, 0.02771172, 
    0.003183774, -3.342164e-05, 2.190968e-06, -2.249189e-05, 0.007396148, 
    0.03501562, 0.03726856, 0.07982661, 0.01791155, 0.001147725, 
    2.967328e-05, -2.262117e-05,
  0.03922241, 0.04261111, 0.09594743, 0.07989924, 0.0841069, 0.03595049, 
    0.1404299, 0.03384746, 0.01848296, 0.05996491, 0.1007583, 0.08758847, 
    0.168722, 0.1942816, 0.1737569, 0.1772642, 0.1101936, 0.1220423, 
    0.04952168, 0.1497605, 0.1692445, 0.09155139, 0.1084331, 0.1817056, 
    0.1872193, 0.1260593, 0.0962467, 0.0635981, 0.04459443,
  0.09447286, 0.124369, 0.0919962, 0.1070076, 0.1269204, 0.1819872, 
    0.1567194, 0.1902067, 0.162024, 0.1092444, 0.2337198, 0.1893506, 
    0.1989357, 0.07426332, 0.1415455, 0.2155668, 0.2771896, 0.2135816, 
    0.1260178, 0.1521492, 0.1629983, 0.1332535, 0.1345149, 0.2372344, 
    0.2245649, 0.1696984, 0.1172178, 0.1845459, 0.1504535,
  0.1858848, 0.1374863, 0.08397242, 0.2293086, 0.2523182, 0.1847185, 
    0.2291024, 0.2836293, 0.2405838, 0.2179106, 0.1550295, 0.2631649, 
    0.1878601, 0.1971422, 0.1738687, 0.3290404, 0.2589009, 0.4376729, 
    0.2489562, 0.1690531, 0.1434684, 0.1616225, 0.05714628, 0.243512, 
    0.1345002, 0.3174025, 0.2510505, 0.1667424, 0.1231167,
  0.2506115, 0.1492415, 0.1693983, 0.09695737, 0.1545895, 0.2015883, 
    0.1207779, 0.2979882, 0.2053477, 0.2120064, 0.1044909, 0.1057873, 
    0.100727, 0.05153377, 0.05645467, 0.1810543, 0.1976516, 0.1731975, 
    0.08708756, 0.1016045, 0.06852605, 0.05110878, 0.1028399, 0.1006824, 
    0.05644296, 0.1825431, 0.1623111, 0.211827, 0.2631498,
  0.07716425, 0.1235153, 0.1932561, 0.2788536, 0.222564, 0.1860937, 
    0.1187435, 0.1560886, 0.1752882, 0.1398821, 0.1210819, 0.1241737, 
    0.2563379, 0.3099282, 0.322514, 0.3061439, 0.2857561, 0.196631, 
    0.1305153, 0.06867637, 0.05874915, 0.09405805, 0.05774135, 0.04419881, 
    0.03314571, 0.04646013, 0.07422678, 0.07880288, 0.0790941,
  0.2365951, 0.235928, 0.2352609, 0.2345938, 0.2339268, 0.2332597, 0.2325926, 
    0.230465, 0.2337214, 0.2369779, 0.2402343, 0.2434907, 0.2467472, 
    0.2500036, 0.2288052, 0.2322092, 0.2356132, 0.2390171, 0.2424211, 
    0.245825, 0.249229, 0.2559595, 0.2499662, 0.2439729, 0.2379796, 
    0.2319863, 0.225993, 0.2199997, 0.2371287,
  0.0607516, 0.002980232, -0.0003709366, 0, 0, -0.0004704371, 0, 0, 0, 
    5.370382e-05, 0.01912832, 0.1685901, 0.192488, 0.3536036, 0.2813194, 
    0.2524238, 0.2153077, 0.2066018, 0.2321192, 0.2741541, 0.4352454, 
    0.5111104, 0.333803, 0.2792017, 0.2129111, 0.1346076, 0.08878717, 
    0.07351282, 0.05981415,
  0.3179186, 0.4035793, 0.423049, 0.2899843, 0.1791379, 0.06553802, 
    0.2638962, 0.3199246, 0.3269794, 0.3860629, 0.3817465, 0.2967629, 
    0.1624587, 0.1956648, 0.2882868, 0.2409213, 0.2818858, 0.2872551, 
    0.3600112, 0.3594923, 0.4302439, 0.4201106, 0.3592381, 0.3785615, 
    0.38438, 0.2078879, 0.1532069, 0.2080938, 0.3895988,
  0.2320417, 0.2955049, 0.2489041, 0.2797572, 0.3013349, 0.3269636, 0.330947, 
    0.3118108, 0.3013995, 0.3286505, 0.3882799, 0.2703768, 0.2693276, 
    0.2852175, 0.2172192, 0.242812, 0.2476502, 0.2725729, 0.3221798, 
    0.3580115, 0.3331153, 0.2764585, 0.2896362, 0.2956507, 0.3584688, 
    0.4009981, 0.2653198, 0.1597818, 0.2288861,
  0.2710178, 0.236643, 0.1858833, 0.1687503, 0.128229, 0.1661132, 0.1499196, 
    0.2030619, 0.2262098, 0.2356365, 0.212781, 0.2269631, 0.154841, 
    0.1377076, 0.1044043, 0.1047927, 0.1676827, 0.1366344, 0.1582041, 
    0.207854, 0.2211888, 0.1610219, 0.1844089, 0.2198657, 0.1279851, 
    0.1581277, 0.1820671, 0.2717744, 0.2513323,
  0.1847639, 0.06676202, 0.07540171, 0.08880618, 0.1344778, 0.08646506, 
    0.1483357, 0.0932452, 0.06878012, 0.1139491, 0.1195074, 0.1294506, 
    0.1566375, 0.1045603, 0.2027329, 0.1888376, 0.1179025, 0.107794, 
    0.1418817, 0.1742992, 0.1704543, 0.1209071, 0.1300951, 0.1434741, 
    0.04576887, 0.09751257, 0.1357944, 0.1427129, 0.2156358,
  0.02795631, 0.001735536, 0.09039535, 0.03296021, 0.05585314, 0.04460908, 
    0.02427418, 0.0258912, 0.105225, 0.05116307, 0.01151873, 0.02119947, 
    0.06834086, 0.04833708, 0.1196991, 0.1632053, 0.1274413, 0.1439791, 
    0.1461254, 0.07295369, 0.04312452, 0.04948836, 0.04417235, 0.009791108, 
    0.06014279, 0.02372295, 0.03891528, 0.05747509, 0.05357246,
  9.916905e-08, 0.009068388, 0.03587351, 0.01808581, 0.1310295, 0.05859457, 
    0.03871551, 0.007665778, 0.07535739, 0.0006549702, 2.56881e-07, 
    4.179774e-05, 0.03984138, 0.05534525, 0.02901912, 0.007492375, 
    0.06597272, 0.03427827, 0.05196395, 0.0317738, 0.0104786, 0.001471546, 
    -0.0002162966, 2.114656e-05, 0.03047978, 0.001922333, 0.01228854, 
    0.02242592, -1.658769e-06,
  5.867803e-06, 0.006422543, 0.02781361, 0.10235, 0.1008862, 0.06130243, 
    0.09825675, 0.02377577, 0.06256833, 0.02932633, 0.04013412, 0.01782601, 
    0.235436, 0.04525111, 0.03466067, 0.03091283, 0.03178639, 0.04869692, 
    0.03570979, 0.01997085, 0.001585927, 1.174942e-06, 7.57482e-06, 
    0.04724174, 0.009004644, 0.07436261, 0.09806458, 0.0004962381, 
    3.922134e-07,
  0.01162829, 0.1416176, 0.1893983, 0.05147413, 0.004462234, 0.007171847, 
    0.008631037, 0.006725177, 0.1484329, 0.2105148, 0.0288794, 0.01829621, 
    0.01422986, 0.009624807, 0.01642744, 0.01711833, 0.01410707, 0.008016867, 
    0.004983856, 0.004139753, 0.01246174, 0.002879835, 0.04010796, 0.2367367, 
    0.199017, 0.1575906, 0.1406601, 0.02577598, 0.009127988,
  0.03002405, 0.009985811, 0.01900192, 0.1548828, 0.01042749, 0.00441355, 
    0.001702068, 0.003942468, 0.005716672, 0.003903792, 0.008481793, 
    0.01201858, 0.07398619, 0.1347955, 0.2071987, 0.1145885, 0.1194295, 
    0.03547788, 0.06186296, 0.05603848, 0.01291745, 0.02036072, 0.08360829, 
    0.06801223, 0.01417435, 0.002899957, 0.006406839, 0.0007168327, 0.06397404,
  4.607451e-07, 0.0002678837, 5.268368e-06, -2.614733e-05, 0.0001736699, 
    9.636144e-06, 6.113474e-05, 0.004698048, 0.1258295, 0.1512532, 
    0.008891284, 0.01188208, 0.04828819, 0.01204671, 0.02430559, 0.02298316, 
    0.03983224, 0.02872213, 2.217255e-05, 1.385977e-05, 4.06784e-06, 
    0.03537936, 0.005026414, 0.02921288, 0.03120737, 0.014762, 0.000176724, 
    4.647556e-06, 2.303813e-06,
  8.144297e-05, 0.001384923, 0.002067053, 0.001054669, 0.01977304, 
    0.0002638053, -0.0009510433, 0.04963476, 0.311666, 0.05660853, 0.1026535, 
    0.1889494, 0.08599905, 0.02444652, 0.04268221, 0.02799559, 0.04056873, 
    0.002258698, 0.005327164, 3.579682e-06, -0.0001480601, 0.008764223, 
    0.03182047, 0.03885293, 0.07041317, 0.02841174, 0.003249842, 5.60967e-05, 
    -2.644778e-05,
  0.02938585, 0.04893157, 0.1046655, 0.08357636, 0.07898824, 0.03318411, 
    0.1379365, 0.02095104, 0.008163569, 0.03771368, 0.1068759, 0.09619261, 
    0.174096, 0.2033819, 0.1709278, 0.1966042, 0.1105111, 0.1257877, 
    0.06505983, 0.1646156, 0.163353, 0.09301573, 0.1499603, 0.1865701, 
    0.190575, 0.1413262, 0.1044689, 0.0889364, 0.06189698,
  0.1221184, 0.1274037, 0.1174187, 0.1303061, 0.1462277, 0.1892176, 
    0.1554848, 0.2165862, 0.1413344, 0.1150949, 0.2557936, 0.1965635, 
    0.2299673, 0.08868449, 0.1299962, 0.2472976, 0.2913462, 0.2191591, 
    0.105443, 0.1608104, 0.1763884, 0.1431346, 0.1231994, 0.2647419, 
    0.2493396, 0.2251014, 0.1507226, 0.1917345, 0.1666444,
  0.2537963, 0.1605448, 0.1465191, 0.2349964, 0.2658635, 0.2431452, 
    0.2643197, 0.2658896, 0.2762989, 0.2553826, 0.2608552, 0.3352344, 
    0.1818926, 0.2157421, 0.2805316, 0.4950522, 0.3584804, 0.4589258, 
    0.2463786, 0.1976555, 0.1416458, 0.1712828, 0.09580933, 0.2750149, 
    0.2003058, 0.320433, 0.2724718, 0.1999401, 0.1624569,
  0.2990792, 0.1431689, 0.1930929, 0.08043285, 0.1963628, 0.2594685, 
    0.09995956, 0.2711315, 0.2183892, 0.2306402, 0.1675515, 0.1634277, 
    0.1246671, 0.08702584, 0.09937721, 0.2446766, 0.2858998, 0.1890627, 
    0.1007279, 0.1068818, 0.08527037, 0.04242534, 0.1116374, 0.111645, 
    0.05045627, 0.1861541, 0.1548553, 0.2013289, 0.349192,
  0.08517937, 0.1636944, 0.1792335, 0.2238968, 0.2402022, 0.1762485, 
    0.1445016, 0.1794942, 0.2102112, 0.1516783, 0.1353661, 0.1442613, 
    0.301117, 0.3828958, 0.3852794, 0.349033, 0.2121807, 0.1699455, 
    0.1147763, 0.07293624, 0.1132077, 0.1305997, 0.08672138, 0.05657648, 
    0.05173772, 0.04790034, 0.0644707, 0.114682, 0.1320717,
  0.2527589, 0.2539192, 0.2550794, 0.2562396, 0.2573999, 0.2585601, 
    0.2597203, 0.2549865, 0.2575714, 0.2601563, 0.2627412, 0.2653261, 
    0.267911, 0.270496, 0.2616542, 0.2683358, 0.2750175, 0.2816991, 
    0.2883807, 0.2950624, 0.301744, 0.3402299, 0.3298031, 0.3193763, 
    0.3089496, 0.2985228, 0.288096, 0.2776692, 0.2518308,
  0.1002498, 0.03602106, 0.01169187, -3.167781e-05, 0, -0.003589754, 
    -1.059941e-05, -2.338721e-05, 6.897345e-06, 0.0069311, 0.08770656, 
    0.1516761, 0.238071, 0.3482469, 0.1644833, 0.1761079, 0.1917385, 
    0.1530909, 0.1656108, 0.2253156, 0.4774626, 0.5535511, 0.3466633, 
    0.2676304, 0.2250524, 0.1207745, 0.0823253, 0.08426204, 0.06245217,
  0.2954314, 0.3897161, 0.3924506, 0.2646905, 0.2078453, 0.0607509, 
    0.2956592, 0.3344909, 0.3756418, 0.3811811, 0.4067681, 0.2914767, 
    0.1429195, 0.2261582, 0.279401, 0.2620231, 0.2501831, 0.242047, 
    0.3076166, 0.3068546, 0.4314465, 0.3344983, 0.3161911, 0.3604918, 
    0.3281239, 0.1888342, 0.127209, 0.1734215, 0.3658467,
  0.2466127, 0.2688145, 0.2571447, 0.2923837, 0.2770335, 0.341161, 0.3373353, 
    0.3069623, 0.3195248, 0.36854, 0.3578355, 0.2934951, 0.2698973, 
    0.2864694, 0.2268666, 0.2677507, 0.2644829, 0.2815823, 0.3493395, 
    0.3795419, 0.3187629, 0.2628437, 0.3063265, 0.2766837, 0.3342271, 
    0.3437216, 0.2703343, 0.1370809, 0.2279946,
  0.2599768, 0.248499, 0.2073061, 0.1782671, 0.1415474, 0.1999119, 0.179307, 
    0.2209684, 0.2480479, 0.260551, 0.2310437, 0.2479682, 0.1803882, 
    0.1276084, 0.1381399, 0.1385678, 0.1853441, 0.1644122, 0.2041837, 
    0.2208612, 0.2406503, 0.1733726, 0.2293703, 0.2312086, 0.1212859, 
    0.1726429, 0.196811, 0.2977049, 0.2558508,
  0.1929203, 0.08241491, 0.08887863, 0.09636253, 0.1628727, 0.09571597, 
    0.1498284, 0.1130551, 0.1159934, 0.1518708, 0.1401963, 0.1374591, 
    0.1727723, 0.1331649, 0.2302913, 0.2412869, 0.1619723, 0.118289, 
    0.1567699, 0.1850544, 0.1850513, 0.129178, 0.1434207, 0.153411, 
    0.05943934, 0.1162675, 0.1584804, 0.1631853, 0.2370118,
  0.03735573, 0.003309583, 0.05503256, 0.04516986, 0.0422426, 0.04937851, 
    0.03730917, 0.03660565, 0.1114391, 0.0346125, 0.006936722, 0.008781403, 
    0.0790183, 0.05472626, 0.1148681, 0.1577751, 0.1146032, 0.1723343, 
    0.1597978, 0.07775436, 0.05604767, 0.07805355, 0.04382665, 0.008665849, 
    0.07355032, 0.0341805, 0.05275943, 0.06066084, 0.0646119,
  8.973507e-07, 0.0003727646, 0.0627862, 0.02281004, 0.1241531, 0.05200046, 
    0.05686208, 0.0245949, 0.07239089, 0.0008776482, 1.064619e-07, 
    0.001035841, 0.04142675, 0.07072981, 0.02634622, 0.01033194, 0.07081439, 
    0.04583336, 0.05085379, 0.06554641, 0.01588435, 0.01291649, 0.009088163, 
    7.243196e-06, 0.03673194, 0.006169897, 0.02839165, 0.04301665, 
    0.0009527809,
  3.881833e-06, 0.01765137, 0.02713366, 0.09635022, 0.09683616, 0.06367189, 
    0.09100296, 0.03091985, 0.06037546, 0.03192313, 0.0501749, 0.02790468, 
    0.2407637, 0.04547544, 0.03671219, 0.03204866, 0.03046656, 0.05143461, 
    0.03560217, 0.02127232, 0.0008898982, 0.0001932, 2.686022e-06, 
    0.04639974, 0.01086876, 0.2112223, 0.1343646, 0.001524238, 5.671258e-07,
  0.01284104, 0.1178012, 0.168978, 0.0854567, 0.005653055, 0.007629774, 
    0.01028189, 0.007351078, 0.1664003, 0.2300715, 0.0301844, 0.02020148, 
    0.01579597, 0.01100041, 0.01810072, 0.02070935, 0.01581088, 0.01160175, 
    0.01225794, 0.008183459, 0.00342124, 0.001994841, 0.0364035, 0.2384162, 
    0.191932, 0.1409865, 0.1410879, 0.0323556, 0.01129893,
  0.02158838, 0.007904638, 0.009695003, 0.1323155, 0.01106447, 0.004458527, 
    0.002510212, 0.004541294, 0.005602754, 0.00490694, 0.01517904, 
    0.01465064, 0.07015564, 0.1249659, 0.1758517, 0.1107719, 0.1199733, 
    0.0477266, 0.07902029, 0.06562643, 0.01860602, 0.01883996, 0.087169, 
    0.06302419, 0.01969049, 0.004582844, 0.00806549, 3.977917e-05, 0.04509008,
  6.455727e-07, 2.734483e-05, 2.694698e-06, -1.97016e-05, 2.919335e-05, 
    6.138524e-06, 4.297598e-05, 0.001721317, 0.1402674, 0.1380682, 
    0.01369215, 0.01462202, 0.04977402, 0.02526913, 0.02723142, 0.03541302, 
    0.0388081, 0.03532825, 4.388077e-06, 4.262721e-06, 1.24596e-06, 
    0.0345977, 0.005942939, 0.02580977, 0.02833887, 0.03113515, 0.006222345, 
    2.1049e-06, 5.820618e-07,
  1.090607e-05, 0.0008058799, 0.0005797259, 0.0001325569, 0.0110872, 
    2.269978e-05, -0.0007671798, 0.03389212, 0.286307, 0.06430803, 
    0.08429386, 0.1762461, 0.08122527, 0.03932353, 0.04516497, 0.02980548, 
    0.05188828, 0.005931426, 0.005286629, 2.457808e-05, -6.918817e-05, 
    0.008196412, 0.0208679, 0.0638035, 0.06402214, 0.0330145, 0.007902059, 
    8.954723e-05, -2.908874e-06,
  0.01985136, 0.03552181, 0.1045689, 0.09104817, 0.04409564, 0.01290627, 
    0.1231369, 0.01703238, 0.002932254, 0.02684931, 0.1193193, 0.09927738, 
    0.1743696, 0.1933581, 0.148694, 0.1936653, 0.1141723, 0.1348874, 
    0.08173075, 0.1785595, 0.1380063, 0.1042998, 0.1656037, 0.1798685, 
    0.1923351, 0.1576426, 0.1185557, 0.09558214, 0.07400671,
  0.1772147, 0.1405014, 0.1211509, 0.1580358, 0.1478094, 0.153711, 0.1298047, 
    0.215511, 0.1152915, 0.1119953, 0.2544423, 0.2449552, 0.2152432, 
    0.09144856, 0.1326036, 0.2425322, 0.2602959, 0.2459883, 0.1077202, 
    0.1720828, 0.1730263, 0.0952253, 0.1559838, 0.2551297, 0.2209135, 
    0.2437786, 0.1794901, 0.2029545, 0.1640356,
  0.2935513, 0.2079663, 0.1640397, 0.2668491, 0.3077522, 0.2918573, 
    0.2896087, 0.2682517, 0.2408024, 0.2550725, 0.2620836, 0.352354, 
    0.1947421, 0.2054762, 0.1926575, 0.3974137, 0.4223817, 0.475986, 
    0.2036954, 0.1901839, 0.1219386, 0.1456959, 0.1145292, 0.2619502, 
    0.1357814, 0.3010169, 0.2578211, 0.2255952, 0.243403,
  0.2338981, 0.1194026, 0.2218512, 0.1128891, 0.1841804, 0.2364917, 
    0.08764271, 0.2762721, 0.2622761, 0.2385449, 0.1916906, 0.167849, 
    0.09002902, 0.1132616, 0.1075868, 0.189314, 0.2098909, 0.1571044, 
    0.09104355, 0.1042187, 0.07955824, 0.05254781, 0.1765908, 0.1331145, 
    0.05865643, 0.188706, 0.1495235, 0.181247, 0.3499921,
  0.09919968, 0.1407987, 0.1602099, 0.1561459, 0.1574941, 0.1365937, 
    0.1101316, 0.1386276, 0.1675776, 0.1185692, 0.1090744, 0.1233484, 
    0.2355277, 0.3441114, 0.2635581, 0.3230933, 0.1868718, 0.1457228, 
    0.07305375, 0.05065285, 0.07032768, 0.2039542, 0.1371755, 0.1235049, 
    0.0746962, 0.06099052, 0.07670094, 0.1103108, 0.1032463,
  0.3013707, 0.3044307, 0.3074907, 0.3105508, 0.3136108, 0.3166708, 
    0.3197309, 0.330064, 0.3359181, 0.3417721, 0.3476262, 0.3534802, 
    0.3593343, 0.3651883, 0.3486566, 0.351932, 0.3552075, 0.358483, 
    0.3617584, 0.3650339, 0.3683093, 0.3738808, 0.3616913, 0.3495017, 
    0.3373122, 0.3251226, 0.3129331, 0.3007435, 0.2989227,
  0.1283372, 0.1003454, 0.03436863, 0.01160169, -0.001377295, 0.0002432973, 
    -0.002616363, -0.0007647023, 0.001273462, 0.02798119, 0.1542528, 
    0.1712876, 0.2600492, 0.3032303, 0.2214101, 0.2311022, 0.1962228, 
    0.1519821, 0.1093698, 0.2053743, 0.5383394, 0.5483487, 0.3200155, 
    0.2466118, 0.2775078, 0.1032421, 0.08228271, 0.08692188, 0.09166024,
  0.378256, 0.4111258, 0.3400834, 0.253464, 0.2240623, 0.05941621, 0.3038222, 
    0.3611006, 0.4040587, 0.3651265, 0.439558, 0.2901806, 0.1461201, 
    0.2327086, 0.3003352, 0.2857377, 0.2414205, 0.286794, 0.338251, 
    0.2750801, 0.4073521, 0.2947029, 0.3047874, 0.3191599, 0.2984383, 
    0.1511746, 0.1300064, 0.2005543, 0.3889647,
  0.2727666, 0.2701465, 0.2604422, 0.2693652, 0.2579924, 0.3430851, 
    0.3441791, 0.3358035, 0.310921, 0.3487104, 0.2930847, 0.32321, 0.3056549, 
    0.2945356, 0.2454229, 0.2734111, 0.2717134, 0.2963935, 0.3195132, 
    0.3723928, 0.3409869, 0.2594361, 0.2840646, 0.2463216, 0.2817224, 
    0.2856458, 0.2121802, 0.1089709, 0.2372934,
  0.2377741, 0.2879961, 0.2254301, 0.1945422, 0.1674159, 0.2190233, 
    0.2021222, 0.2634141, 0.2799706, 0.260448, 0.2595443, 0.2936663, 
    0.1898645, 0.1471283, 0.1863425, 0.1720361, 0.2255831, 0.1976425, 
    0.2281418, 0.2400527, 0.2444136, 0.1815867, 0.2037393, 0.2389075, 
    0.1283849, 0.2122701, 0.2037646, 0.2904208, 0.2396466,
  0.1982478, 0.09868079, 0.09524684, 0.1208627, 0.1729321, 0.09858453, 
    0.1319281, 0.1185123, 0.1667615, 0.1926939, 0.1857295, 0.1311584, 
    0.1677128, 0.1518183, 0.1797113, 0.2582758, 0.1721643, 0.1418634, 
    0.1916951, 0.1946723, 0.1975905, 0.1402794, 0.1575602, 0.172835, 
    0.05500113, 0.1439475, 0.1770401, 0.2016604, 0.2432833,
  0.05016872, 0.003441417, 0.01309108, 0.05534358, 0.03922467, 0.05847643, 
    0.03600115, 0.06470495, 0.1350175, 0.0406528, 0.0143484, 0.004171883, 
    0.04798774, 0.05736431, 0.1033945, 0.1411918, 0.1166077, 0.1829928, 
    0.1888689, 0.07806521, 0.06064628, 0.08232046, 0.0449636, 0.009117099, 
    0.06597814, 0.04104071, 0.07102253, 0.06168472, 0.06590105,
  8.089454e-06, 5.535432e-05, 0.06148732, 0.02301193, 0.1144436, 0.04727379, 
    0.0543539, 0.0333247, 0.06801753, 0.001721165, 2.707876e-08, 0.005164245, 
    0.0494814, 0.06876157, 0.02623627, 0.014344, 0.06254409, 0.05125996, 
    0.0399307, 0.05804979, 0.05000995, 0.04028248, 0.01062711, 3.10349e-05, 
    0.04567373, 0.01490326, 0.03986537, 0.05489719, 0.04382519,
  1.600011e-05, 0.0121761, 0.02394777, 0.1012517, 0.0836555, 0.06585192, 
    0.08773378, 0.03471557, 0.06377593, 0.05349434, 0.07709265, 0.04978388, 
    0.2353817, 0.04140964, 0.03624398, 0.03149893, 0.02791932, 0.05119932, 
    0.03555741, 0.02191922, 0.002803713, 0.002488139, 1.001748e-06, 
    0.04525853, 0.01438785, 0.1128855, 0.1366878, 0.003705426, 3.639068e-06,
  0.02295423, 0.1033512, 0.1404108, 0.0962632, 0.007192689, 0.009002625, 
    0.01118064, 0.008557356, 0.1672826, 0.2334616, 0.02993776, 0.01980227, 
    0.01612522, 0.0117238, 0.01811972, 0.02189784, 0.01600241, 0.01411679, 
    0.01417412, 0.01197985, 0.004267834, 0.003891753, 0.02377061, 0.2337143, 
    0.1835075, 0.1198079, 0.1363504, 0.04452864, 0.01243315,
  0.01750054, 0.006282357, 0.003865829, 0.09824371, 0.008826292, 0.005207932, 
    0.008083924, 0.006676107, 0.007490786, 0.008122698, 0.02272252, 
    0.01617333, 0.07221688, 0.1129931, 0.1493189, 0.1078317, 0.1253098, 
    0.05458426, 0.09961205, 0.06431702, 0.02356771, 0.01925262, 0.08822077, 
    0.06911378, 0.02294184, 0.009106234, 0.009697059, -4.799686e-05, 
    0.02855569,
  5.170709e-07, 1.778356e-06, 1.834724e-06, -1.154055e-05, 4.15095e-06, 
    3.049046e-06, 2.778405e-05, 0.0002200242, 0.1453187, 0.1415465, 
    0.02000713, 0.02133732, 0.04473605, 0.03252042, 0.04169358, 0.02897815, 
    0.04662639, 0.06171869, 0.0003277522, 1.481747e-06, 1.142831e-06, 
    0.03359808, 0.006939804, 0.02365135, 0.0244623, 0.04461702, 0.02443109, 
    -1.153744e-05, 1.3588e-07,
  -3.727884e-05, 0.0001817515, 3.212171e-05, 1.141963e-05, 0.004135448, 
    6.500413e-06, -0.0005911925, 0.01761205, 0.2708232, 0.08463187, 
    0.08946908, 0.1694204, 0.0859779, 0.06860339, 0.04437622, 0.0544798, 
    0.05527668, 0.007396611, 0.006015139, 0.0003651694, -1.235919e-05, 
    0.008661098, 0.01730676, 0.061105, 0.06294804, 0.03315069, 0.01733039, 
    0.003495612, -0.0001262322,
  0.01146728, 0.02767091, 0.09891458, 0.09939735, 0.01558695, 0.007258988, 
    0.1178906, 0.01153867, 0.004812788, 0.01963766, 0.1201161, 0.09306382, 
    0.1916682, 0.1738234, 0.1554332, 0.1975961, 0.1366371, 0.1375042, 
    0.07476501, 0.1777209, 0.1224078, 0.1135415, 0.1676056, 0.1782719, 
    0.191011, 0.1505322, 0.1141769, 0.1204326, 0.07394515,
  0.1416432, 0.1489811, 0.1313753, 0.1722363, 0.06881931, 0.1165087, 
    0.08148362, 0.2175788, 0.09339105, 0.08814635, 0.2620348, 0.2688667, 
    0.2305151, 0.08142198, 0.115531, 0.2332071, 0.2903963, 0.2245197, 
    0.114411, 0.2134098, 0.1530646, 0.06749186, 0.1669662, 0.2893337, 
    0.2116338, 0.2485378, 0.2112011, 0.2291999, 0.1779588,
  0.2479124, 0.2700918, 0.134233, 0.3036998, 0.2860319, 0.2203235, 0.2372854, 
    0.2360635, 0.2293904, 0.256356, 0.2299991, 0.3746438, 0.1898296, 
    0.164183, 0.1786034, 0.2607772, 0.4003207, 0.4941377, 0.2013229, 
    0.1746156, 0.1200364, 0.1241411, 0.08925283, 0.1808173, 0.1030396, 
    0.2699462, 0.2379681, 0.1861857, 0.2186362,
  0.2357818, 0.1549377, 0.2696312, 0.1298706, 0.1427801, 0.152814, 0.1655687, 
    0.2871414, 0.2813672, 0.19358, 0.1540135, 0.1482672, 0.05957081, 
    0.06541747, 0.07650798, 0.1112376, 0.09891458, 0.1091347, 0.07820776, 
    0.08946086, 0.1272969, 0.0459533, 0.1456434, 0.1703762, 0.0530094, 
    0.1903129, 0.146196, 0.1721036, 0.2862174,
  0.05496738, 0.08173295, 0.1052399, 0.1169154, 0.1031677, 0.1453164, 
    0.07589625, 0.09753743, 0.1058621, 0.08805548, 0.1006996, 0.08559469, 
    0.1770411, 0.243267, 0.1648011, 0.2262387, 0.1794704, 0.09741195, 
    0.09527408, 0.07643177, 0.1212728, 0.2220197, 0.1663842, 0.07042626, 
    0.04765902, 0.07254659, 0.1150612, 0.1071843, 0.1312753,
  0.3261281, 0.3284515, 0.3307749, 0.3330983, 0.3354217, 0.3377451, 
    0.3400685, 0.3394687, 0.3461449, 0.3528211, 0.3594974, 0.3661736, 
    0.3728498, 0.379526, 0.370472, 0.374307, 0.378142, 0.381977, 0.3858119, 
    0.3896469, 0.3934819, 0.4225768, 0.4097423, 0.3969077, 0.384073, 
    0.3712384, 0.3584038, 0.3455692, 0.3242694,
  0.1389281, 0.1957614, 0.05401098, 0.0364733, 0.006224372, 0.02714524, 
    0.006853419, -0.0005627868, 0.008737089, 0.04670482, 0.1663568, 
    0.2002166, 0.2913143, 0.2661961, 0.2219125, 0.2596098, 0.197989, 
    0.1392545, 0.09100711, 0.1928163, 0.552188, 0.5596476, 0.3009397, 
    0.2391378, 0.2256592, 0.1195305, 0.1029252, 0.09818723, 0.09215626,
  0.3874147, 0.4308186, 0.3508195, 0.2395739, 0.2402284, 0.064004, 0.2710185, 
    0.3760414, 0.4637498, 0.3860041, 0.4548364, 0.2914363, 0.1504779, 
    0.2403577, 0.300882, 0.2953888, 0.2337835, 0.2992595, 0.3730502, 
    0.3103999, 0.4233466, 0.3357, 0.3757783, 0.3603218, 0.299752, 0.1678432, 
    0.1090277, 0.2076623, 0.3942606,
  0.3314268, 0.3214526, 0.3310663, 0.2910306, 0.2700261, 0.3603272, 
    0.3827499, 0.3884386, 0.3508393, 0.3530035, 0.2992615, 0.3741588, 
    0.3363483, 0.3290839, 0.2941169, 0.3223301, 0.3317877, 0.3352798, 
    0.3480198, 0.3850805, 0.3465172, 0.2797318, 0.3331905, 0.2515717, 
    0.3119624, 0.2751536, 0.1829258, 0.1476124, 0.3166594,
  0.2724655, 0.3134796, 0.2782064, 0.2366357, 0.1955779, 0.2241896, 
    0.2255801, 0.3220789, 0.3132691, 0.2902073, 0.2917083, 0.3006395, 
    0.2286697, 0.2037315, 0.1959094, 0.2069649, 0.272714, 0.2473829, 
    0.2785975, 0.2497534, 0.2672587, 0.1973149, 0.2089089, 0.2639443, 
    0.1702765, 0.2666942, 0.2660755, 0.3390869, 0.25537,
  0.2197278, 0.1232131, 0.1037892, 0.1354892, 0.1570202, 0.1059817, 
    0.1497601, 0.1410309, 0.2151348, 0.2278801, 0.2036544, 0.1347018, 
    0.1738281, 0.173553, 0.2037794, 0.2489241, 0.1788072, 0.1738832, 
    0.2166139, 0.2010666, 0.201099, 0.1518066, 0.1557279, 0.1860785, 
    0.05080973, 0.1667349, 0.2209828, 0.2104804, 0.2390638,
  0.08872972, 0.004626177, 0.008176446, 0.0588158, 0.03841573, 0.09651741, 
    0.04745529, 0.08731142, 0.1630243, 0.08199623, 0.02437492, 0.00754085, 
    0.03855472, 0.08695287, 0.09025399, 0.1657129, 0.1399328, 0.2061262, 
    0.1990366, 0.07789812, 0.06694469, 0.1085796, 0.05539586, 0.009610285, 
    0.05224065, 0.05593732, 0.09323523, 0.1068585, 0.09553718,
  0.005867685, 9.892851e-06, 0.01443969, 0.02540797, 0.1045559, 0.04163225, 
    0.05950842, 0.03151823, 0.06966008, 0.03989494, 3.812326e-09, 
    6.686941e-06, 0.06345841, 0.08360112, 0.03098229, 0.04241585, 0.06810749, 
    0.05429853, 0.02759043, 0.03757517, 0.08527692, 0.0872611, 0.03256943, 
    4.064468e-05, 0.07426629, 0.021393, 0.04087031, 0.06641554, 0.06813952,
  0.000128785, 0.003767411, 0.02428659, 0.1143866, 0.07241131, 0.05495609, 
    0.07714676, 0.03583997, 0.05970125, 0.06159888, 0.08996229, 0.05310867, 
    0.2262049, 0.03381461, 0.03120016, 0.03111514, 0.02471499, 0.0452444, 
    0.03121297, 0.02388241, 0.01225932, 0.0115557, -1.592674e-05, 0.04648091, 
    0.01675542, 0.0234875, 0.1201359, 0.01518526, 0.0006844891,
  0.03248475, 0.1044203, 0.1126518, 0.08394268, 0.008884, 0.01067334, 
    0.01358657, 0.0124408, 0.1533221, 0.228358, 0.02874146, 0.01831966, 
    0.01643933, 0.01261448, 0.01820738, 0.02158915, 0.01736093, 0.01413868, 
    0.01424024, 0.01126758, 0.0093834, 0.005175801, 0.01195924, 0.222444, 
    0.1765456, 0.09893259, 0.1201838, 0.03100987, 0.01759264,
  0.01421513, 0.004597525, 0.00175789, 0.06418556, 0.003475814, 0.007175102, 
    0.02038384, 0.01128201, 0.0137416, 0.01574021, 0.02541298, 0.02333173, 
    0.0645199, 0.09516395, 0.1201157, 0.09234756, 0.119546, 0.06833512, 
    0.1247713, 0.06493041, 0.03142579, 0.02159994, 0.08539728, 0.0776231, 
    0.02727883, 0.02662895, 0.01454569, -9.482105e-05, 0.01843118,
  4.151072e-07, 1.444019e-06, 1.262122e-06, -6.843341e-06, 1.930912e-06, 
    9.897229e-07, 1.426883e-05, -0.0001529027, 0.1424664, 0.149715, 
    0.02518125, 0.01899405, 0.03936008, 0.02983376, 0.03475303, 0.0252756, 
    0.03857737, 0.07346743, 0.008847758, 2.014677e-06, 7.350757e-07, 
    0.0381437, 0.01118457, 0.02044897, 0.02218255, 0.0370606, 0.04111334, 
    -5.19399e-05, 5.551929e-08,
  6.847655e-07, 3.971269e-05, 5.786486e-05, 4.815741e-06, 0.001280907, 
    2.108195e-06, -0.0004251991, 0.009835927, 0.2687708, 0.08573404, 
    0.09107836, 0.1698212, 0.09810649, 0.1044598, 0.0631754, 0.1014528, 
    0.0650505, 0.0406393, 0.03501366, 0.007226119, -2.327885e-06, 0.01174691, 
    0.0236002, 0.04865725, 0.06076169, 0.04713594, 0.02732296, 0.01952791, 
    -9.513178e-05,
  0.003179383, 0.01277332, 0.07645977, 0.1022707, 0.003480041, 0.002840014, 
    0.1097539, 0.005657841, 0.003367113, 0.01132799, 0.1142894, 0.09647723, 
    0.1917578, 0.1670745, 0.1721738, 0.2447047, 0.1972513, 0.1531917, 
    0.06454445, 0.1583575, 0.1164968, 0.1265625, 0.2006055, 0.1656924, 
    0.2283858, 0.171718, 0.1285392, 0.1377189, 0.0852254,
  0.1019296, 0.1693667, 0.151548, 0.1683651, 0.03064592, 0.08421286, 
    0.06922536, 0.2110336, 0.08822899, 0.05676334, 0.2698038, 0.2701739, 
    0.2394328, 0.08419553, 0.1540374, 0.2615293, 0.332498, 0.2578397, 
    0.1213449, 0.1779484, 0.1441873, 0.06353036, 0.1282207, 0.2241849, 
    0.2147389, 0.2733892, 0.2147891, 0.2751748, 0.1944069,
  0.258793, 0.269412, 0.1792294, 0.3074397, 0.2705587, 0.1748096, 0.2269278, 
    0.2791477, 0.2409719, 0.2204445, 0.1662661, 0.3047421, 0.1967996, 
    0.1564272, 0.1701412, 0.2249711, 0.3815553, 0.511143, 0.1935295, 
    0.1677858, 0.09214105, 0.08206253, 0.04737596, 0.2075427, 0.1213886, 
    0.2389066, 0.3152648, 0.2478924, 0.2610752,
  0.3117996, 0.1600135, 0.3069948, 0.1677469, 0.1906482, 0.1317093, 
    0.1380073, 0.2541087, 0.2251899, 0.1922533, 0.1752063, 0.08832522, 
    0.06439577, 0.03545571, 0.04927021, 0.1066967, 0.1353762, 0.07313062, 
    0.05063781, 0.112333, 0.1558739, 0.04054984, 0.1388451, 0.1339293, 
    0.04296568, 0.1674987, 0.1344001, 0.1835063, 0.2861029,
  0.1042245, 0.05946048, 0.07924336, 0.145268, 0.1242033, 0.1649162, 
    0.175766, 0.1767905, 0.1217952, 0.08921666, 0.06927264, 0.1586205, 
    0.2467145, 0.2680953, 0.2714671, 0.2181162, 0.1773615, 0.127512, 
    0.06199504, 0.06069528, 0.1869491, 0.1199898, 0.1454112, 0.0741569, 
    0.0503184, 0.0864728, 0.09900227, 0.133188, 0.1316731,
  0.3658895, 0.3689875, 0.3720854, 0.3751834, 0.3782814, 0.3813793, 
    0.3844773, 0.3835487, 0.3902487, 0.3969488, 0.4036488, 0.4103488, 
    0.4170489, 0.4237489, 0.4275773, 0.4302805, 0.4329838, 0.435687, 
    0.4383902, 0.4410935, 0.4437967, 0.4411659, 0.4286646, 0.4161634, 
    0.4036621, 0.3911609, 0.3786597, 0.3661585, 0.3634111,
  0.1516593, 0.2509073, 0.1227579, 0.05232412, 0.02425944, 0.04828389, 
    0.06222037, 0.01243207, 0.01363669, 0.09542697, 0.1717432, 0.2749303, 
    0.3099597, 0.2201975, 0.1601937, 0.2324197, 0.1749835, 0.09937323, 
    0.08043413, 0.1669652, 0.5882341, 0.5719039, 0.3156867, 0.1738738, 
    0.1994386, 0.1334019, 0.1180545, 0.09422206, 0.1028491,
  0.3578251, 0.4501359, 0.3475645, 0.2142105, 0.2388207, 0.0874081, 
    0.2579746, 0.396312, 0.46909, 0.399881, 0.4587604, 0.2859349, 0.1454786, 
    0.2763284, 0.3008522, 0.3355913, 0.2386192, 0.3721672, 0.5132708, 
    0.3410607, 0.447077, 0.3890856, 0.4015913, 0.3814157, 0.286072, 
    0.1695089, 0.1678638, 0.2100001, 0.4335171,
  0.384598, 0.3497989, 0.372737, 0.3292073, 0.2949869, 0.3973187, 0.4425925, 
    0.4790529, 0.4399322, 0.4615051, 0.3485719, 0.3459603, 0.3933447, 
    0.364125, 0.363466, 0.3592322, 0.3740835, 0.3608331, 0.3422553, 
    0.3539154, 0.3645677, 0.2925179, 0.3978371, 0.3700201, 0.3829805, 
    0.3008029, 0.2115024, 0.2603563, 0.4281087,
  0.3770401, 0.3261272, 0.3041377, 0.2759075, 0.2323648, 0.3032103, 
    0.2533843, 0.3840003, 0.3153708, 0.29092, 0.2991953, 0.3058972, 
    0.2484014, 0.286456, 0.1861819, 0.2126949, 0.2861177, 0.2842605, 
    0.3018016, 0.2677729, 0.2847334, 0.2415374, 0.2370617, 0.2645881, 
    0.2290383, 0.3423219, 0.3743338, 0.3557911, 0.3470343,
  0.2271953, 0.1688054, 0.1225673, 0.142327, 0.1492931, 0.1756009, 0.2235945, 
    0.2436335, 0.2200033, 0.2063949, 0.1632892, 0.1236205, 0.1627743, 
    0.2047975, 0.2346765, 0.2346212, 0.2130762, 0.2082684, 0.2377228, 
    0.2138165, 0.2359045, 0.1582288, 0.1763727, 0.2173764, 0.06605611, 
    0.2207156, 0.2492123, 0.1769526, 0.2167685,
  0.1566048, 0.04711614, 0.005385261, 0.07861097, 0.06633365, 0.08050294, 
    0.1483731, 0.1472276, 0.1928098, 0.1099411, 0.008579644, 0.0004530864, 
    0.01950136, 0.1504139, 0.08731787, 0.1685271, 0.1491838, 0.2037985, 
    0.1958251, 0.1095848, 0.1047958, 0.1614807, 0.1166145, 0.008886503, 
    0.07212247, 0.05791544, 0.131243, 0.1503771, 0.145883,
  0.1097344, 5.025603e-06, 0.00319863, 0.04882016, 0.09636935, 0.04829863, 
    0.07448856, 0.04578364, 0.07678495, 0.015727, 1.477433e-09, 
    -1.858342e-06, 0.08977975, 0.1062566, 0.05349201, 0.06839386, 0.1207271, 
    0.06530214, 0.03188239, 0.04151176, 0.07049818, 0.169895, 0.05681224, 
    0.0005851639, 0.08049165, 0.03075856, 0.04553192, 0.0977201, 0.1059175,
  7.375417e-05, 0.0005173173, 0.03427668, 0.1452882, 0.06262328, 0.04475773, 
    0.06234465, 0.03448788, 0.06177329, 0.05869043, 0.09877977, 0.0603675, 
    0.2068336, 0.02954308, 0.02949901, 0.03241765, 0.02412725, 0.04185901, 
    0.03200817, 0.02648845, 0.03421932, 0.03492964, 0.001454037, 0.04520736, 
    0.01872965, 0.006384591, 0.1035696, 0.02881014, 0.01092744,
  0.04354543, 0.1073454, 0.09735069, 0.05827074, 0.01245455, 0.01281379, 
    0.01808402, 0.01782194, 0.1258673, 0.2272645, 0.0301673, 0.01915058, 
    0.01854114, 0.01643718, 0.02151461, 0.02404105, 0.02094036, 0.01351914, 
    0.01741118, 0.01328572, 0.01334243, 0.008075756, 0.00723936, 0.1966885, 
    0.1650838, 0.08428328, 0.1002892, 0.02888142, 0.0259135,
  0.01202828, 0.003921143, 0.0007492448, 0.04153678, 0.002655936, 0.01376969, 
    0.03435577, 0.0197032, 0.02267235, 0.02227238, 0.02632569, 0.02684972, 
    0.05723091, 0.07589091, 0.08988839, 0.08212288, 0.09745996, 0.08562761, 
    0.1299503, 0.06863396, 0.04164007, 0.02274975, 0.07753275, 0.06504758, 
    0.03290671, 0.04672639, 0.0298645, -2.699959e-05, 0.01130656,
  3.30535e-07, 1.298066e-06, 8.61288e-07, -4.683007e-06, 1.303029e-06, 
    4.612656e-07, 5.035213e-06, 0.0006967203, 0.1514238, 0.1357485, 
    0.03505655, 0.02044614, 0.0385384, 0.03418903, 0.03361647, 0.03134048, 
    0.04002086, 0.06727005, 0.04720795, 0.0001636391, 3.214968e-07, 
    0.04338009, 0.01569686, 0.0185619, 0.02418424, 0.03979906, 0.1258357, 
    0.001205407, 3.831842e-08,
  2.246174e-06, 1.189168e-05, -2.180309e-05, 1.97639e-06, 0.0003338599, 
    1.310201e-06, -0.0003072672, 0.003889032, 0.2531041, 0.05960122, 
    0.1002659, 0.1672447, 0.1321886, 0.1465703, 0.113994, 0.110261, 
    0.08881115, 0.1222183, 0.09767094, 0.06465838, -1.232551e-06, 0.01868694, 
    0.01685324, 0.05006488, 0.07084911, 0.06731353, 0.05497446, 0.07192, 
    0.002136302,
  0.0009649437, 0.00691784, 0.04669308, 0.1021645, -0.00150548, 0.00194591, 
    0.09664086, 0.002854764, 0.001732809, 0.009805934, 0.1208402, 0.09408745, 
    0.2022253, 0.1934813, 0.2774097, 0.2946781, 0.2516924, 0.2384338, 
    0.1632185, 0.1429473, 0.1047321, 0.139965, 0.1471698, 0.1521143, 
    0.2527566, 0.2371935, 0.1700352, 0.1571327, 0.08674757,
  0.0865164, 0.2236724, 0.110963, 0.08807801, 0.01959386, 0.07886678, 
    0.07054302, 0.1932201, 0.06431249, 0.03980239, 0.2598782, 0.303037, 
    0.2913838, 0.09330859, 0.2961038, 0.3017806, 0.3997447, 0.3399935, 
    0.1425249, 0.1589779, 0.1390197, 0.04077357, 0.08251998, 0.196384, 
    0.2031315, 0.311068, 0.2345904, 0.3034505, 0.2154264,
  0.294817, 0.2855174, 0.1681603, 0.2759064, 0.2004951, 0.1223395, 0.20085, 
    0.2361223, 0.2243209, 0.2093055, 0.1632124, 0.2382895, 0.2305272, 
    0.1780816, 0.1954308, 0.2371474, 0.3612643, 0.5084726, 0.2401246, 
    0.2041723, 0.07091079, 0.08452808, 0.0345353, 0.2401009, 0.1397909, 
    0.2180449, 0.4485221, 0.3383938, 0.2583148,
  0.3765223, 0.2330658, 0.374809, 0.2872618, 0.1962803, 0.2292197, 0.2238703, 
    0.2256606, 0.1556439, 0.1495915, 0.1387367, 0.09419412, 0.06283436, 
    0.03251665, 0.02185203, 0.1439103, 0.126059, 0.0672866, 0.05954328, 
    0.1458435, 0.1991894, 0.03359504, 0.1637005, 0.1437981, 0.04029339, 
    0.1910473, 0.1227797, 0.2671501, 0.404762,
  0.1674273, 0.170558, 0.1463417, 0.1473974, 0.1710153, 0.1733625, 0.1638826, 
    0.1887989, 0.111613, 0.08962073, 0.07167788, 0.1543156, 0.261858, 
    0.320401, 0.3540891, 0.3119326, 0.1993857, 0.1480977, 0.08302936, 
    0.1669258, 0.1369928, 0.1316475, 0.1515418, 0.1120218, 0.08669009, 
    0.08953417, 0.07458161, 0.1605256, 0.2316472,
  0.4102564, 0.4145253, 0.4187942, 0.4230631, 0.427332, 0.4316009, 0.4358698, 
    0.3934885, 0.3993524, 0.4052162, 0.4110801, 0.416944, 0.4228078, 
    0.4286717, 0.4436453, 0.4447422, 0.4458391, 0.446936, 0.4480329, 
    0.4491298, 0.4502268, 0.4567815, 0.4455519, 0.4343222, 0.4230925, 
    0.4118628, 0.4006331, 0.3894034, 0.4068412,
  0.1815312, 0.3070099, 0.2124377, 0.06413906, 0.03501394, 0.1147765, 
    0.07277018, 0.05708095, 0.01536856, 0.1305374, 0.187021, 0.297104, 
    0.3295856, 0.1826082, 0.127429, 0.1434928, 0.1480094, 0.0644626, 
    0.07103977, 0.1613222, 0.599491, 0.5845106, 0.359441, 0.1252703, 
    0.2017566, 0.1352722, 0.1143429, 0.1075297, 0.1171603,
  0.3786405, 0.4358296, 0.3807952, 0.1888353, 0.2454467, 0.1192411, 
    0.2420426, 0.4159935, 0.4542102, 0.4198997, 0.4462915, 0.259718, 
    0.1561533, 0.291171, 0.3053184, 0.2841656, 0.3592549, 0.4886366, 
    0.5043494, 0.3947059, 0.4584332, 0.4372689, 0.3965821, 0.3772353, 
    0.2727997, 0.1536526, 0.2024222, 0.2730936, 0.4142127,
  0.2936313, 0.3371158, 0.3389827, 0.3361426, 0.312163, 0.3936537, 0.4789932, 
    0.4387653, 0.3537566, 0.4985967, 0.427305, 0.3410729, 0.3823938, 
    0.3998894, 0.3691946, 0.353508, 0.3548364, 0.3425254, 0.3265828, 
    0.3185181, 0.3520287, 0.3153875, 0.3791392, 0.3625494, 0.4128022, 
    0.3335582, 0.2799574, 0.34498, 0.4460401,
  0.3856568, 0.2993212, 0.3044122, 0.2930427, 0.2701972, 0.3337225, 
    0.2830777, 0.3246734, 0.2810876, 0.2691912, 0.247159, 0.2838986, 
    0.3024301, 0.2982828, 0.2050739, 0.2546416, 0.2695303, 0.3012905, 
    0.268081, 0.2947907, 0.2725683, 0.2720229, 0.2817739, 0.252486, 
    0.1867509, 0.4061108, 0.484702, 0.4330896, 0.3158284,
  0.270465, 0.2806962, 0.1593625, 0.2025309, 0.2046342, 0.1917366, 0.2914124, 
    0.3104788, 0.2276826, 0.1409389, 0.1717158, 0.101838, 0.156624, 
    0.1609226, 0.2614584, 0.2005799, 0.2058211, 0.2368107, 0.2391462, 
    0.2133343, 0.2271513, 0.17151, 0.1894686, 0.2573759, 0.07774414, 
    0.1908358, 0.2040565, 0.1717587, 0.2642734,
  0.1512524, 0.04496279, 0.007539972, 0.08912909, 0.09599225, 0.08869923, 
    0.1412804, 0.1459781, 0.2259789, 0.1278538, 0.0006538633, 4.266573e-05, 
    0.01322214, 0.08772183, 0.08876397, 0.1201734, 0.104239, 0.1911385, 
    0.2099718, 0.08242856, 0.1224289, 0.170772, 0.2152067, 0.0116765, 
    0.07182388, 0.08617213, 0.1041207, 0.07886998, 0.1700294,
  0.07514365, -1.810302e-05, 0.001220974, 0.05324063, 0.1098964, 0.06335183, 
    0.0686061, 0.07995309, 0.07967193, 0.009735825, 9.371318e-10, 
    2.163489e-07, 0.1014666, 0.126139, 0.06466402, 0.08380756, 0.1141194, 
    0.1208328, 0.06228524, 0.06449185, 0.06697969, 0.1709563, 0.3481245, 
    0.00074783, 0.09139315, 0.02751946, 0.08023132, 0.1314355, 0.1260284,
  0.001570813, 0.0005207143, 0.02544479, 0.155734, 0.06135665, 0.05063142, 
    0.06551787, 0.03814198, 0.07005971, 0.08765136, 0.1078795, 0.1106204, 
    0.1948446, 0.03213366, 0.042415, 0.0404967, 0.04240323, 0.04195278, 
    0.04984761, 0.05562761, 0.0426313, 0.1090475, 0.03271919, 0.0405737, 
    0.02575534, 0.001192999, 0.102788, 0.08222017, 0.1234502,
  0.05304328, 0.08642869, 0.07999379, 0.03741904, 0.02645171, 0.02429927, 
    0.02667636, 0.0384415, 0.1131426, 0.2006042, 0.03444643, 0.02379419, 
    0.03015486, 0.02554495, 0.04586862, 0.03903926, 0.02836503, 0.01569787, 
    0.01980419, 0.01925468, 0.0186157, 0.02013621, 0.006975483, 0.1600772, 
    0.1356554, 0.07701159, 0.08606828, 0.03102081, 0.03454409,
  0.009218211, 0.002404459, 0.0002988068, 0.02459437, 0.002094339, 
    0.03730555, 0.04548194, 0.03220751, 0.01447093, 0.03839802, 0.0411888, 
    0.03374989, 0.05555103, 0.06707123, 0.07433288, 0.07689253, 0.08555648, 
    0.09202768, 0.1458949, 0.07982231, 0.05549552, 0.06507012, 0.07762528, 
    0.07101551, 0.03820343, 0.06137626, 0.07546303, 0.0006845155, 0.006864072,
  2.780038e-07, 1.152086e-06, 5.619834e-07, -1.001763e-06, 1.020043e-06, 
    2.648923e-07, -1.256225e-07, 0.002494839, 0.1440474, 0.128096, 
    0.07092132, 0.02634813, 0.06717058, 0.04104874, 0.04404486, 0.06715862, 
    0.04947535, 0.07348504, 0.2430792, 0.02656584, 2.075773e-08, 0.04366918, 
    0.01915404, 0.02244551, 0.0497165, 0.06535211, 0.1539564, 0.0525031, 
    2.910325e-08,
  1.264145e-06, 6.243826e-06, -0.0001637445, 1.541653e-06, 6.195704e-05, 
    8.686703e-07, -0.0002407059, 0.0006187533, 0.2524133, 0.04827197, 
    0.1452967, 0.2125636, 0.1924731, 0.1737634, 0.2244473, 0.1585756, 
    0.1992825, 0.1932083, 0.3602808, 0.1473003, -5.462347e-06, 0.03057021, 
    0.04322157, 0.07724784, 0.08448754, 0.09503189, 0.103537, 0.2046627, 
    0.002669855,
  0.001069777, 0.003864081, 0.0399639, 0.100786, -0.001511924, 0.0005148472, 
    0.09574617, 0.002436598, 0.001112783, 0.01015292, 0.1339656, 0.09091791, 
    0.197993, 0.2431193, 0.3262906, 0.3429217, 0.296324, 0.3669647, 
    0.2617304, 0.1274055, 0.09894886, 0.2369674, 0.1418635, 0.1577891, 
    0.2829866, 0.3204657, 0.2363988, 0.2146465, 0.119021,
  0.1082947, 0.154552, 0.09806477, 0.05216946, 0.02870146, 0.05405245, 
    0.06717937, 0.18513, 0.04638433, 0.0295862, 0.2352314, 0.3014856, 
    0.3108337, 0.2425941, 0.4310516, 0.4273516, 0.4422388, 0.3947687, 
    0.2271758, 0.1595093, 0.1226568, 0.04880549, 0.05689178, 0.1862082, 
    0.1988784, 0.3982046, 0.235804, 0.2816181, 0.2089682,
  0.2195344, 0.2606163, 0.1103819, 0.2464695, 0.1609249, 0.1086245, 
    0.1706795, 0.2038602, 0.1906347, 0.1851663, 0.163917, 0.2260506, 
    0.2217705, 0.1915992, 0.2504462, 0.3944507, 0.3763184, 0.5228803, 
    0.2218712, 0.1696282, 0.05076484, 0.08039055, 0.07969485, 0.2881899, 
    0.1597467, 0.2264031, 0.5440406, 0.4007128, 0.2927196,
  0.5072591, 0.3175387, 0.3897179, 0.3784933, 0.3571909, 0.2551556, 
    0.1224304, 0.1886702, 0.1296909, 0.1512599, 0.1014045, 0.09845763, 
    0.03760955, 0.03149537, 0.05722574, 0.248308, 0.1145575, 0.08402097, 
    0.06264078, 0.1226832, 0.1973436, 0.07577451, 0.1446869, 0.1800961, 
    0.153689, 0.2414517, 0.1241134, 0.3723131, 0.6174492,
  0.2067223, 0.2164584, 0.1819392, 0.2227379, 0.2117433, 0.2564303, 0.198363, 
    0.1789732, 0.2222669, 0.1724263, 0.2008182, 0.1797115, 0.3397751, 
    0.4019881, 0.3835946, 0.3483218, 0.2716649, 0.1766972, 0.1676088, 
    0.2155637, 0.1815875, 0.1723884, 0.1334032, 0.261101, 0.1347569, 
    0.1160614, 0.082012, 0.2401027, 0.2871497,
  0.4384012, 0.4430297, 0.4476582, 0.4522866, 0.4569151, 0.4615435, 0.466172, 
    0.4143759, 0.4202605, 0.4261451, 0.4320297, 0.4379143, 0.443799, 
    0.4496836, 0.4590657, 0.4565721, 0.4540784, 0.4515848, 0.4490911, 
    0.4465975, 0.4441038, 0.4564127, 0.4483932, 0.4403738, 0.4323544, 
    0.4243349, 0.4163155, 0.4082961, 0.4346984,
  0.2070991, 0.3335978, 0.2577789, 0.090419, 0.04840971, 0.1684358, 0.108021, 
    0.06254244, 0.0160684, 0.1469968, 0.2202599, 0.319783, 0.3533949, 
    0.1236386, 0.1313651, 0.1446501, 0.1459885, 0.05107095, 0.06718339, 
    0.1819562, 0.6418731, 0.6247611, 0.3591562, 0.1460915, 0.2176787, 
    0.1347399, 0.1543213, 0.1316068, 0.1886202,
  0.3849415, 0.3879499, 0.3651227, 0.1723977, 0.2283957, 0.1175729, 
    0.2114676, 0.4365023, 0.4512847, 0.4404771, 0.4195229, 0.2290962, 
    0.1686898, 0.2835536, 0.3137324, 0.2995464, 0.4737716, 0.5198853, 
    0.4039297, 0.3925095, 0.4765498, 0.5210032, 0.4102612, 0.3940819, 
    0.2982877, 0.1487441, 0.2185943, 0.3258285, 0.3816748,
  0.2535053, 0.2780024, 0.2734782, 0.3240876, 0.3354486, 0.390305, 0.4813549, 
    0.3455161, 0.300264, 0.4377804, 0.3994159, 0.3338198, 0.4114965, 
    0.3865837, 0.345707, 0.3578816, 0.3351542, 0.3146096, 0.2829847, 
    0.3092855, 0.3362835, 0.314966, 0.3713599, 0.3756725, 0.4700442, 
    0.4660946, 0.3615226, 0.3954551, 0.3459186,
  0.4297257, 0.389544, 0.3691764, 0.3320192, 0.3021176, 0.3047995, 0.2999375, 
    0.2897104, 0.2673211, 0.2422764, 0.2497, 0.2745912, 0.2717873, 0.2857803, 
    0.2574599, 0.2705987, 0.2650603, 0.29366, 0.2375563, 0.250809, 0.2681, 
    0.2600388, 0.2671672, 0.2751379, 0.1742402, 0.4358656, 0.3798465, 
    0.4419283, 0.3588446,
  0.3328204, 0.2606442, 0.1293111, 0.1881156, 0.1936599, 0.2018561, 
    0.3102618, 0.2306246, 0.1562103, 0.1319063, 0.1601318, 0.1022266, 
    0.1063476, 0.1009569, 0.2922109, 0.1408149, 0.179629, 0.2503178, 
    0.1924007, 0.2047973, 0.1798702, 0.1765048, 0.1710161, 0.2891715, 
    0.08208199, 0.1382899, 0.1732645, 0.1300062, 0.2611144,
  0.1783934, 0.07405662, 0.008823313, 0.06533574, 0.07571604, 0.1096883, 
    0.08823472, 0.1115414, 0.1955526, 0.04212079, -3.038347e-05, 
    -2.441885e-05, 0.009364204, 0.05297277, 0.09993643, 0.1180283, 
    0.06172785, 0.1593608, 0.1909836, 0.05768691, 0.08531513, 0.1082863, 
    0.1668744, 0.01548057, 0.07161311, 0.06340419, 0.05662567, 0.04543299, 
    0.09212328,
  0.3671913, -3.718736e-05, 0.0007293187, 0.04313591, 0.1284354, 0.06582336, 
    0.08801997, 0.09167483, 0.07415353, 0.03742055, 8.457542e-10, 
    8.720605e-08, 0.06387673, 0.1605151, 0.08044591, 0.05785743, 0.08632073, 
    0.08566832, 0.07623494, 0.04666485, 0.04322185, 0.08833872, 0.3455537, 
    -0.000646441, 0.1202388, 0.0153449, 0.05040896, 0.09424407, 0.1599304,
  0.1805998, 0.0002987396, 0.007767458, 0.1195802, 0.08198484, 0.09725022, 
    0.09510121, 0.05162318, 0.06301412, 0.04496915, 0.05674752, 0.07507779, 
    0.1828773, 0.05844403, 0.04572859, 0.07697952, 0.05156478, 0.06119455, 
    0.05381386, 0.04413923, 0.03643677, 0.1264642, 0.2539994, 0.04413415, 
    0.007465579, 0.0002757853, 0.09463046, 0.09867968, 0.3193894,
  0.08328731, 0.05373174, 0.06408419, 0.02973324, 0.2645345, 0.1616885, 
    0.1485244, 0.1111768, 0.07222933, 0.164732, 0.09684017, 0.0614224, 
    0.03256725, 0.1708796, 0.05084775, 0.05136792, 0.06415673, 0.0402621, 
    0.05008866, 0.03411351, 0.03196882, 0.06026387, 0.00937205, 0.1275634, 
    0.09065733, 0.07664108, 0.1142219, 0.1265524, 0.05923942,
  0.00561043, 0.001335636, 7.293616e-05, 0.01683194, 0.01006069, 0.1340733, 
    0.06172644, 0.154171, 0.02707692, 0.2621556, 0.09124825, 0.1438356, 
    0.07939602, 0.09064638, 0.0840582, 0.07527452, 0.0924574, 0.127028, 
    0.1408982, 0.1558936, 0.1561558, 0.09266127, 0.06840705, 0.05354875, 
    0.04803928, 0.1065261, 0.1652866, 0.01064405, 0.00323826,
  2.517205e-07, 1.044057e-06, 4.268027e-07, 6.405563e-06, 9.225481e-07, 
    -6.806734e-07, -2.587418e-06, 0.01692806, 0.1234539, 0.1289994, 
    0.08901392, 0.06113808, 0.08415717, 0.07790718, 0.06974651, 0.07087777, 
    0.03354774, 0.04501536, 0.2689831, 0.3146057, -1.750559e-06, 0.04206586, 
    0.0571646, 0.04068615, 0.06091131, 0.06882311, 0.06808674, 0.1210191, 
    2.208986e-08,
  9.977374e-07, 4.595572e-06, -0.0002896556, 1.567771e-06, -2.038956e-05, 
    6.464228e-07, -0.0001737431, 0.002332166, 0.2580658, 0.04813316, 
    0.1485441, 0.2949875, 0.2105789, 0.2069583, 0.1746334, 0.1795804, 
    0.2340894, 0.2154558, 0.4498286, 0.1944124, -1.440681e-05, 0.03321107, 
    0.03620594, 0.1405085, 0.1476637, 0.1853485, 0.214006, 0.3435919, 
    0.007903122,
  0.002675696, 0.002451167, 0.03254949, 0.1045914, 0.005938393, 0.0002803331, 
    0.09979986, 0.003727949, 0.0006507965, 0.009671037, 0.1498697, 0.0850062, 
    0.2518451, 0.379714, 0.3997986, 0.3768789, 0.3761941, 0.4427993, 
    0.2461571, 0.121567, 0.0875215, 0.2578462, 0.1451364, 0.1693667, 
    0.302591, 0.3273033, 0.2974263, 0.2745294, 0.1447649,
  0.1149417, 0.1136034, 0.0829142, 0.0363679, 0.02400283, 0.03960593, 
    0.07090836, 0.1694911, 0.03328882, 0.02400939, 0.2154355, 0.3133644, 
    0.3195571, 0.4589223, 0.4047404, 0.4047101, 0.473037, 0.4055209, 
    0.2960533, 0.128824, 0.1156394, 0.04734189, 0.04207942, 0.1877688, 
    0.1903539, 0.5237657, 0.2630841, 0.2987239, 0.2532636,
  0.1684526, 0.2003542, 0.09098397, 0.2187922, 0.1345573, 0.1017397, 
    0.1459078, 0.1900288, 0.1737549, 0.1565986, 0.140875, 0.2060535, 
    0.2083322, 0.1842109, 0.3171198, 0.4550242, 0.3748819, 0.5276288, 
    0.2137048, 0.1366203, 0.05393329, 0.08896419, 0.2156717, 0.3131038, 
    0.2435046, 0.2087342, 0.5665413, 0.3749738, 0.3439942,
  0.4686298, 0.2831442, 0.3363791, 0.2362234, 0.3544052, 0.1853645, 
    0.06399335, 0.1681534, 0.09375317, 0.1204404, 0.09824225, 0.09196834, 
    0.04002599, 0.026205, 0.1244668, 0.409528, 0.1526636, 0.07224427, 
    0.07838217, 0.09033264, 0.1735892, 0.08393688, 0.1429399, 0.2866035, 
    0.2687025, 0.2593098, 0.1215386, 0.3273806, 0.6050363,
  0.3655011, 0.2575891, 0.2557642, 0.2846488, 0.3212608, 0.2324274, 
    0.2094542, 0.2085463, 0.2394096, 0.265743, 0.218881, 0.2510707, 
    0.3850789, 0.474674, 0.4437079, 0.3457943, 0.3259876, 0.2831137, 
    0.2956325, 0.2375024, 0.2228003, 0.2263417, 0.174555, 0.3028723, 
    0.2092933, 0.1945087, 0.1423746, 0.3370647, 0.294479,
  0.4339935, 0.4381829, 0.4423721, 0.4465615, 0.4507508, 0.4549401, 
    0.4591294, 0.4178836, 0.4243389, 0.4307942, 0.4372496, 0.4437049, 
    0.4501603, 0.4566156, 0.4544036, 0.4501111, 0.4458185, 0.441526, 
    0.4372334, 0.4329409, 0.4286483, 0.4559607, 0.4496086, 0.4432565, 
    0.4369044, 0.4305523, 0.4242002, 0.4178481, 0.4306421,
  0.2452309, 0.3665509, 0.2969489, 0.1050328, 0.05696812, 0.1840162, 
    0.1352746, 0.06149384, 0.009832429, 0.1544529, 0.2196326, 0.322246, 
    0.4471426, 0.07869685, 0.1429196, 0.1635182, 0.2123651, 0.05460689, 
    0.06364612, 0.2138962, 0.6695626, 0.6480166, 0.3623843, 0.1344524, 
    0.1727303, 0.1357799, 0.1448471, 0.1538845, 0.2196674,
  0.3544871, 0.3245151, 0.3034615, 0.1394382, 0.1769487, 0.1071998, 
    0.1668133, 0.4545942, 0.4476739, 0.4348499, 0.4174682, 0.210616, 
    0.1674535, 0.2616486, 0.2969936, 0.3318889, 0.4559021, 0.4503923, 
    0.2883731, 0.3924555, 0.5004369, 0.5339798, 0.4410254, 0.3959019, 
    0.3521386, 0.1916623, 0.2424966, 0.4012958, 0.3790728,
  0.2224432, 0.2283089, 0.2518579, 0.3347622, 0.3719033, 0.4154622, 
    0.4282689, 0.2694283, 0.2477241, 0.3569356, 0.3483258, 0.3532409, 
    0.4125233, 0.3663205, 0.354454, 0.381092, 0.341777, 0.3101631, 0.2441542, 
    0.2909599, 0.3074921, 0.3300566, 0.3831324, 0.3455574, 0.5434937, 
    0.5616822, 0.4102809, 0.3465571, 0.2443842,
  0.4076779, 0.3867918, 0.4404356, 0.382791, 0.3294747, 0.3156455, 0.2950125, 
    0.261495, 0.2567184, 0.2137419, 0.2554226, 0.2691404, 0.2417952, 
    0.2362685, 0.2387916, 0.2065988, 0.2430668, 0.252024, 0.2020442, 
    0.2182826, 0.2430888, 0.2167314, 0.2137957, 0.3045077, 0.1721755, 
    0.3773195, 0.3281096, 0.3620747, 0.3735179,
  0.2638228, 0.1773031, 0.08467457, 0.1246698, 0.2055106, 0.216159, 
    0.3079577, 0.214563, 0.1626291, 0.1035276, 0.1362234, 0.08233404, 
    0.0524142, 0.1000732, 0.345187, 0.1244765, 0.1361488, 0.1553612, 
    0.1428727, 0.2115311, 0.2063936, 0.155709, 0.1313467, 0.3301331, 
    0.06103915, 0.1243336, 0.1127689, 0.09673055, 0.2338799,
  0.08242799, 0.07898533, 0.006565363, 0.04312624, 0.03321388, 0.06610839, 
    0.08673975, 0.04802642, 0.1499557, 0.0220649, 2.472597e-05, -3.90648e-05, 
    0.007004356, 0.02283689, 0.05807133, 0.08902102, 0.04944856, 0.1318638, 
    0.1702048, 0.05359408, 0.03985502, 0.05014726, 0.07087939, 0.02081552, 
    0.04720268, 0.03065815, 0.03950024, 0.0173746, 0.04245182,
  0.2363444, 0.0001681701, 0.001669817, 0.05486058, 0.06123659, 0.0489586, 
    0.03063129, 0.032973, 0.06039569, 0.005829087, 9.487693e-10, 
    4.470731e-08, 0.02189383, 0.07423741, 0.03823838, 0.04313948, 0.1466262, 
    0.05465464, 0.02543995, 0.01216934, 0.01755692, 0.03177887, 0.1209911, 
    0.02536913, 0.1171099, 0.0122404, 0.01897685, 0.02797505, 0.1154497,
  0.3340344, 0.0003084198, 0.002932837, 0.07942684, 0.0626215, 0.02913306, 
    0.05013361, 0.03037682, 0.04249103, 0.007601214, 0.02925731, 0.01671661, 
    0.1539655, 0.080405, 0.02845736, 0.02131949, 0.02720916, 0.03366604, 
    0.02960389, 0.01238939, 0.009969804, 0.0315829, 0.4214161, 0.02493876, 
    0.001384301, 5.665189e-05, 0.04942723, 0.01854068, 0.1266166,
  0.1493215, 0.03043483, 0.05478672, 0.02494141, 0.0484413, 0.03172017, 
    0.04345584, 0.02247969, 0.04051998, 0.1041694, 0.05043671, 0.1376133, 
    0.01640238, 0.02574392, 0.01714419, 0.03028131, 0.05268881, 0.07435739, 
    0.06314277, 0.0610089, 0.08204292, 0.1909797, 0.06410718, 0.0948067, 
    0.05856673, 0.07289445, 0.08022341, 0.1425794, 0.2337148,
  0.002458826, 0.0007847449, -3.27454e-05, 0.01047366, 0.007066306, 
    0.03252429, 0.06146864, 0.0248961, 0.003129469, 0.04413025, 0.03504647, 
    0.04932433, 0.04951252, 0.06051468, 0.06755754, 0.06159428, 0.06299461, 
    0.0715395, 0.0967706, 0.08919124, 0.1057288, 0.07422397, 0.1351925, 
    0.04084248, 0.01967133, 0.0313221, 0.09424494, 0.3507681, 0.001407086,
  2.428851e-07, 9.589568e-07, 3.702755e-07, 5.867512e-05, 8.605954e-07, 
    -0.000391572, -4.118811e-05, 0.03939389, 0.08382808, 0.1595761, 
    0.1063576, 0.1455002, 0.0336986, 0.02475344, 0.02827528, 0.01366637, 
    0.01315761, 0.008610402, 0.08499238, 0.5356069, 0.01180165, 0.04060704, 
    0.01403669, 0.02676626, 0.05202071, 0.01608633, 0.01129903, 0.1085991, 
    1.787896e-08,
  9.35272e-07, -1.320091e-05, -8.573863e-05, 1.565818e-06, -3.833454e-05, 
    5.242961e-07, -0.0001428994, 0.004300157, 0.2786853, 0.04941817, 
    0.1914606, 0.2433512, 0.286588, 0.194005, 0.1469609, 0.1913141, 
    0.2086035, 0.09914207, 0.246475, 0.1773401, -7.309312e-06, 0.02521786, 
    0.02829347, 0.1912142, 0.1653382, 0.1826058, 0.1946776, 0.1400882, 
    0.005024101,
  0.007857283, 0.004289452, 0.02830162, 0.1027475, 0.01451536, -1.406765e-05, 
    0.09794199, 0.0040885, 0.0002903549, 0.008891574, 0.1583777, 0.1115922, 
    0.2760486, 0.3809776, 0.4302306, 0.3565937, 0.4137959, 0.4055412, 
    0.3209982, 0.1241624, 0.08052608, 0.1969883, 0.1329937, 0.1852976, 
    0.2575929, 0.321531, 0.3091279, 0.2213062, 0.1293776,
  0.09725791, 0.1042734, 0.07737325, 0.03145942, 0.02282291, 0.03445952, 
    0.06540412, 0.1459261, 0.02545765, 0.02174329, 0.2192207, 0.3143516, 
    0.3566742, 0.3950859, 0.2846638, 0.3298354, 0.4332233, 0.3808718, 
    0.302727, 0.1103175, 0.113954, 0.04256821, 0.03822669, 0.1699124, 
    0.2107809, 0.4873285, 0.2643666, 0.2864948, 0.2769445,
  0.1444674, 0.1789479, 0.08300791, 0.1914507, 0.1107425, 0.09442408, 
    0.1360041, 0.181753, 0.1727037, 0.1555568, 0.1251921, 0.1668357, 
    0.1847048, 0.1695525, 0.2654731, 0.4878361, 0.3762927, 0.5133263, 
    0.2233783, 0.1219073, 0.06377047, 0.1175139, 0.2379547, 0.3151075, 
    0.2326604, 0.2005875, 0.5143278, 0.3149433, 0.3662257,
  0.3803077, 0.2085235, 0.2696148, 0.09311689, 0.2296546, 0.1824532, 
    0.08200444, 0.1477103, 0.05586223, 0.1152058, 0.09567436, 0.06968278, 
    0.03115398, 0.03948009, 0.226728, 0.5825467, 0.2161558, 0.0811996, 
    0.05965266, 0.08918044, 0.1618584, 0.11817, 0.1215455, 0.3696305, 
    0.3005912, 0.232194, 0.1331965, 0.2214223, 0.5625818,
  0.4056242, 0.2559476, 0.3668705, 0.2855704, 0.405775, 0.2969833, 0.2376844, 
    0.2418053, 0.2265657, 0.2672934, 0.3040848, 0.3928955, 0.4556228, 
    0.5479511, 0.5492071, 0.3941844, 0.435089, 0.3621542, 0.3369318, 
    0.2568164, 0.2208873, 0.2779042, 0.1392726, 0.2353898, 0.1609853, 
    0.1556129, 0.13169, 0.2887351, 0.2925901,
  0.3853813, 0.3901182, 0.394855, 0.3995918, 0.4043287, 0.4090655, 0.4138023, 
    0.3708212, 0.3792619, 0.3877027, 0.3961434, 0.4045841, 0.4130249, 
    0.4214656, 0.4560623, 0.4506646, 0.445267, 0.4398693, 0.4344717, 
    0.429074, 0.4236763, 0.4308228, 0.4230429, 0.415263, 0.407483, 0.3997031, 
    0.3919232, 0.3841433, 0.3815919,
  0.2860303, 0.365562, 0.2857846, 0.1090773, 0.04794043, 0.1730224, 
    0.1313513, 0.0667918, 0.009426826, 0.1215926, 0.2174812, 0.2979626, 
    0.4810877, 0.04129631, 0.1649699, 0.2440844, 0.2526227, 0.06423635, 
    0.06915077, 0.2242202, 0.6878245, 0.6721112, 0.3424037, 0.0903864, 
    0.126004, 0.1544142, 0.1631807, 0.1956778, 0.2484832,
  0.3123604, 0.2529864, 0.2571186, 0.1014131, 0.1249141, 0.09140746, 
    0.1223198, 0.4343849, 0.4621917, 0.4249337, 0.4201273, 0.2274926, 
    0.1649274, 0.2181373, 0.2763266, 0.3604457, 0.4618286, 0.3466057, 
    0.2050218, 0.4015612, 0.5255373, 0.5526772, 0.4782319, 0.3894301, 
    0.3662826, 0.2213084, 0.2898442, 0.3924813, 0.3615663,
  0.1780193, 0.193367, 0.2343769, 0.3585246, 0.3567455, 0.3967131, 0.3576969, 
    0.205608, 0.1965207, 0.2777498, 0.3158512, 0.3342503, 0.4011756, 
    0.395107, 0.3500755, 0.3743983, 0.3395522, 0.2993505, 0.2141115, 
    0.2654697, 0.2826082, 0.2841082, 0.3610636, 0.3273849, 0.5370166, 
    0.6313936, 0.4924172, 0.2408017, 0.1795515,
  0.3499472, 0.3818897, 0.4104744, 0.3881889, 0.3433022, 0.3424587, 
    0.2925839, 0.2436532, 0.2413829, 0.1968851, 0.2381793, 0.2747484, 
    0.2170877, 0.1736258, 0.1831416, 0.213986, 0.2323427, 0.2183638, 
    0.1654505, 0.1845284, 0.2125299, 0.1965563, 0.1885362, 0.2974998, 
    0.1519752, 0.3236946, 0.297798, 0.3042606, 0.3454888,
  0.2412546, 0.1179991, 0.06496316, 0.0830039, 0.1795239, 0.174613, 
    0.2211642, 0.1844385, 0.1436397, 0.0715033, 0.09668991, 0.0400694, 
    0.01500824, 0.09263363, 0.364283, 0.1022162, 0.09858796, 0.110921, 
    0.1090447, 0.2052535, 0.1801251, 0.1243007, 0.109895, 0.3494503, 
    0.03430353, 0.1141548, 0.08569995, 0.08437409, 0.2335258,
  0.02943716, 0.03009978, 0.00534627, 0.02864849, 0.01436018, 0.03503062, 
    0.0363051, 0.02253732, 0.0814814, 0.0131398, 2.029161e-05, -3.620456e-05, 
    0.003332854, 0.006089109, 0.04818261, 0.07560851, 0.03784536, 0.1016292, 
    0.162382, 0.08593591, 0.0484789, 0.01953542, 0.03274832, 0.03343501, 
    0.04136258, 0.01460894, 0.04723332, 0.01148431, 0.01389865,
  0.09178349, 0.00403792, 0.0004727559, 0.006829378, 0.03144345, 0.02315872, 
    0.01142612, 0.007615114, 0.06686568, 0.001635124, 1.263238e-09, 
    2.476483e-08, 0.006466587, 0.03539058, 0.01333106, 0.01725316, 
    0.04779425, 0.02282516, 0.005860875, 0.0009898437, 0.00186052, 
    0.008069754, 0.03780738, 0.02996079, 0.08693077, 0.01408902, 0.002368655, 
    0.00793861, 0.04091286,
  0.1716135, 0.0002121345, 0.001042421, 0.06194873, 0.0213637, 0.007881154, 
    0.02163513, 0.00731063, 0.0129645, 0.001403692, 0.01523735, 0.001937695, 
    0.14047, 0.02061745, 0.007371688, 0.00472817, 0.006097736, 0.02027461, 
    0.01222062, 0.00187034, 0.001082979, 0.006900527, 0.1559356, 0.008029024, 
    0.0003137164, 9.615504e-06, 0.01763209, 0.004221625, 0.04253396,
  0.06390513, 0.02761705, 0.04355657, 0.02027416, 0.009540818, 0.005580401, 
    0.007076877, 0.003525371, 0.03651785, 0.06605638, 0.01415146, 0.02554245, 
    0.001680561, 0.004939791, 0.001574048, 0.003857251, 0.007446626, 
    0.01620191, 0.01836577, 0.03001111, 0.05174918, 0.1206516, 0.3967993, 
    0.081546, 0.04045469, 0.05841026, 0.07040082, 0.0309681, 0.0937712,
  0.001101589, 0.0005489873, -3.688049e-05, 0.00506265, 0.004046817, 
    0.006195709, 0.0361551, 0.005561276, 5.736081e-06, 0.009397152, 
    0.006844611, 0.01327917, 0.01914053, 0.03107642, 0.04084633, 0.04139746, 
    0.03011892, 0.02962703, 0.04276064, 0.0347191, 0.02859941, 0.01602686, 
    0.1927449, 0.03597475, 0.002071462, 0.00899887, 0.0294924, 0.2079806, 
    -0.0003247511,
  2.370659e-07, 8.870317e-07, 3.468301e-07, 0.00315784, 8.171677e-07, 
    0.001141422, -0.0001303843, 0.03703759, 0.05237813, 0.1815854, 
    0.04741554, 0.02195192, 0.004746841, 0.00401648, 0.00917655, 0.002110874, 
    0.002917027, 0.001073977, 0.02968585, 0.237235, 0.003895444, 0.03688657, 
    0.00219042, 0.01171116, 0.009215607, 0.001732159, 0.002354677, 
    0.02602168, 1.597047e-08,
  9.023854e-07, -8.202226e-05, -4.373019e-05, 1.291521e-06, -4.537782e-05, 
    4.617573e-07, -0.0001341697, 0.00521593, 0.2945915, 0.03911463, 
    0.1751875, 0.2582572, 0.2863948, 0.1964472, 0.2367224, 0.1580068, 
    0.1280973, 0.0234774, 0.1140143, 0.1106853, -1.759253e-06, 0.03756625, 
    0.04679357, 0.1152826, 0.08611531, 0.07350098, 0.06772771, 0.04283242, 
    0.01009015,
  0.01061853, 0.002604549, 0.01908744, 0.1134715, 0.01780683, -2.115787e-06, 
    0.09009428, 0.003776985, 0.0001845052, 0.007429245, 0.168058, 0.1351134, 
    0.276994, 0.3182833, 0.3541362, 0.3099501, 0.3364818, 0.366011, 
    0.2323515, 0.1192727, 0.0681928, 0.1546489, 0.1278728, 0.1932371, 
    0.2301794, 0.29371, 0.2504066, 0.1570443, 0.1029879,
  0.08383651, 0.1164026, 0.06508175, 0.03503713, 0.01914496, 0.03327756, 
    0.0540878, 0.1210293, 0.01820048, 0.01942658, 0.2069411, 0.3010462, 
    0.3732454, 0.2540753, 0.166214, 0.2580612, 0.3762912, 0.3574741, 
    0.2405929, 0.09826148, 0.09016337, 0.03810172, 0.03154742, 0.1470869, 
    0.17734, 0.4423328, 0.2212543, 0.2710717, 0.3011143,
  0.1457615, 0.1597232, 0.07676566, 0.1731785, 0.08878258, 0.08203843, 
    0.1230373, 0.1556311, 0.1629445, 0.1503289, 0.1156766, 0.1369658, 
    0.160961, 0.1173806, 0.1737387, 0.5633661, 0.3437856, 0.509174, 
    0.2049755, 0.1068775, 0.06344063, 0.08270667, 0.1818579, 0.3121656, 
    0.318848, 0.1915517, 0.3745642, 0.2603475, 0.346258,
  0.3630903, 0.159841, 0.2325432, 0.04565562, 0.1430656, 0.2572638, 
    0.09915292, 0.08827762, 0.03378029, 0.1022822, 0.08289511, 0.0555477, 
    0.03670201, 0.08808706, 0.2312054, 0.5852671, 0.2617172, 0.09176124, 
    0.06424102, 0.09453952, 0.2003894, 0.09033968, 0.1149108, 0.3459098, 
    0.2559564, 0.1807098, 0.1409137, 0.1522045, 0.5230691,
  0.2824006, 0.2020348, 0.284912, 0.2860066, 0.447071, 0.3981566, 0.3292318, 
    0.3136186, 0.3006996, 0.2880749, 0.3038669, 0.419844, 0.4783727, 
    0.5631391, 0.6088851, 0.4681771, 0.4273601, 0.4165919, 0.2660033, 
    0.2482121, 0.2865126, 0.3044928, 0.1372833, 0.1889276, 0.1197919, 
    0.129329, 0.1230678, 0.2546602, 0.2131758,
  0.2851419, 0.2876454, 0.2901489, 0.2926524, 0.2951559, 0.2976593, 
    0.3001629, 0.2642801, 0.2733125, 0.2823449, 0.2913774, 0.3004098, 
    0.3094422, 0.3184746, 0.3759879, 0.3735506, 0.3711133, 0.368676, 
    0.3662388, 0.3638015, 0.3613642, 0.3455783, 0.3364796, 0.327381, 
    0.3182823, 0.3091837, 0.300085, 0.2909864, 0.2831391,
  0.3023286, 0.3388455, 0.2285225, 0.09194328, 0.04447735, 0.13489, 
    0.1136703, 0.06064174, 0.003868844, 0.05426341, 0.1835727, 0.2726294, 
    0.5095472, 0.01403929, 0.2170537, 0.3277678, 0.3322854, 0.07832265, 
    0.07906473, 0.2579488, 0.6913624, 0.6814758, 0.295541, 0.06989575, 
    0.107579, 0.1765536, 0.2125632, 0.2083135, 0.2785164,
  0.2753304, 0.185952, 0.2228425, 0.07557475, 0.09838104, 0.07765427, 
    0.08937319, 0.4075386, 0.4562003, 0.4059867, 0.4088637, 0.2449198, 
    0.1539322, 0.1687814, 0.2837679, 0.4051055, 0.4446906, 0.2735014, 
    0.1376871, 0.3917834, 0.504499, 0.5792207, 0.4652055, 0.3948413, 
    0.365146, 0.2946151, 0.3760649, 0.3716251, 0.344181,
  0.1466995, 0.1595842, 0.2091328, 0.3049849, 0.2832891, 0.3434416, 
    0.2994609, 0.1526395, 0.1597804, 0.2196813, 0.272899, 0.2923645, 
    0.3495276, 0.3971769, 0.3308384, 0.3501311, 0.3164994, 0.2652723, 
    0.1773911, 0.2361217, 0.2622247, 0.2252022, 0.3270463, 0.2923557, 
    0.5077398, 0.6266709, 0.5477241, 0.1758207, 0.1342941,
  0.2992108, 0.3911341, 0.3604296, 0.3655807, 0.3468952, 0.3627947, 
    0.2764201, 0.2108874, 0.2209075, 0.1771333, 0.2098726, 0.2490438, 
    0.1923718, 0.1321438, 0.1569947, 0.2025336, 0.1993394, 0.1822233, 
    0.1357254, 0.1601775, 0.1690041, 0.1625187, 0.1595456, 0.2563438, 
    0.13957, 0.2843844, 0.2641026, 0.2615916, 0.2860997,
  0.2013235, 0.08452138, 0.05054041, 0.0505326, 0.1647963, 0.1341353, 
    0.1502143, 0.1282405, 0.09737261, 0.04530467, 0.06206818, 0.01803673, 
    0.00569055, 0.05825179, 0.3405928, 0.07528733, 0.0800062, 0.0872456, 
    0.09260561, 0.1765408, 0.154011, 0.09384092, 0.09331281, 0.3393243, 
    0.021164, 0.09962557, 0.06716719, 0.07797643, 0.2204779,
  0.0127066, 0.008455426, 0.003770658, 0.01544942, 0.004711784, 0.02279824, 
    0.01874967, 0.01379693, 0.04124696, 0.008731585, -2.272333e-07, 
    -3.692667e-05, 0.001032618, 0.002452009, 0.03177366, 0.06044085, 
    0.02929349, 0.07032092, 0.1332818, 0.05309949, 0.02623663, 0.00856877, 
    0.01544391, 0.04590402, 0.03171435, 0.005219243, 0.01805107, 0.006822979, 
    0.005149138,
  0.03489866, 0.007683563, 2.131064e-06, 0.002390898, 0.0134566, 0.009731956, 
    0.002338164, 0.001738907, 0.04034117, 0.0007297699, 1.619336e-09, 
    2.114693e-08, 0.002004773, 0.01903391, 0.005506731, 0.003878433, 
    0.01904209, 0.006105592, 0.001626013, 0.0002906531, 0.0003053996, 
    0.001667498, 0.01550173, 0.04309144, 0.05912253, 0.02716905, 
    0.0009738208, 0.002322531, 0.01318408,
  0.08160808, 0.0007926305, 0.0002308436, 0.05522599, 0.006960947, 
    0.00127112, 0.007134729, 0.0008127094, 0.004756312, 0.0001454701, 
    0.00651491, 0.0006203596, 0.1031634, 0.003391882, 0.002614646, 
    0.0005192168, 0.001340437, 0.01360093, 0.006584607, 0.0006350387, 
    0.0003991352, 0.0027044, 0.06507289, 0.002470147, 0.0001047683, 
    3.534717e-06, 0.008824917, 0.001713601, 0.01745484,
  0.0114406, 0.02611543, 0.04211048, 0.02090504, 0.003771833, 0.001998596, 
    0.002190508, 0.001297346, 0.03621079, 0.05243974, 0.002591318, 
    0.007720911, 0.0002258336, 0.001902129, 0.0001828507, 0.0005236731, 
    0.001673305, 0.003575332, 0.002166893, 0.003154387, 0.01155353, 
    0.03042437, 0.3053831, 0.07984857, 0.03564284, 0.05395185, 0.03657685, 
    0.006049541, 0.01879152,
  0.000347749, 0.0002497751, -2.899186e-05, 0.004879121, 0.002064192, 
    0.002270342, 0.0124077, 0.002142005, -5.431197e-05, 0.004079604, 
    0.001140723, 0.003934377, 0.004831993, 0.01073876, 0.01492191, 
    0.01918416, 0.01516398, 0.01306429, 0.01728634, 0.0115541, 0.008940696, 
    0.004805195, 0.1547692, 0.03832309, 5.937305e-05, 0.002636121, 
    0.01102063, 0.07935669, -0.00115573,
  2.271413e-07, 8.403388e-07, 3.369851e-07, 0.004050099, 7.99018e-07, 
    6.376056e-05, -0.000132247, 0.0152149, 0.03563502, 0.0927469, 0.01050148, 
    0.00659166, 0.001026112, 0.001062776, 0.00111857, 0.0008363614, 
    0.000447974, 9.645968e-05, 0.01379935, 0.1172277, 0.001706756, 
    0.02772511, 0.0009370795, -0.0001486724, 0.003006259, 0.0005370785, 
    0.0009137788, 0.01194759, 1.492094e-08,
  8.855823e-07, -0.000188324, -1.286221e-05, 9.035662e-07, -6.788217e-05, 
    4.276382e-07, -0.0001289863, 0.005727567, 0.3073771, 0.02341546, 
    0.1553635, 0.2446949, 0.2382983, 0.1757542, 0.1937499, 0.1422693, 
    0.07340798, 0.009185741, 0.05439317, 0.06301007, -6.785687e-07, 
    0.04685709, 0.03584488, 0.07118148, 0.04030953, 0.03528121, 0.02629412, 
    0.01675721, 0.008622495,
  0.009267236, 0.003837507, 0.01107207, 0.1263102, 0.008280487, 8.91685e-07, 
    0.08251007, 0.002239951, 8.891174e-05, 0.005921626, 0.1663472, 0.1134668, 
    0.2858272, 0.2961242, 0.2677696, 0.2513686, 0.2581837, 0.340193, 
    0.1423785, 0.1125058, 0.05703574, 0.1397939, 0.1051281, 0.1753348, 
    0.1727852, 0.233311, 0.1864134, 0.1110794, 0.09790684,
  0.06526856, 0.1201438, 0.05490343, 0.03224695, 0.01436104, 0.02554481, 
    0.04265609, 0.09971894, 0.01357767, 0.01564812, 0.1896009, 0.2724389, 
    0.4440382, 0.1780362, 0.09761036, 0.2108751, 0.3183015, 0.3073474, 
    0.1888254, 0.08869992, 0.07104839, 0.02887147, 0.02441415, 0.1226186, 
    0.1636666, 0.4093913, 0.1670263, 0.2440349, 0.3046442,
  0.1650588, 0.1504295, 0.07004623, 0.146541, 0.07452695, 0.07432076, 
    0.1094343, 0.1323599, 0.1428961, 0.1428838, 0.111464, 0.08683632, 
    0.1283493, 0.07541534, 0.1070106, 0.5561872, 0.2942567, 0.4300878, 
    0.1770367, 0.09486513, 0.049644, 0.05229388, 0.1048169, 0.259791, 
    0.2711632, 0.1779436, 0.2971086, 0.2421805, 0.3232015,
  0.3643444, 0.1280827, 0.2022448, 0.0268529, 0.09284986, 0.2617, 0.09288007, 
    0.03591628, 0.02028179, 0.09008158, 0.08377596, 0.05589582, 0.02147302, 
    0.1421089, 0.2524064, 0.5031952, 0.3337005, 0.08621802, 0.05735851, 
    0.1008174, 0.180048, 0.09882767, 0.09087345, 0.3564781, 0.219015, 
    0.1236793, 0.1321521, 0.1201115, 0.5262609,
  0.1991001, 0.1395603, 0.2256895, 0.2858401, 0.3457645, 0.329752, 0.3659478, 
    0.3379112, 0.2672216, 0.3241835, 0.3189661, 0.4004164, 0.5054736, 
    0.5478305, 0.5714173, 0.4854736, 0.4383653, 0.427557, 0.2315675, 
    0.2768194, 0.3048467, 0.2721214, 0.1882809, 0.1358823, 0.1029901, 
    0.0974534, 0.0927225, 0.2314513, 0.1587506,
  0.2236998, 0.2233455, 0.2229912, 0.222637, 0.2222827, 0.2219284, 0.2215741, 
    0.1796542, 0.1921897, 0.2047252, 0.2172607, 0.2297962, 0.2423318, 
    0.2548673, 0.3380937, 0.3357836, 0.3334734, 0.3311633, 0.3288532, 
    0.3265431, 0.324233, 0.269086, 0.2592149, 0.2493438, 0.2394727, 
    0.2296015, 0.2197304, 0.2098593, 0.2239832,
  0.3218701, 0.2817795, 0.1335417, 0.05776772, 0.03801143, 0.07651259, 
    0.05052511, 0.04858177, 0.002766277, 0.01718576, 0.1087566, 0.264251, 
    0.5066445, 0.002603155, 0.3197264, 0.3937566, 0.4931969, 0.1583188, 
    0.07687608, 0.2909162, 0.6926274, 0.7111261, 0.2646719, 0.05818103, 
    0.1234991, 0.2240198, 0.2365674, 0.1915946, 0.3002182,
  0.2430674, 0.1488363, 0.1794609, 0.0499017, 0.09115095, 0.07311146, 
    0.05944632, 0.367376, 0.4384135, 0.3790184, 0.3912472, 0.2477724, 
    0.1345117, 0.1284344, 0.3059495, 0.3892798, 0.4226245, 0.2138039, 
    0.09605918, 0.3324485, 0.4495677, 0.5128634, 0.4277811, 0.3996252, 
    0.3598483, 0.3314609, 0.4563174, 0.344292, 0.2966309,
  0.1056226, 0.1272935, 0.1743841, 0.2343461, 0.2158895, 0.2698056, 
    0.2451126, 0.1149871, 0.1268246, 0.1677421, 0.2350962, 0.2500619, 
    0.301148, 0.3493551, 0.2546507, 0.28104, 0.2585034, 0.2182243, 0.1426038, 
    0.2037733, 0.2266231, 0.1597615, 0.2648229, 0.2484706, 0.4621207, 
    0.5755507, 0.4657215, 0.1332875, 0.09971169,
  0.2621436, 0.3576995, 0.3102936, 0.3308237, 0.3428495, 0.3203278, 
    0.2373689, 0.1737737, 0.18973, 0.1398791, 0.1617222, 0.1746137, 
    0.1412087, 0.09561601, 0.1363335, 0.1647777, 0.1618617, 0.1269386, 
    0.09839166, 0.1362203, 0.1245055, 0.1204976, 0.1198029, 0.2131294, 
    0.1256762, 0.2416464, 0.2095147, 0.2092882, 0.2363982,
  0.1437885, 0.05677748, 0.02583457, 0.02943445, 0.1196416, 0.08293079, 
    0.09439593, 0.08541059, 0.05858081, 0.02920323, 0.04226463, 0.01066605, 
    0.002938128, 0.03178363, 0.2926719, 0.05632469, 0.06217831, 0.073768, 
    0.07721489, 0.133508, 0.1226923, 0.0614801, 0.06182242, 0.3081831, 
    0.01375185, 0.07628501, 0.05128644, 0.05497933, 0.1948658,
  0.006446648, 0.003902951, 0.002427634, 0.006512812, 0.001678943, 
    0.01382178, 0.01321397, 0.008316241, 0.02272944, 0.006127802, 
    1.121536e-06, -7.685931e-06, 0.001382893, 0.001154041, 0.01589389, 
    0.04026488, 0.01951564, 0.04128531, 0.09332272, 0.02438468, 0.01369184, 
    0.003806994, 0.006592113, 0.03946365, 0.02294645, 0.001993123, 
    0.007466719, 0.003317789, 0.002527474,
  0.01957875, 0.005456572, -5.279628e-05, 0.001235473, 0.005534925, 
    0.004829166, 0.00099508, 0.0007627293, 0.01594924, 0.0004205982, 
    1.610348e-09, 1.655961e-08, 0.000880159, 0.009957592, 0.002001565, 
    0.001137467, 0.007227654, 0.002063982, 0.0007025098, 0.0001658879, 
    0.000112393, 0.0008543115, 0.008365133, 0.03230658, 0.03880245, 
    0.04336666, 0.000571319, 0.001243178, 0.00693763,
  0.04419643, 0.0001712152, -2.959583e-05, 0.03306968, 0.002140159, 
    0.0006535113, 0.002946527, 0.0001196505, 0.001541115, -0.00017876, 
    0.003217236, 0.0003375301, 0.05974269, 0.0009269932, 0.0008496365, 
    0.0001597866, 0.0005304562, 0.006736023, 0.002092232, 0.0002119144, 
    0.0002032196, 0.001432911, 0.03449629, 0.001940589, 6.243172e-05, 
    2.347829e-06, 0.00274396, 0.0009235058, 0.00967741,
  0.004402154, 0.03096976, 0.04874497, 0.0158091, 0.002031623, 0.00110314, 
    0.001116983, 0.0007133916, 0.02677713, 0.07396123, 0.0009332985, 
    0.00418498, 0.0001177599, 0.001027407, 8.064696e-05, 0.000259185, 
    0.0008062631, 0.001693716, 0.0007333106, 0.0007796132, 0.002838064, 
    0.01115449, 0.1356447, 0.07962979, 0.03737505, 0.03691573, 0.02038164, 
    0.002730345, 0.006813355,
  0.000129147, 0.000118556, -2.048614e-05, 0.005999994, 0.001937064, 
    0.001270761, 0.003246679, 0.001218117, 2.367666e-06, 0.002338699, 
    0.0004996178, 0.001974813, 0.001317486, 0.003328279, 0.003984845, 
    0.00602681, 0.007629887, 0.007549788, 0.003977518, 0.004832749, 
    0.004627493, 0.002404866, 0.1178142, 0.03997925, 2.712675e-05, 
    0.001132551, 0.004294555, 0.04194258, -0.001634002,
  2.189581e-07, 8.10418e-07, 3.322008e-07, 0.002741734, 7.857533e-07, 
    8.136922e-08, -9.086695e-05, 0.001990015, 0.02750543, 0.04610385, 
    0.004479406, 0.003152171, 0.0004760243, 0.0004850255, 0.0004816759, 
    0.0004954532, 0.0001277353, 2.803184e-05, 0.008250435, 0.07119559, 
    0.001021765, 0.0223295, 0.0005402176, -0.0006822616, 0.001547016, 
    0.0002939911, 0.0005018123, 0.006978573, 1.415776e-08,
  8.816457e-07, -0.0001695161, -3.047412e-06, 5.654657e-07, -7.371025e-05, 
    4.087032e-07, -0.0001324957, 0.005482828, 0.2987669, 0.01555305, 
    0.1517693, 0.1727439, 0.1820107, 0.1090168, 0.1004534, 0.08108523, 
    0.04691282, 0.005432867, 0.03161125, 0.03607392, -3.337958e-07, 
    0.04368327, 0.01783395, 0.03145706, 0.0206095, 0.0161781, 0.01480864, 
    0.009644989, 0.008210404,
  0.006663489, 0.001903435, 0.00622878, 0.1295401, 0.00383899, 1.022174e-06, 
    0.06925035, 0.001309491, 4.201458e-05, 0.005270202, 0.1604019, 0.1004168, 
    0.2656631, 0.2641362, 0.2128198, 0.2090367, 0.2089122, 0.3073347, 
    0.08938069, 0.1043285, 0.04578569, 0.1185175, 0.08244523, 0.1453418, 
    0.116575, 0.1736683, 0.1159129, 0.06013392, 0.08536325,
  0.04325598, 0.1015728, 0.03937341, 0.02315457, 0.010216, 0.01813758, 
    0.03179676, 0.08006009, 0.00935299, 0.01648176, 0.1745986, 0.2436961, 
    0.4340209, 0.1181661, 0.05879503, 0.1659589, 0.2569779, 0.2508994, 
    0.1555624, 0.07432854, 0.05369638, 0.0202096, 0.01866038, 0.1021993, 
    0.1468149, 0.3768243, 0.1124439, 0.1817074, 0.2602886,
  0.1832607, 0.1343918, 0.06293275, 0.1256803, 0.06215139, 0.06339017, 
    0.09947786, 0.1074883, 0.120115, 0.1277973, 0.1025882, 0.05920396, 
    0.1026561, 0.05386594, 0.06840835, 0.4780252, 0.2492059, 0.3349437, 
    0.1359163, 0.08391555, 0.03342645, 0.03485915, 0.08282328, 0.2202023, 
    0.1979603, 0.1566756, 0.2620753, 0.2012884, 0.2690619,
  0.3319059, 0.09962419, 0.1709276, 0.01914128, 0.0723597, 0.2239254, 
    0.07749166, 0.01716706, 0.01114338, 0.08201993, 0.07503895, 0.0496787, 
    0.04539651, 0.1271116, 0.2771769, 0.4111869, 0.3786433, 0.1012922, 
    0.06733625, 0.1022417, 0.1614871, 0.2151777, 0.07568351, 0.3187171, 
    0.2050492, 0.07821111, 0.1273835, 0.09830603, 0.5036988,
  0.1404479, 0.09790557, 0.1344803, 0.2359096, 0.2544562, 0.260512, 
    0.3354387, 0.2845236, 0.241283, 0.3095272, 0.3176177, 0.3841507, 
    0.4486449, 0.4922847, 0.5281994, 0.4545854, 0.3937937, 0.4109274, 
    0.2499442, 0.3143778, 0.2658269, 0.2269424, 0.1759902, 0.1016938, 
    0.08798245, 0.07224357, 0.07131135, 0.1856382, 0.1251528,
  0.1599583, 0.156792, 0.1536257, 0.1504595, 0.1472932, 0.1441269, 0.1409607, 
    0.1097276, 0.1238201, 0.1379127, 0.1520053, 0.1660978, 0.1801904, 
    0.194283, 0.2652265, 0.2658286, 0.2664306, 0.2670327, 0.2676347, 
    0.2682367, 0.2688388, 0.2331404, 0.2216121, 0.2100837, 0.1985554, 
    0.187027, 0.1754987, 0.1639703, 0.1624913,
  0.3757266, 0.2360641, 0.05164206, 0.01969273, 8.071572e-06, 0.03214131, 
    0.004549421, -0.0001014838, 0.02620312, 0.02640208, 0.07583938, 
    0.2407866, 0.4375501, -0.001350056, 0.3658754, 0.4494294, 0.5424489, 
    0.183112, 0.06805417, 0.3483344, 0.6986187, 0.7603091, 0.231124, 
    0.04390514, 0.124176, 0.2632831, 0.2880972, 0.1708416, 0.3093643,
  0.1992507, 0.1253505, 0.147197, 0.03475864, 0.0849314, 0.06923636, 
    0.04263158, 0.330023, 0.4035926, 0.3507943, 0.3681757, 0.2671973, 
    0.1095979, 0.102338, 0.2918929, 0.3418169, 0.3882598, 0.1676094, 
    0.06809865, 0.2963366, 0.3903537, 0.4359918, 0.3635997, 0.366957, 
    0.3345623, 0.360963, 0.4737811, 0.290753, 0.2719727,
  0.07597123, 0.09999871, 0.1356868, 0.1819322, 0.1659321, 0.2071963, 
    0.1881306, 0.08241527, 0.09745201, 0.1247961, 0.1865816, 0.1940892, 
    0.2544586, 0.2721439, 0.1950908, 0.2112208, 0.1988428, 0.1689933, 
    0.1151275, 0.1660558, 0.1777259, 0.1084711, 0.1983405, 0.2050858, 
    0.3929928, 0.5045494, 0.3831435, 0.1041761, 0.0732904,
  0.2133211, 0.293946, 0.2442149, 0.2809034, 0.3026184, 0.2659915, 0.2017553, 
    0.1358045, 0.1507831, 0.09968606, 0.1109479, 0.1116283, 0.08321349, 
    0.06187252, 0.1036592, 0.117135, 0.1221356, 0.08843447, 0.06546158, 
    0.1027517, 0.09290852, 0.08267639, 0.07729314, 0.1816185, 0.1028094, 
    0.1913411, 0.161771, 0.1578394, 0.1930053,
  0.09777394, 0.03814035, 0.01335554, 0.01826653, 0.07591912, 0.04691238, 
    0.05627166, 0.0531486, 0.03189942, 0.02012072, 0.02487621, 0.005510709, 
    0.001886541, 0.01608203, 0.2470717, 0.03676543, 0.04147114, 0.05458411, 
    0.05230538, 0.08746205, 0.09107392, 0.0373529, 0.03414761, 0.2819014, 
    0.008282644, 0.05226382, 0.03097633, 0.03324859, 0.1437713,
  0.00426787, 0.00250038, 0.005003713, 0.003027775, 0.0009560328, 
    0.005464192, 0.009315963, 0.004697922, 0.01047379, 0.004056591, 
    -1.142361e-05, -1.019707e-05, 0.001658401, 0.0007803814, 0.007095396, 
    0.02167055, 0.01059929, 0.01914911, 0.05334643, 0.01064399, 0.004560267, 
    0.002207016, 0.003553813, 0.02588602, 0.01513908, 0.001031448, 
    0.004412735, 0.001460108, 0.001604109,
  0.01309754, 0.004036564, -4.837972e-05, 0.00080141, 0.001666271, 
    0.002146903, 0.0006591083, 0.0004700803, 0.005391202, 0.0002931476, 
    -5.192407e-09, 1.361179e-08, 0.0006262168, 0.004123865, 0.0005734778, 
    0.000641409, 0.003559269, 0.0009730573, 0.0004131414, 0.0001125882, 
    6.20139e-05, 0.0005673765, 0.005485931, 0.02693081, 0.02585856, 
    0.04580515, 0.0003897681, 0.0008363599, 0.004639852,
  0.02812258, 4.366684e-05, -1.353481e-05, 0.01727966, 0.0008684325, 
    0.000436224, 0.001235316, 5.87109e-05, 0.0007804381, -0.0001739563, 
    0.001788098, 0.0002083004, 0.03247232, 0.0004819267, 0.00029248, 
    0.0001257295, 0.0002668536, 0.002852445, 0.0007056777, 0.0001049651, 
    0.0001247793, 0.0009155373, 0.02200141, 0.001869168, 0.0006293138, 
    1.445486e-06, 0.0005056037, 0.0005902021, 0.006394125,
  0.002609601, 0.02932206, 0.04890946, 0.01075033, 0.001299976, 0.0007192781, 
    0.0006921963, 0.0004647656, 0.02450157, 0.08673001, 0.0005618723, 
    0.002755024, 7.755709e-05, 0.0006541493, 4.824252e-05, 0.0001629837, 
    0.0005111299, 0.001024636, 0.0004072367, 0.0004314274, 0.001529318, 
    0.00640631, 0.07830907, 0.06946225, 0.03445637, 0.01819188, 0.009673162, 
    0.001709069, 0.003931846,
  6.185631e-05, 6.850099e-05, -1.341028e-05, 0.006659422, 0.0009167417, 
    0.0008437434, 0.0006597842, 0.000804558, 1.041673e-05, 0.001557101, 
    0.0003153098, 0.001293858, 0.0004841827, 0.001119477, 0.001099821, 
    0.002051624, 0.003611662, 0.003417189, 0.001058111, 0.002289584, 
    0.003112878, 0.00121527, 0.08663449, 0.04104239, 1.515627e-05, 
    0.000682409, 0.002326349, 0.02638026, -0.0008944828,
  2.109423e-07, 7.903659e-07, 3.295646e-07, 0.001475273, 7.761794e-07, 
    -1.3765e-06, -5.608168e-05, 0.0008189903, 0.02777839, 0.0208787, 
    0.002742165, 0.001974563, 0.0003064974, 0.0003019626, 0.0002995142, 
    0.0003375308, 6.923365e-05, 1.356612e-05, 0.00573092, 0.049741, 
    0.0007169366, 0.01725944, 0.0003615721, -0.0006194602, 0.0009998321, 
    0.0001920598, 0.0003310951, 0.004700931, 1.407352e-08,
  8.817613e-07, -7.23726e-05, -2.078298e-06, 6.723294e-08, -3.996936e-05, 
    3.926055e-07, -0.0001351278, 0.00551035, 0.2814927, 0.01076708, 
    0.1312781, 0.1062583, 0.1148203, 0.05855054, 0.07790433, 0.0380506, 
    0.02704069, 0.003787328, 0.02174969, 0.02478639, -1.722092e-07, 
    0.0357466, 0.01049893, 0.01413381, 0.01117506, 0.007641439, 0.0103568, 
    0.006689331, 0.008035469,
  0.004619498, 0.001249014, 0.003631326, 0.1160912, 0.001455182, 
    9.975552e-07, 0.05846968, 0.0009380649, 2.098112e-05, 0.004878341, 
    0.1471534, 0.09056395, 0.2294838, 0.2275159, 0.1704179, 0.1619669, 
    0.1507993, 0.246513, 0.05645773, 0.09257015, 0.03635172, 0.1002861, 
    0.06523681, 0.1155728, 0.07278305, 0.1129258, 0.06062346, 0.0284677, 
    0.06209734,
  0.04294065, 0.08221857, 0.02777627, 0.01597943, 0.007705322, 0.01316661, 
    0.02327447, 0.06630295, 0.006975504, 0.0148714, 0.1545127, 0.2184637, 
    0.3788959, 0.08283456, 0.04332866, 0.1335484, 0.1894735, 0.1989234, 
    0.1129249, 0.06164977, 0.0366783, 0.01440557, 0.01352562, 0.08698949, 
    0.1370343, 0.3306814, 0.06924406, 0.1223083, 0.191312,
  0.1477194, 0.1136779, 0.05196105, 0.0998716, 0.05118874, 0.05330057, 
    0.08760057, 0.08600685, 0.09838685, 0.1062988, 0.08936255, 0.04482149, 
    0.07917199, 0.04057062, 0.0462616, 0.3517165, 0.203699, 0.2595874, 
    0.09857079, 0.07424358, 0.02297475, 0.02585986, 0.09760578, 0.1739938, 
    0.1550815, 0.1246907, 0.1896028, 0.1280593, 0.2020011,
  0.2895123, 0.07261168, 0.1438916, 0.01545563, 0.05103374, 0.1539494, 
    0.07332444, 0.01245249, 0.009380063, 0.07257312, 0.07326383, 0.04819987, 
    0.07174603, 0.1148112, 0.2358609, 0.2875691, 0.3536474, 0.09294832, 
    0.07379454, 0.09465759, 0.1809196, 0.2745744, 0.06855402, 0.2767865, 
    0.1807691, 0.05767552, 0.1140632, 0.07993931, 0.4359086,
  0.1122337, 0.09643249, 0.1044284, 0.1833997, 0.1900677, 0.1944751, 
    0.2600592, 0.2291117, 0.2358803, 0.2817927, 0.2928586, 0.3331766, 
    0.340963, 0.3909777, 0.4436547, 0.3849201, 0.3343893, 0.3455529, 
    0.2540784, 0.2997889, 0.251229, 0.1735394, 0.1462983, 0.09418167, 
    0.06861039, 0.05274925, 0.05607148, 0.1659507, 0.09200612,
  0.1298458, 0.1275699, 0.125294, 0.1230181, 0.1207423, 0.1184664, 0.1161905, 
    0.09684664, 0.1070957, 0.1173448, 0.1275939, 0.1378429, 0.148092, 
    0.1583411, 0.1883202, 0.1891809, 0.1900417, 0.1909024, 0.1917631, 
    0.1926239, 0.1934846, 0.1832568, 0.1744229, 0.165589, 0.1567551, 
    0.1479212, 0.1390873, 0.1302533, 0.1316665,
  0.4501016, 0.1901356, 0.04221844, 0.003741551, 0.001572451, 0.00750882, 
    0.00596017, 0.001993569, 0.0001326191, 0.02003828, 0.05529343, 0.2172111, 
    0.3797147, -0.003253396, 0.3927169, 0.4767308, 0.5878987, 0.2158434, 
    0.06599796, 0.3988501, 0.7005682, 0.818873, 0.2242158, 0.03841154, 
    0.140116, 0.2835388, 0.3145162, 0.1542275, 0.3240189,
  0.1751154, 0.1089839, 0.1398291, 0.03009016, 0.0770539, 0.06593312, 
    0.03488743, 0.2851362, 0.3710999, 0.3259119, 0.3797706, 0.2945379, 
    0.09478977, 0.08850059, 0.2972188, 0.3075845, 0.3506303, 0.1343184, 
    0.05413575, 0.2700202, 0.346357, 0.382533, 0.3244562, 0.3245956, 
    0.2980686, 0.3442816, 0.4342013, 0.2485782, 0.2549367,
  0.06142992, 0.08226186, 0.1068202, 0.1496234, 0.1366829, 0.1671575, 
    0.1519317, 0.06449989, 0.07756785, 0.1015469, 0.1504428, 0.1510066, 
    0.2138735, 0.2152101, 0.1536192, 0.1660815, 0.1597195, 0.13946, 
    0.09543712, 0.1338231, 0.1419436, 0.08198972, 0.1532896, 0.1611479, 
    0.3336791, 0.4192776, 0.3186031, 0.08735955, 0.05654716,
  0.1736649, 0.2476125, 0.2025002, 0.234811, 0.2654417, 0.2183046, 0.1707753, 
    0.1084242, 0.1240589, 0.07639185, 0.07956672, 0.08144607, 0.05576551, 
    0.04167605, 0.07541087, 0.0852677, 0.08860103, 0.06326137, 0.04507205, 
    0.07775225, 0.07144684, 0.05969552, 0.05315609, 0.1667065, 0.07732463, 
    0.1417289, 0.1282805, 0.126009, 0.1623573,
  0.06524689, 0.02465837, 0.00847696, 0.01263742, 0.04809478, 0.02748469, 
    0.0348398, 0.03639947, 0.01741202, 0.0138973, 0.0133783, 0.002783367, 
    0.001442335, 0.009060706, 0.2171031, 0.02142756, 0.02665985, 0.03793932, 
    0.03509126, 0.05559039, 0.06422029, 0.02335188, 0.02173477, 0.2532252, 
    0.006499548, 0.03317068, 0.01774251, 0.02008869, 0.0998814,
  0.003144836, 0.001866415, 0.006158669, 0.001619333, 0.000710926, 
    0.00277016, 0.005229148, 0.003072943, 0.006284789, 0.002579811, 
    -0.000123632, -6.763747e-06, 0.002725184, 0.0006192328, 0.003951053, 
    0.01090344, 0.004954112, 0.01007172, 0.03017257, 0.005526857, 
    0.002177382, 0.001530221, 0.002590854, 0.01902243, 0.0130138, 
    0.0006613384, 0.003258328, 0.0007659834, 0.001163315,
  0.009887439, 0.003205813, -3.749125e-05, 0.0005879954, 6.27313e-05, 
    0.001057224, 0.0005020593, 0.0003401678, 0.002817088, 0.0002257341, 
    -1.677342e-07, 1.18194e-08, 0.0004946538, 0.001902192, 0.0002848202, 
    0.0004543575, 0.002100915, 0.0006090709, 0.0002946465, 8.651941e-05, 
    4.136129e-05, 0.000428113, 0.004093534, 0.0229885, 0.02061445, 
    0.04206672, 0.0002951878, 0.0006332488, 0.003471782,
  0.02039213, 4.447426e-06, 0.0002923622, 0.01330338, 0.0005722728, 
    0.0003288983, 0.0007031093, 3.850019e-05, 0.000413373, -0.000151258, 
    0.001146841, 0.0001520975, 0.01760923, 0.0002796915, 0.000191483, 
    0.0001028389, 0.0001757478, 0.001265948, 0.0004097601, 6.791593e-05, 
    8.865103e-05, 0.0006684447, 0.01600122, 0.003604906, 0.002220142, 
    3.073055e-06, 3.814752e-05, 0.0004307619, 0.004781053,
  0.00171942, 0.02809139, 0.03678098, 0.007131091, 0.0009396888, 
    0.0005257276, 0.0004899832, 0.0003375613, 0.02057269, 0.08133366, 
    0.0003854644, 0.002029652, 5.836298e-05, 0.0004697308, 3.403015e-05, 
    0.0001192402, 0.0003727486, 0.0007230557, 0.0002751768, 0.000298424, 
    0.001040028, 0.004430695, 0.05196194, 0.05241948, 0.02960987, 0.00837539, 
    0.004591846, 0.001240371, 0.002732675,
  4.77782e-05, 1.863015e-05, -7.569256e-06, 0.006898197, 0.0005036927, 
    0.0006208565, -0.0005645193, 0.0005859671, 4.118736e-08, 0.00115914, 
    0.0002288435, 0.0009581366, 0.0002649486, 0.000557213, 0.0004285114, 
    0.0007400958, 0.001722497, 0.001680053, 0.0005116157, 0.001379125, 
    0.002372258, 0.0008015328, 0.07808616, 0.03870444, 1.03109e-05, 
    0.0004841115, 0.001561352, 0.01912436, -0.0005378634,
  2.033635e-07, 7.779288e-07, 3.276972e-07, 0.001007643, 7.667069e-07, 
    -1.385188e-06, -3.483595e-05, 0.0005633415, 0.03646442, 0.01078794, 
    0.001986622, 0.001417658, 0.0002279093, 0.0002173555, 0.0002186271, 
    0.0002562323, 4.655341e-05, 9.050447e-06, 0.00443967, 0.03844832, 
    0.0005556704, 0.01381789, 0.0002708707, -0.0008480726, 0.0007332431, 
    0.0001427213, 0.0002483994, 0.003547079, 1.394014e-08,
  8.823856e-07, -4.279372e-05, -1.426925e-06, 4.300488e-07, -2.345504e-05, 
    3.821649e-07, -0.0001338828, 0.005187079, 0.2659992, 0.008299121, 
    0.1183069, 0.06266674, 0.06889372, 0.03611191, 0.05863427, 0.02290396, 
    0.01563733, 0.002949754, 0.01678875, 0.01911987, -7.783618e-08, 
    0.03050556, 0.01148356, 0.0083553, 0.006232912, 0.004405636, 0.008072243, 
    0.005204481, 0.006359056,
  0.003279773, 0.0002269898, 0.002385771, 0.1071477, 0.0006742689, 
    9.741497e-07, 0.04897751, 0.0007437818, 1.086886e-05, 0.004479812, 
    0.1350473, 0.07534112, 0.1837661, 0.1884137, 0.1325334, 0.123858, 
    0.1085731, 0.1768838, 0.03693365, 0.08228777, 0.03038565, 0.08484314, 
    0.05134044, 0.09171322, 0.04849067, 0.07223717, 0.03414695, 0.01467893, 
    0.042976,
  0.05169709, 0.06766944, 0.02017995, 0.01154141, 0.005950202, 0.01039791, 
    0.01811491, 0.05739613, 0.005925813, 0.01365331, 0.1336614, 0.1949769, 
    0.2882476, 0.06823695, 0.04149118, 0.1091983, 0.1474988, 0.1471821, 
    0.08172788, 0.05553209, 0.02835599, 0.01142658, 0.01105015, 0.07860254, 
    0.1251491, 0.2664159, 0.04481979, 0.07876261, 0.1322044,
  0.1157649, 0.09164577, 0.04566716, 0.08074689, 0.04508371, 0.04486249, 
    0.08313368, 0.07323331, 0.08741487, 0.09251196, 0.0783233, 0.04735408, 
    0.07408672, 0.0355753, 0.0362727, 0.2612292, 0.1724624, 0.2122401, 
    0.1014566, 0.06449469, 0.0177191, 0.02477229, 0.09618445, 0.1487769, 
    0.1230334, 0.1033218, 0.1311461, 0.07880118, 0.1434634,
  0.2170868, 0.05173146, 0.1253148, 0.0133362, 0.03977225, 0.1046398, 
    0.08320764, 0.01459463, 0.0144389, 0.0653553, 0.07160429, 0.04967058, 
    0.1151575, 0.1140159, 0.1932855, 0.2242699, 0.3404692, 0.08300229, 
    0.08105184, 0.1170439, 0.1830359, 0.2893897, 0.08916031, 0.2591182, 
    0.1790049, 0.05000546, 0.1238351, 0.07297238, 0.3583075,
  0.1103508, 0.1168626, 0.08235699, 0.140119, 0.1386837, 0.1446992, 
    0.1889526, 0.1720703, 0.1988627, 0.2305793, 0.2491111, 0.2622458, 
    0.2608078, 0.316266, 0.3515013, 0.3005782, 0.277997, 0.2852958, 
    0.2142128, 0.2666549, 0.2481597, 0.1403183, 0.126357, 0.0849287, 
    0.0565095, 0.04309114, 0.04336843, 0.1564074, 0.0844741,
  0.1142291, 0.1111387, 0.1080483, 0.1049578, 0.1018674, 0.09877702, 
    0.09568661, 0.09896562, 0.1095164, 0.1200671, 0.1306179, 0.1411686, 
    0.1517194, 0.1622701, 0.1760827, 0.1776361, 0.1791895, 0.1807429, 
    0.1822963, 0.1838497, 0.1854031, 0.1792216, 0.1702078, 0.1611941, 
    0.1521803, 0.1431666, 0.1341529, 0.1251391, 0.1167014,
  0.3889688, 0.1094372, 0.02380452, 0.003926403, 0.0008987734, 0.005293367, 
    0.005082765, 0.001534852, 9.771952e-05, 0.01677429, 0.05299937, 
    0.1867943, 0.3654442, -0.003872392, 0.4205222, 0.4805417, 0.5778924, 
    0.2758497, 0.07923865, 0.4391133, 0.6649759, 0.835078, 0.2481565, 
    0.04615059, 0.1403892, 0.2800215, 0.3466277, 0.1632668, 0.3144901,
  0.1668466, 0.1042618, 0.1297714, 0.03340607, 0.1075668, 0.06110083, 
    0.03179587, 0.2693032, 0.3620613, 0.3222315, 0.3680567, 0.3086273, 
    0.08873668, 0.08058225, 0.3058838, 0.2870069, 0.3344603, 0.1178759, 
    0.04661036, 0.2520925, 0.3260164, 0.3559992, 0.3039555, 0.295264, 
    0.2748332, 0.3241748, 0.4026427, 0.2202291, 0.2316495,
  0.05382342, 0.06927019, 0.09079247, 0.1327851, 0.1217011, 0.144405, 
    0.1310022, 0.05437953, 0.0663799, 0.08877224, 0.1328548, 0.1278255, 
    0.1836577, 0.1825615, 0.1298938, 0.1400961, 0.1387295, 0.1242416, 
    0.08318663, 0.1114477, 0.1200841, 0.06899299, 0.1283495, 0.1277634, 
    0.2831761, 0.3569706, 0.2827878, 0.0783613, 0.04814629,
  0.1453833, 0.2039289, 0.1645622, 0.1853738, 0.2285107, 0.1808328, 
    0.1434556, 0.09157152, 0.1075084, 0.06372109, 0.06379626, 0.066947, 
    0.04387895, 0.03123013, 0.05868764, 0.06344168, 0.06771199, 0.04672335, 
    0.03415096, 0.06373052, 0.05946506, 0.04741064, 0.04150009, 0.1912793, 
    0.06049864, 0.1085084, 0.1101311, 0.1084088, 0.1403536,
  0.04936937, 0.0167241, 0.006376709, 0.009671693, 0.03285327, 0.01904111, 
    0.0249674, 0.02780281, 0.01163715, 0.01022713, 0.007774242, 0.002104445, 
    0.001227614, 0.006326307, 0.2339239, 0.01322555, 0.01906338, 0.02842465, 
    0.02719857, 0.04166181, 0.04549719, 0.01671762, 0.01545131, 0.2512605, 
    0.005031301, 0.02294186, 0.01182073, 0.0128805, 0.07383064,
  0.002630349, 0.001564011, 0.005967437, 0.001071369, 0.0005932553, 
    0.001907903, 0.003622675, 0.002097066, 0.004860678, 0.00190141, 
    -0.0001520632, -3.487572e-06, 0.01294394, 0.0005387686, 0.002626463, 
    0.00666323, 0.003118, 0.006740224, 0.01907268, 0.003690993, 0.001576682, 
    0.001246604, 0.002211293, 0.01610046, 0.03157598, 0.0005178128, 
    0.002710124, 0.0005804445, 0.0009674369,
  0.00828471, 0.002800422, -7.332312e-05, 0.0004800437, -0.0006172937, 
    0.0006889601, 0.0004246017, 0.0002845486, 0.001805817, 0.0001903099, 
    -4.347579e-07, 1.07264e-08, 0.0004230275, 0.001163027, 0.0002083776, 
    0.0003716401, 0.001603618, 0.0004672036, 0.0002405935, 7.437604e-05, 
    3.264442e-05, 0.0003599649, 0.00341484, 0.02051663, 0.02233272, 
    0.04371436, 0.0002473527, 0.0005303818, 0.00285626,
  0.01661268, -1.587421e-05, 0.005086375, 0.03028422, 0.000453934, 
    0.0002732883, 0.0005220705, 3.095882e-05, 0.0002917794, -0.0002704552, 
    0.0009235626, 0.0001281133, 0.01106874, 0.0002153464, 0.0001644321, 
    8.74008e-05, 0.000137934, 0.0007550081, 0.000312974, 5.158679e-05, 
    7.335515e-05, 0.0005532543, 0.01312232, 0.04693352, 0.03189736, 
    0.0005883768, -8.382256e-05, 0.0003561069, 0.00399442,
  0.001356532, 0.04590253, 0.03683059, 0.006052608, 0.0007485761, 
    0.0004241099, 0.000390336, 0.0002757749, 0.02406403, 0.08244108, 
    0.0003051363, 0.001653701, 4.862404e-05, 0.0003759481, 2.755653e-05, 
    9.82444e-05, 0.0003046251, 0.0005779826, 0.0002169916, 0.0002351877, 
    0.0008366598, 0.003490533, 0.03997412, 0.07754975, 0.0577202, 
    0.005127654, 0.002913213, 0.001010702, 0.002174228,
  0.002135935, -3.842429e-05, -1.220768e-05, 0.01020058, 0.0002558878, 
    0.0005105145, -0.002420088, 0.0004793591, -0.0003695176, 0.0009635169, 
    0.0001867721, 0.0007878217, 0.0001874458, 0.0004196891, 0.0002992065, 
    0.0004485226, 0.001000478, 0.001092009, 0.000402091, 0.001059248, 
    0.001972203, 0.0006248767, 0.1183095, 0.04503543, 8.559496e-06, 
    0.000398672, 0.001240008, 0.01551222, 0.02518468,
  2.002633e-07, 7.691814e-07, 3.267408e-07, 0.0007887669, 7.620156e-07, 
    -1.243373e-06, -2.341092e-05, 0.000462298, 0.09300543, 0.005895814, 
    0.001595837, 0.00113877, 0.0001913541, 0.0001802731, 0.0001785426, 
    0.0002159015, 3.714962e-05, 7.38518e-06, 0.003814137, 0.03258916, 
    0.0004706553, 0.01242919, 0.0002232043, -0.001710625, 0.000601188, 
    0.0001202128, 0.0002105745, 0.003006797, 1.417907e-08,
  8.840386e-07, -2.298818e-05, -1.039283e-06, 6.98882e-07, -1.815484e-05, 
    3.746135e-07, -0.0001404182, 0.006092978, 0.2709701, 0.009922839, 
    0.08524878, 0.03944307, 0.043518, 0.02454329, 0.04482286, 0.01497894, 
    0.00988273, 0.002521496, 0.01425872, 0.01611591, -9.344707e-09, 
    0.07195821, 0.03778772, 0.005616492, 0.004336256, 0.003313658, 
    0.006834057, 0.00445551, 0.004680655,
  0.002554906, 0.0001300595, 0.001838306, 0.1056548, 0.0003069248, 
    9.653697e-07, 0.04256311, 0.0006499609, 4.005506e-06, 0.004076219, 
    0.1337805, 0.06094531, 0.1466221, 0.1488101, 0.1019739, 0.09308641, 
    0.08072709, 0.1298402, 0.02807775, 0.0789689, 0.02682514, 0.08618566, 
    0.04873573, 0.07909338, 0.03742735, 0.04615896, 0.02261606, 0.00919482, 
    0.03534452,
  0.04400703, 0.06577811, 0.01826607, 0.009076271, 0.005019068, 0.00889249, 
    0.0156241, 0.05622635, 0.006113926, 0.01519975, 0.1341644, 0.2010705, 
    0.2123491, 0.05890588, 0.03650357, 0.09332231, 0.1189571, 0.1145983, 
    0.06174707, 0.06277268, 0.02490179, 0.0097124, 0.0125646, 0.09217874, 
    0.1159112, 0.2113916, 0.03454702, 0.0554505, 0.1005281,
  0.08408095, 0.09143731, 0.0445746, 0.07645033, 0.04807056, 0.0460154, 
    0.09715645, 0.07744624, 0.09757461, 0.09757305, 0.07722007, 0.08148714, 
    0.1128946, 0.04363911, 0.03085663, 0.2156849, 0.1590872, 0.1892063, 
    0.1327448, 0.07202175, 0.01678251, 0.04305496, 0.1097747, 0.1461951, 
    0.1057143, 0.09190481, 0.1015629, 0.05850084, 0.1161977,
  0.1674874, 0.03465379, 0.1161884, 0.0121142, 0.03492526, 0.0804406, 
    0.1117083, 0.03733999, 0.03346968, 0.09385383, 0.08889219, 0.06124326, 
    0.1960868, 0.1366629, 0.1908994, 0.1900247, 0.3343122, 0.08180868, 
    0.0918924, 0.1302301, 0.1698653, 0.3060817, 0.1574262, 0.2710875, 
    0.1603433, 0.04786262, 0.1769427, 0.0625013, 0.2912948,
  0.1305575, 0.1212392, 0.09577704, 0.1268598, 0.1224154, 0.1186837, 
    0.1577516, 0.1570891, 0.1868457, 0.199757, 0.2183763, 0.2037303, 
    0.2181299, 0.2686846, 0.298996, 0.2569416, 0.2424883, 0.2507157, 
    0.1924961, 0.2395472, 0.2410456, 0.1278573, 0.1172247, 0.08286147, 
    0.05066213, 0.0361388, 0.03805861, 0.1476355, 0.1021395,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -8.812913e-06, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.001126177, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3.072968e-06, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0004607148, 0, 0, 0.0007469145, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -7.097198e-05, 0.001711336, 0, 0, 0, 0, 0, 
    0, 0, -1.039074e-05, -4.399705e-05, 2.66796e-06, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.001485464, 0, 0.0001795419, -5.566732e-06, 
    -1.225321e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, -7.492964e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.455063e-05, -2.068371e-05, 
    5.107669e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001913651, 0, 0, 0.005784527, 5.758918e-06, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  -4.00477e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0002182072, 0.008717751, 
    -6.493764e-06, 0, 0, 0, 0, 0, -1.59005e-05, -5.453753e-05, 0.0001015678, 
    3.59322e-05, 0, 0, -1.406776e-06, 0, 0.0001345728, 0,
  0, 0, 0, 0, 0, 0, -2.648189e-05, 0.003051016, 0, 0.001044546, 0.0006177453, 
    0.0002994577, -0.0001033149, 0, 0, 0, 0, 0, 0, 0, 0, 0.001060594, 0, 0, 
    0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, -4.495779e-05, -2.612166e-05, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, -3.016967e-05, 0, 0, -0.0001113879, -7.745618e-06, 0, 0, 0, 
    -2.791674e-05, 0.001611058, -8.714134e-05, 0.0009348636, 3.131247e-06, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, -1.736889e-05, 0, 0, 2.192422e-06, 0.003969975, 0, 0, 
    0.0105859, -9.345046e-07, 0, 0, 0, -7.065328e-05, 0, 0, 0, 0, 0, 
    2.373664e-05, 0.0006741537, 0, 0, 0, 0,
  -5.103788e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0002704248, 0.02178077, 
    0.00286543, -5.807375e-06, 0.002249037, -2.518434e-05, 0, 0, 
    -8.188379e-05, 0.0001088384, 0.001182713, 0.003019504, 1.833559e-05, 
    0.000853706, -4.497881e-05, 0.0001715081, 0.0006482143, 0,
  0, 0, 0, 0, 0, 0, 0.00187856, 0.007853636, 0, 0.002036522, 0.003361192, 
    0.001213068, -0.0001050592, 0, 0, 0, 0, 0, 0, 0, 0, 0.001348212, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, -0.0001223688, -6.166745e-05, 0.0002568707, 
    -2.306517e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3.135618e-08, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.000440832, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, -7.867676e-05, 0, 0, 0.000500045, -3.872809e-05, 0, 0, 0, 
    -0.0002325778, 0.004737918, -0.0001181356, 0.004881943, 0.0002463477, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -7.554071e-06, 0, 0, 0.000113764, 0, 0, 3.188452e-06, 0.004528897, 0, 
    0.001328706, 0.01929879, 1.450389e-05, 4.462772e-06, 0, 0, -3.418969e-05, 
    0, 0, 0, 0, 0, 0.0004894147, 0.002997298, 0, 0, 0, 0,
  -2.579701e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0005725634, 0.03978977, 
    0.006203149, -7.360354e-05, 0.004251489, -0.0001114491, 0, -1.112699e-05, 
    -0.0001125049, 0.0005197799, 0.002563111, 0.01197691, 7.334235e-05, 
    0.00328777, 0.001909112, 0.0009069921, 0.002165241, 0,
  0, 0, 0, 0, 0, 0, 0.003826058, 0.01555133, 0, 0.004269961, 0.005865844, 
    0.002802784, 0.005049002, 0, 0, 0, 0, 0, 0, 0, 0, 0.002947324, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, -0.000200454, 0.003874191, 0.001932493, 0.0009619064, 
    -3.890341e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -6.204598e-05, -7.061278e-08, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, -3.71543e-05, 0, 0, 2.691951e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -2.65506e-07, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002215964, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, -0.0001292789, 1.81767e-05, -3.688933e-05, 0.001596696, 
    -0.0001124185, 0, 0, -1.943388e-05, 0.0006295716, 0.0091664, 
    0.0001580991, 0.00733267, 0.001915493, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -1.541661e-05, 0, 0, 0.0004439107, 0, 0, 3.049409e-07, 0.00512745, 0, 
    0.002980052, 0.04194767, -6.473747e-05, -9.365085e-06, -2.332121e-06, 0, 
    5.79933e-05, 0, 0, 0, 0, 0, 0.001688375, 0.006597427, 0, 0, 0, 0,
  -3.573859e-05, 0, 0, 0, 0, 0, 0, -5.708266e-06, 2.571615e-06, 0, 0, 
    0.0002791985, 0.06215868, 0.01330028, 0.0004630955, 0.005518581, 
    -0.000303302, -1.072781e-05, 0.0005230149, -0.000176292, 0.008042683, 
    0.01250442, 0.02130225, 0.0002265248, 0.005401774, 0.002368147, 
    0.002434707, 0.009364825, -1.594308e-05,
  0, 0, 0, 0, 0, 0, 0.0047994, 0.02351489, -9.429266e-06, 0.008291571, 
    0.008940105, 0.005420444, 0.01458835, 0, 0, 0, 0, 0, 0, 0, 0, 0.00606632, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, -0.0003087553, 0.01400593, 0.004625904, 0.006323732, 
    -4.762689e-05, -2.917326e-10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -1.37033e-05, 0.001768179, 0.003031929, 
    -4.494741e-05, 8.756015e-06, 7.969885e-05, 0, 0, 0, 0, 0, 0, 
    0.0003742935, 0, 0, 0.00190959, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002679513, 0, 0, 0, 0, 0, 0, 0, 
    -4.016853e-05, 0.001734353, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -4.822121e-07, 
    0.002528579, 0, 0, 0, 0, 0.0008002101, 0, -2.096956e-05, 0.003316031,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.471572e-07, 0.0002375201, 0, 
    -9.563856e-05, -5.686458e-05, 0, 0, 0, 0, 0, 0, -8.902511e-06, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.006025166, 0, 0, 0, 0, 
    -4.126627e-09, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, -0.0001754203, 0.0003856457, -0.0001677053, 0.004332033, 
    -0.0002614227, 0, 0, -0.0002234396, 0.006507819, 0.01941207, 9.72456e-05, 
    0.01749239, 0.005401969, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -5.639642e-05, 0, 0, 0.001913337, 0, 0, 1.019459e-05, 0.005025782, 0, 
    0.006353386, 0.06708563, 0.0001454974, 5.645428e-06, -1.126806e-05, 
    -1.307145e-05, 0.002124347, 0, 0, 0, 0, 0, 0.003550505, 0.01006483, 0, 0, 
    0, 0,
  0.0003114966, 0, 0, 0, 0, -1.999958e-05, 9.179555e-05, 6.898072e-07, 
    0.0003182669, 0.0001254631, 0.0001283146, 0.00840639, 0.08429749, 
    0.02629396, 0.001253625, 0.01068789, 0.0008973192, -8.503233e-05, 
    0.001058523, -4.158341e-05, 0.01400103, 0.02989782, 0.0312487, 
    0.004000712, 0.009300601, 0.003189696, 0.003510545, 0.0198777, 
    -5.492814e-05,
  0, 0, 0, 0, 0, 5.801567e-07, 0.007078798, 0.02952389, 0.001243916, 
    0.02740009, 0.0149193, 0.01214285, 0.03040791, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.01019956, -6.529292e-05, -1.521649e-05, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -3.825652e-05, -0.0002327443, 0.02280442, 0.007728377, 
    0.02111208, -9.737257e-05, 7.603579e-07, 0, -5.373785e-06, 0, 0, 0, 0, 0, 
    0, -3.111571e-05, 6.487492e-07, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0.0005424768, 0.001385731, 0.01068401, 0.01207614, 
    -0.0001761414, 0.004943595, 0.004188805, -3.985412e-05, 0, 0, 0, 0, 0, 
    0.003870136, 0.0005508916, -5.507961e-05, 0.004716563, 0.01387311, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0003852807, -0.0001918041, 0.001407804, 
    0.002505748, 0, -3.634679e-05, -1.924175e-06, 0, 0, 0, 0.0004250486, 
    0.0007515991, 0.004650165, -8.773209e-05, 0.00161688, 0.00227152, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.001607398, 0,
  0, 0, 0, 0, 0.003298384, -6.134189e-06, 0, 0, 0, 0, -3.140813e-05, 0, 0, 0, 
    0, 0.0005190606, 0, 0, -2.526301e-05, -3.17146e-05, 0.01347898, 
    -0.0001051554, 0, 0, 0, 0.00500027, 0.004339239, 0.001797626, 0.005058169,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.149762e-05, -2.053543e-06, 0, 0, 
    0.0001989743, 0.006616048, 0, 0.001273005, 0.0008004965, 0.0003647441, 
    -6.322654e-06, 0, 0, 0, 0, 0.001807916, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01324337, 0.000370434, 
    -1.936161e-05, 0, 0, -1.955618e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, -0.0002287878, 0.009233164, 0.0001619766, 0.009847146, 
    0.001452162, -0.0001949453, -1.418609e-10, -0.0004745057, 0.01918051, 
    0.03593089, 0.0002348461, 0.03283753, 0.01381665, 0.0002832123, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, -1.533119e-05, -0.0001177039, 0, 0, 0.003632499, 3.868117e-06, 
    1.381752e-06, 0.001393284, 0.005012417, 4.994254e-05, 0.01302333, 
    0.1050376, 0.007918759, 0.008530801, -3.222611e-05, -4.388954e-05, 
    0.008138332, 0, 0, 0, 0, 3.133558e-06, 0.008727384, 0.01464276, 
    -3.395895e-05, -3.276829e-05, 0, -5.192304e-05,
  0.004892287, 0.0001428289, 0.0004297913, 0, -2.413709e-06, 0.0006639606, 
    0.003166629, 0.001521295, 0.0005672073, 0.001777423, 0.00252263, 
    0.0259768, 0.1118562, 0.05002065, 0.006699939, 0.01609475, 0.01194593, 
    0.0005500433, 0.001591829, 0.001544865, 0.02268576, 0.05809182, 
    0.0421467, 0.01459562, 0.01452575, 0.006942828, 0.005418816, 0.05928662, 
    -0.0001649661,
  0, 0, 0, 1.449786e-05, -6.456632e-09, 7.261078e-05, 0.01174909, 0.04835826, 
    0.004016621, 0.05210299, 0.04031753, 0.01700041, 0.06832215, 
    3.970212e-07, 0.0004390777, -3.206565e-05, 0, 2.999835e-05, 0, 
    -8.03875e-09, -5.98128e-07, 0.01698637, 1.22349e-05, 0.00227408, 0, 0, 0, 
    0, 0,
  0, -2.374385e-05, 0, 0, 0, 0, 0.001001362, 0.0001324303, 0.03795752, 
    0.01539922, 0.04455755, 0.008184058, 0.0008777739, 0, -1.230738e-05, 
    -3.066928e-06, 0, 0, 0, 0, 0, 0.0008238099, 0.0005072411, 0, 
    -7.427429e-06, 0, 0, 0, 0,
  -2.255601e-06, -7.838865e-05, 0, 0, 0, 0, -3.517768e-06, -3.640487e-09, 
    0.003616599, 0.009160783, 0.02201179, 0.02460274, 0.01139226, 
    0.009027487, 0.007341367, -6.74392e-05, 0, 0, 0, 0, 0, 0.006913357, 
    0.002212253, 0.0006566066, 0.009237014, 0.01846541, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0.004270971, 0.004882706, 0.008494841, 
    0.008444238, 0.005845699, 0.0002018274, 0.004001668, -6.151557e-06, 0, 0, 
    0, 0.006793748, 0.005579601, 0.01440861, -0.0001526478, 0.003347034, 
    0.004668495, 0, -3.596171e-05, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -7.661251e-06, 0, -1.148957e-06, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  -1.261634e-05, 0, 0, 0.0009884898, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0007464708, 0, 0, 0, 0, 0, 0, 0, 6.173459e-05, 0, 0, 0, -5.020009e-06, 
    0.00362167, -8.6217e-06,
  0, 0, -2.334288e-06, -1.848392e-05, 0.005304106, 0.0001013384, 0, 
    -4.228759e-06, 0, 0, 0.00252223, 0, -2.946447e-06, -2.149371e-08, 0, 
    0.005517758, 0.001283064, 0.0004798514, 0.0002198353, 1.25872e-05, 
    0.0292991, 0.00824781, -1.755197e-05, 0.0009727097, -2.845441e-05, 
    0.01058677, 0.0121091, 0.006582431, 0.007337105,
  0, 0, 0, 0, -1.794271e-06, -3.109493e-05, 0, 0, 0, 0.0002599108, 
    0.001055656, 0.0006289412, 0, -5.822773e-08, 0.005067479, 0.0238074, 
    0.001106947, 0.0141112, 0.005261109, 0.004652286, 0.0008500753, 0, 0, 0, 
    0, 0.005509277, -4.082713e-05, 0, 0,
  0, 0, 0, 0, 1.376321e-08, 0, 0, 0, -9.867575e-06, -2.511498e-05, 0, 0, 0, 
    -3.107593e-09, 0.01961061, 0.008015948, 0.007694762, 0.0001588573, 
    0.0001234453, 0.002366066, 0, 0, 0, -1.712747e-06, 0, 0, 0, 0, 0,
  0, 0, 0, 0, -0.0001937068, 0.02369696, 0.004703358, 0.02136326, 
    0.002794651, 0.0001324746, 4.739884e-06, 0.002778428, 0.03789591, 
    0.05812293, 0.01118132, 0.06770382, 0.03857833, 0.000740663, 0, 
    -5.796879e-08, 1.251279e-09, 0, -1.565992e-06, 5.164917e-08, 0, 
    -5.335785e-05, 0, 0, 2.834061e-06,
  1.691072e-06, 2.953944e-05, -0.0001821945, 0, 0, 0.01290924, 0.001012413, 
    9.551435e-05, 0.007518171, 0.005230449, 0.004893206, 0.03131245, 
    0.1356885, 0.03139951, 0.02316392, 0.0001937456, -0.0001576528, 
    0.01227307, 0, -3.978839e-06, -2.684295e-06, 3.777059e-05, 0.0002233733, 
    0.04687778, 0.02613538, -8.623623e-05, 2.335495e-06, -4.035147e-05, 
    -0.000165381,
  0.0141648, 0.0003530949, 0.0005331247, -3.008266e-08, -3.862392e-05, 
    0.004261693, 0.01956249, 0.03278329, 0.02270257, 0.00507956, 0.004360642, 
    0.04128829, 0.1547857, 0.07567371, 0.02073114, 0.02311915, 0.05084749, 
    0.006302748, 0.004608923, 0.0109649, 0.04280092, 0.1094543, 0.09285641, 
    0.03074518, 0.02103555, 0.01575487, 0.01040097, 0.08287054, 0.003678333,
  -1.073193e-07, 0, 0, 0.0001157219, 3.177475e-06, 0.01395778, 0.03124498, 
    0.1723916, 0.02826252, 0.1003945, 0.07950205, 0.03376449, 0.08878803, 
    5.52268e-05, 0.0002037256, 0.003226799, -4.078108e-05, 0.001512526, 
    0.001718316, 8.965466e-05, 0.00126421, 0.02559478, 0.002420522, 
    0.01255902, 0, 8.637326e-08, 0, 0, 0.001328761,
  0, -0.0001283355, 0, 0, -2.399602e-08, 0, 0.00988489, 0.002917299, 
    0.09199912, 0.04712857, 0.07316633, 0.02425399, 0.003725512, 
    0.0004316658, 0.000332923, 0.001400443, 0, 0, 0, 0, 0, 0.008729665, 
    0.001637855, 0, -5.797084e-05, 0, 0, 0, -1.51632e-11,
  2.268714e-05, 0.00137664, -1.041077e-09, -5.181694e-13, -8.192053e-06, 
    -9.715495e-05, 7.770761e-05, 0.0001035591, 0.006591741, 0.01383535, 
    0.02974583, 0.04442681, 0.03329359, 0.01652637, 0.01207813, 2.081548e-05, 
    0, 0, 0, 0, 0, 0.01496595, 0.007818178, 0.001715718, 0.01327575, 
    0.02389848, -2.8922e-06, -4.509328e-06, 0,
  0, -7.911193e-06, 0.001315095, -6.589963e-05, 4.213269e-06, 3.077276e-05, 
    0, 0, 0.001012472, 0.007137371, 0.008456485, 0.01620307, 0.02711721, 
    0.01067294, 0.002806312, 0.006830609, -3.954246e-06, 0, 0, -1.214408e-05, 
    0.01584968, 0.01137159, 0.02291385, 0.004644112, 0.003958816, 
    0.009040401, 0, 0.0005332427, 0,
  0, 0, 0, -5.629237e-05, 0, -3.689745e-06, 0, 0, 0, 0, 0, -3.587229e-06, 
    -0.0001271111, -3.4094e-06, -3.512397e-05, 0, -5.327747e-05, 0, 0, 0, 0, 
    -6.480088e-05, -0.0002664192, 4.366143e-06, -2.553339e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0, -8.921007e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, -1.708612e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  -5.984889e-05, 0.00492191, -6.684439e-06, 0.003125063, -6.691748e-07, 
    0.0008054859, 0, 0, 0, 0, 0, 0, 0.0002098217, -1.624527e-05, 0.002728772, 
    -2.071431e-06, 0, -1.308881e-05, 0, 0, -0.0001756035, 0.0001254289, 
    0.00095325, 0, 0, 0, 0.003211121, 0.004875921, 0.000581735,
  0, 0, 0.0008551262, -0.0001775621, 0.01127262, 0.005117955, 0, 
    -0.000102761, 0.0004426063, 0, 0.004101741, -9.51966e-05, 0.002232417, 
    0.001826176, -7.868379e-05, 0.01710192, 0.008475858, 0.002721714, 
    0.004757122, 0.006640315, 0.04670865, 0.02966272, 0.006008795, 
    0.009452572, -0.0001070895, 0.0194969, 0.02507688, 0.01090559, 0.01118726,
  0, 0, 0, -5.945453e-06, -7.372398e-05, 0.0001121784, 0, 0, -6.886314e-09, 
    0.003816688, 0.005304267, 0.007865439, 7.406891e-05, -3.443039e-05, 
    0.01241004, 0.04067958, 0.005018565, 0.03704, 0.02658196, 0.02547602, 
    0.003998454, 8.738801e-05, -1.821203e-10, 0.0008060293, 0.000112433, 
    0.01059903, 0.001770083, 0, -1.144106e-06,
  0, 0, 0, 0, 1.952278e-05, 1.026753e-05, -1.831262e-08, 2.045902e-07, 
    0.0003606927, -9.009355e-05, -2.876059e-07, 2.369934e-08, -7.351193e-06, 
    1.324069e-05, 0.03448463, 0.02819225, 0.0302358, 0.007782684, 
    0.003318889, 0.01338746, -5.552068e-06, 3.139207e-07, -2.450789e-07, 
    0.0001566542, 2.272098e-05, -2.416512e-11, 0, -1.230101e-10, -3.276734e-09,
  0, 0, 0, -1.824492e-07, 0.001153735, 0.03396646, 0.0301094, 0.04902705, 
    0.03921635, 0.02340924, 0.0002474889, 0.0136312, 0.1009829, 0.1754346, 
    0.1348992, 0.2316451, 0.1458172, 0.00701337, 7.495617e-07, -5.492733e-05, 
    6.372602e-05, -2.521627e-05, -4.041404e-06, 1.430968e-05, 0.000239259, 
    -6.675543e-05, -8.374704e-09, 2.470479e-08, 0.002266952,
  0.003034451, 0.001496152, 0.0008219455, 0, -5.455722e-06, 0.02268426, 
    0.06111486, 0.05461352, 0.04722575, 0.02751637, 0.06657978, 0.1604927, 
    0.258325, 0.1436739, 0.1737248, 0.02580569, 0.00297426, 0.01765919, 
    0.00073026, 2.612116e-05, 0.0008107654, 0.03629674, 0.04115784, 
    0.1484981, 0.07777499, 0.0006405634, -4.111659e-06, 0.003220622, 0.0150828,
  0.04849494, 0.004570278, 0.0008615789, -1.470901e-05, 0.008793069, 
    0.1867911, 0.3212869, 0.5896968, 0.340271, 0.168748, 0.06220886, 
    0.1355967, 0.3511024, 0.213357, 0.1686587, 0.131778, 0.1397528, 
    0.03339285, 0.02964659, 0.0402282, 0.1344673, 0.2709567, 0.2562635, 
    0.1683589, 0.07487309, 0.02657318, 0.03804309, 0.1586768, 0.03021288,
  1.138825e-05, 0, 1.770546e-05, 0.006966916, 0.01460731, 0.0914845, 
    0.133607, 0.2838689, 0.2351412, 0.3235635, 0.2091955, 0.1576107, 
    0.1670292, 0.02627652, 0.001274416, 0.01250816, 0.00621809, 0.0110518, 
    0.02107185, 0.002267663, 0.03501677, 0.1385363, 0.03288572, 0.0407274, 
    -4.053296e-07, 0.0003876336, 5.53063e-05, 2.489281e-06, 0.004514771,
  0.001083069, 0.001189029, -1.515804e-05, 0, 0.000337186, 2.291022e-06, 
    0.07673273, 0.005086407, 0.1519197, 0.168178, 0.2212566, 0.125053, 
    0.07993901, 0.03654163, 0.001685759, 0.004165648, 0, 1.064234e-08, 0, 
    6.121448e-07, 0, 0.0791624, 0.01606917, -6.644871e-05, 0.001122382, 
    1.720013e-05, 0.001084313, 4.88325e-06, -2.400229e-08,
  0.00595735, 0.01326932, 0.0006928318, 6.23089e-05, -0.0001388057, 
    0.0003152539, 0.003508471, 0.0220679, 0.02693437, 0.02392924, 0.06936861, 
    0.1328408, 0.140054, 0.0762701, 0.0240712, 0.003621516, 0.001484575, 
    -1.373882e-06, 0, -1.317379e-06, -3.831262e-05, 0.02926378, 0.01806265, 
    0.01357592, 0.01795509, 0.0331032, -6.001073e-05, 8.573711e-05, 
    -1.195997e-11,
  -3.198161e-06, 7.748725e-05, 0.02088491, 0.004668912, 0.0007508239, 
    0.0001871577, -9.085136e-06, 1.038351e-06, 0.003275403, 0.01472209, 
    0.02055063, 0.01983938, 0.04226175, 0.02113278, 0.005472669, 0.01477081, 
    0.001876662, 0.002803699, 0, -0.000136934, 0.02552397, 0.01713132, 
    0.03284063, 0.0112078, 0.01633545, 0.02086632, 0.001674436, 0.002778919, 0,
  -1.715997e-05, 0, 0, 0.00215458, 5.90736e-05, 0.001561248, -8.852604e-05, 
    -1.988503e-08, 0, 0, 0.001790204, 0.0005934249, 0.001812615, 
    -6.371216e-05, -0.0001484966, 0, 7.084046e-05, 0.001310251, 0, 0, 
    -9.178986e-05, -0.0002793123, 0.0006825785, 9.443701e-05, -0.0002775019, 
    -0.0001808798, 0.0004241889, 1.147386e-05, 0,
  0, 0, 0, 0, 0, 0.002718655, 0, 0, 0.0009884181, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -9.278428e-06, 0, -0.0001424602, 0.0001581491, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, -5.31191e-06, 0, -1.286617e-06, 0, 0, 6.545571e-05, 0, 0, 0, 
    0.0001011646, -3.76014e-05, -0.0002217324, -1.45349e-05, 0, 0, 0, 0, 0, 
    0, -6.968215e-06, -1.892013e-05, 0, 0, 0, 0, 0, 0,
  -0.0002309828, 0.01047713, 0.0007985387, 0.00373547, 0.0009395826, 
    0.002704088, -6.739482e-05, 0, 0, -7.929578e-06, 0.001143416, 
    0.003485727, 0.003364403, 0.003961558, 0.004088917, 1.060884e-05, 
    -5.02141e-05, 0.003685946, 0.0006299881, 0, 0.003845942, 0.001289943, 
    0.001713086, 3.115897e-05, -8.165151e-06, -2.201438e-05, 0.006790781, 
    0.01568527, 0.001854493,
  0.0007801171, -7.85618e-05, 0.01164724, 0.001731992, 0.01716755, 
    0.02159392, -3.676199e-05, 0.001417759, 0.003154553, -5.06301e-07, 
    0.01322469, 0.003650087, 0.004412979, 0.00767608, 0.003820947, 
    0.03218969, 0.02219266, 0.008955666, 0.01994432, 0.01642084, 0.07465538, 
    0.06703318, 0.02138136, 0.01641341, 0.001235367, 0.03004201, 0.03790345, 
    0.02509853, 0.01444101,
  0.00575536, 0.0003111249, -3.411778e-06, 0.0001005502, 5.354249e-05, 
    0.001760424, -7.915307e-08, -2.906361e-07, -1.307774e-05, 0.002667659, 
    0.02683259, 0.04468166, 0.002350557, 0.001109689, 0.02438779, 0.08393724, 
    0.02816085, 0.07155031, 0.06144312, 0.05959162, 0.009929548, 0.008741512, 
    0.0003110023, 0.006974231, 0.01212102, 0.02603843, 0.01290608, 
    0.0008335199, -5.560875e-05,
  0.0006086521, 8.050304e-05, 7.072007e-07, 1.004041e-08, 0.0001202831, 
    1.255866e-05, 5.491341e-07, -1.25298e-05, -0.0001434534, -0.0001084997, 
    1.823088e-05, -5.23672e-07, 0.0001247427, 0.000105933, 0.08197169, 
    0.1061492, 0.07447921, 0.04762837, 0.01842281, 0.02795231, 2.534889e-05, 
    2.161456e-05, 1.407269e-05, 0.05612361, 0.0005794443, 0.0001829571, 
    3.855406e-05, 6.712153e-06, 4.510402e-06,
  5.408313e-05, 2.662425e-05, 1.534129e-05, 1.031491e-05, 0.004960345, 
    0.08453275, 0.04657682, 0.06421486, 0.06738397, 0.02265089, 0.005762917, 
    0.0192535, 0.0989423, 0.1697066, 0.1252815, 0.2154309, 0.1175573, 
    0.009018534, 1.148528e-05, 0.0006098357, 0.0002300357, 7.707166e-05, 
    0.008884318, 0.0175743, 0.0004943325, 0.004258878, 1.112216e-05, 
    0.0001154482, 0.001754526,
  0.06009059, 0.08358273, 0.20452, 1.384497e-05, 0.0007090911, 0.09711906, 
    0.2279867, 0.08375254, 0.208827, 0.1322393, 0.05696746, 0.1360606, 
    0.2399303, 0.1214236, 0.1432466, 0.01308036, 0.0004539388, 0.01755612, 
    3.712026e-05, 0.002456186, 0.017354, 0.07193669, 0.09932242, 0.3016155, 
    0.1360632, 0.008745321, 0.005655758, 0.04310809, 0.028929,
  0.1962668, 0.06002298, 0.06576005, -1.851503e-05, 0.03998651, 0.1687409, 
    0.341281, 0.5187908, 0.3043158, 0.1455642, 0.0406668, 0.1076132, 
    0.2893751, 0.2031994, 0.1510366, 0.1875596, 0.1230712, 0.02929563, 
    0.03464049, 0.04875088, 0.1220816, 0.2595649, 0.3844069, 0.261323, 
    0.1393203, 0.1200911, 0.06496394, 0.2485097, 0.2117393,
  0.02050458, 1.033027e-05, 0.001345123, 0.003663829, 0.01032488, 0.09276656, 
    0.1258642, 0.247088, 0.1991443, 0.2592397, 0.1898204, 0.1279793, 
    0.1563373, 0.09247985, 0.06746648, 0.0668966, 0.09307504, 0.05425475, 
    0.06429481, 0.02817475, 0.02560037, 0.1846546, 0.1653963, 0.2107585, 
    0.06754348, 0.001807127, 0.0002703803, 0.003840378, 0.03476932,
  0.03184865, 0.03121702, 0.01152851, -1.181951e-08, 0.000261506, 
    2.556267e-06, 0.07203785, 0.01357149, 0.2309601, 0.1789554, 0.2588798, 
    0.1647609, 0.1492643, 0.1454344, 0.181993, 0.07920974, 0.001991325, 
    -5.587866e-07, -1.51992e-05, 0.01065346, -7.035098e-05, 0.1493308, 
    0.1173671, 0.1853245, 0.07896356, 0.02895229, 0.008297461, 0.007039487, 
    7.887976e-05,
  0.01405795, 0.03072166, 0.009164052, 0.001670725, 0.007569872, 0.00589292, 
    0.01443096, 0.04633458, 0.08450768, 0.05803632, 0.1145751, 0.1755546, 
    0.2411429, 0.1692566, 0.09773958, 0.1254255, 0.03046888, 0.003948798, 
    -7.735392e-05, 1.587164e-06, -4.283002e-05, 0.07398898, 0.1020132, 
    0.05748148, 0.05908858, 0.07314818, 0.02506145, 0.02517411, 0.002407075,
  0.01028184, 0.0004204052, 0.03851798, 0.01000891, 0.001739447, 0.002959346, 
    -0.0003801181, 0.0002168661, 0.005626006, 0.02748531, 0.04089435, 
    0.03754204, 0.07261562, 0.09967751, 0.05599416, 0.04267672, 0.0156185, 
    0.01039201, -2.998178e-05, -0.0002777852, 0.03830039, 0.0299807, 
    0.06153512, 0.01923343, 0.04279997, 0.04534591, 0.006321877, 0.01710948, 
    0.01207787,
  -0.000113663, 0.0003996515, -0.0001319006, 0.006669399, 0.0007136085, 
    0.00149775, 0.002181494, 0.000112998, -1.049219e-05, 0, 0.004355544, 
    0.005152368, 0.006651627, 0.002181015, 0.007736786, 3.96338e-06, 
    -7.467181e-05, 0.002626992, -0.0001107671, 0.002676073, 0.008397905, 
    0.002972466, 0.008704387, 0.00528665, 0.0003144038, 0.00460169, 
    0.004355468, 0.001488272, 0.0005358364,
  -3.979324e-05, 0, 0, 0, 0, 0.003691362, 0, 0, 0.002305303, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, -1.469261e-05, -0.0002933273, 0.007787027, 0.0009164382, 0, 
    0, 0.002619352, 0, 0, -0.0001799887, -0.0003109229,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3.579901e-05, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -3.653127e-06, -2.60273e-05, 0.0002017927, 0, 0, 0.0007855099, 0, 0, 
    0, 0.002688669, 0.001003807, -0.00031489, -3.209318e-05, 3.692119e-05, 
    -4.104072e-05, 0, 0, 0, 8.669705e-06, 0.002591235, -0.0002004347, 
    -2.412003e-06, 0, 0, -1.331579e-05, 0, 0,
  0.006621792, 0.01498384, 0.007578727, 0.005127855, 0.001289616, 
    0.008395996, 0.001595647, 0.002307606, 0.002068674, 0.00257014, 
    0.006018571, 0.01175995, 0.01135339, 0.006192538, 0.01220664, 0.00193445, 
    0.006426258, 0.01168008, 0.002277786, -0.0001684796, 0.01036981, 
    0.01740738, 0.01039253, 0.005570021, 0.001569424, 0.001657646, 
    0.01745189, 0.03294523, 0.007125191,
  0.005647736, 5.174306e-07, 0.01825849, 0.01953539, 0.02394824, 0.03067809, 
    0.01026956, 0.01008553, 0.009659258, 0.000594861, 0.01854972, 0.01321097, 
    0.008590183, 0.01640237, 0.0112175, 0.05899841, 0.04887745, 0.03194027, 
    0.03870494, 0.032035, 0.116361, 0.1248039, 0.04856469, 0.03986083, 
    0.008480689, 0.04721514, 0.06813004, 0.05724438, 0.02740161,
  0.008472499, 0.001030651, -7.456896e-05, 0.0003375406, 0.002074927, 
    0.03340058, -0.0001232559, -0.0001084136, 0.000705881, 0.003039793, 
    0.06580044, 0.1050894, 0.02862001, 0.02602778, 0.07010309, 0.1119888, 
    0.07908484, 0.1037558, 0.1321273, 0.1570603, 0.1334512, 0.02015854, 
    0.004736838, 0.01612367, 0.04801403, 0.03856566, 0.08057989, 0.02703418, 
    0.000503285,
  7.066881e-05, 6.351928e-06, 4.585961e-06, -1.521344e-09, 0.0003415809, 
    -3.596703e-06, 1.184256e-05, -1.248942e-06, -0.0001226238, 0.000198641, 
    -1.755489e-05, -1.356565e-07, 2.892475e-05, 4.040665e-05, 0.0752655, 
    0.09501492, 0.1188146, 0.06503114, 0.04143445, 0.04945535, 4.052229e-05, 
    1.513934e-06, 4.520688e-06, 0.008097793, 0.000227642, 0.009421325, 
    3.408146e-06, 2.046852e-07, 8.292051e-07,
  3.251112e-05, 6.330572e-06, 8.523669e-06, -5.203562e-06, 0.002758383, 
    0.05804368, 0.03416622, 0.05823298, 0.05244645, 0.02114866, 0.0005865983, 
    0.00387898, 0.09006728, 0.1457047, 0.0925427, 0.1760644, 0.08504695, 
    0.001178196, 2.829102e-05, 0.0001280462, 2.517277e-06, 1.242418e-05, 
    0.01898179, 0.01227281, -0.0001847457, 0.0004497918, 1.698786e-05, 
    1.329614e-05, 4.574846e-05,
  0.02803143, 0.05033847, 0.1191376, 3.335607e-06, 0.0001261242, 0.05633358, 
    0.1397658, 0.0453006, 0.1846061, 0.1011421, 0.03880498, 0.08537224, 
    0.2239295, 0.09896006, 0.1165853, 0.007397728, 0.0002708854, 0.01695905, 
    3.398737e-06, 0.0002426363, 0.001175728, 0.04210591, 0.09609008, 
    0.267706, 0.08502066, 0.003053315, 0.004388448, 0.01606245, 0.007002498,
  0.1289218, 0.03773333, 0.06454813, 0.01438625, 0.02915362, 0.13959, 
    0.2312857, 0.405002, 0.2574572, 0.1022287, 0.03428116, 0.07975858, 
    0.2563344, 0.1729339, 0.1263626, 0.1532044, 0.1061323, 0.02130857, 
    0.02131233, 0.02033482, 0.09532464, 0.2401934, 0.3342724, 0.1843592, 
    0.09550615, 0.06930032, 0.0365328, 0.2210034, 0.1577918,
  0.01674936, 2.795092e-05, 0.0008973958, 0.002892198, 0.002745218, 
    0.09847222, 0.1368509, 0.2218024, 0.1632432, 0.2195534, 0.1703172, 
    0.08947621, 0.1391288, 0.04725925, 0.04478676, 0.05925564, 0.05732577, 
    0.07403556, 0.06517386, 0.01301479, 0.01542377, 0.150894, 0.1253971, 
    0.1655778, 0.04179882, 0.01103166, -8.249657e-07, 0.006470972, 0.04262674,
  0.067143, 0.0778323, 0.01954624, 0.007670166, 4.006454e-05, -1.143866e-05, 
    0.07086138, 0.08040281, 0.3356051, 0.1607254, 0.2387441, 0.1323865, 
    0.1191117, 0.1172952, 0.1665544, 0.08600742, 0.06345641, 0.01141089, 
    0.01692353, 0.01663018, 0.01328588, 0.1520843, 0.07878168, 0.1520733, 
    0.1274609, 0.1130404, 0.0354858, 0.003543293, 0.0003581113,
  0.03788696, 0.07259389, 0.01540419, 0.012689, 0.04215786, 0.02976893, 
    0.02953739, 0.09117993, 0.173414, 0.1099164, 0.1267927, 0.1892848, 
    0.2426665, 0.1906058, 0.1402172, 0.2497481, 0.197713, 0.1007609, 
    0.03450604, 0.0001832699, -6.726874e-05, 0.1443721, 0.1144944, 
    0.08695222, 0.1223436, 0.1403595, 0.07459314, 0.121471, 0.05219509,
  0.04798694, 0.003127084, 0.062663, 0.02748294, 0.03375799, 0.01935871, 
    0.007379147, 0.00984699, 0.01192416, 0.05190995, 0.1139941, 0.1418275, 
    0.1012606, 0.09629863, 0.1239369, 0.1323308, 0.1339272, 0.1574555, 
    0.09426413, 0.0001997536, 0.05785254, 0.1035585, 0.1313305, 0.06980217, 
    0.1137549, 0.1281374, 0.1332099, 0.09927123, 0.05133209,
  0.02766329, 0.0001248779, 0.000694361, 0.01170101, 0.00615981, 0.0036971, 
    0.0159174, 0.0002744838, -5.943647e-05, 0.001834111, 0.0104091, 
    0.02747546, 0.0139473, 0.01503922, 0.0297227, 0.01569547, 0.01960193, 
    0.02246442, 0.001603302, 0.005396947, 0.02059382, 0.0244069, 0.01130025, 
    0.009853327, 0.04090406, 0.007851991, 0.02413233, 0.03280475, 0.01977967,
  0.0002553773, 1.140556e-05, 0, 0, -1.745823e-05, 0.004461703, 
    -0.0001491081, 0, 0.006159193, 0, 0, 0, -2.053884e-05, 0, 0, 0, 0, 
    -6.041254e-10, -0.0001214606, 0.002091483, 0.03389074, 0.002381786, 0, 0, 
    0.004739853, -1.414575e-06, 0, -0.0003060217, 0.005275434,
  -7.753579e-07, 0, 0, 0, 0, 0, 0, -2.22286e-05, 6.055918e-08, -1.763122e-09, 
    2.065824e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.464139e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, -8.511148e-05, 0, 0, 0, 0, 0, 0, -3.74662e-05, 9.514393e-06, 
    0.001293506, 0, 0, 0, -4.338825e-06, -5.135115e-05, 0, 0, 0, 0, 
    0.0001863649, 0, 0, 0, 0,
  0.001694779, 0.006354516, 0.002392261, 0.004271106, 0.001004133, 
    0.0001719804, 0.0005814545, 0.006912757, -7.939793e-05, -5.571983e-07, 
    -3.875052e-05, 0.01197098, 0.006046934, 0.0004936875, 0.001532887, 
    0.003072828, 0.003330682, 0.0002384521, 0.001303632, -0.0002317675, 
    0.001342022, 0.007448762, 0.01403942, 0.00188765, -8.548377e-05, 
    0.0009183256, 0.002283482, 0.0004488373, 0,
  0.03585406, 0.02816343, 0.01817877, 0.006103572, 0.01109639, 0.01249773, 
    0.003859489, 0.008023949, 0.004991851, 0.005445892, 0.01208876, 
    0.02036224, 0.01883178, 0.01288784, 0.02206188, 0.008877418, 0.04571456, 
    0.02981236, 0.01612253, 0.01962139, 0.03183348, 0.05834231, 0.05651941, 
    0.01774503, 0.01958328, 0.008233109, 0.04235994, 0.08126419, 0.04096382,
  0.1031464, 0.03910688, 0.04615645, 0.03990512, 0.03132395, 0.04488402, 
    0.0331498, 0.03201456, 0.01547398, 0.001873101, 0.03844014, 0.03737335, 
    0.02052747, 0.02680959, 0.02475532, 0.1143751, 0.1492932, 0.08526747, 
    0.0972981, 0.05952676, 0.1652819, 0.2051209, 0.1098518, 0.08422464, 
    0.04823471, 0.127816, 0.1684223, 0.1615446, 0.1387483,
  0.02213277, 0.01114125, -6.643539e-05, 0.002357581, 0.01400616, 0.04249289, 
    0.001169762, -7.410387e-05, 0.01044133, 0.02071139, 0.0792148, 
    0.09999238, 0.04455899, 0.04322498, 0.08358521, 0.117058, 0.07484513, 
    0.1051275, 0.1853379, 0.1878877, 0.0856876, 0.02604905, 0.01443415, 
    0.007757858, 0.05647679, 0.05930311, 0.1154506, 0.08269857, 0.01787033,
  8.009332e-06, 8.639546e-07, 1.350001e-06, 1.382301e-08, 0.0003025186, 
    -0.0001993779, -5.063934e-05, 1.429801e-06, 0.0003811324, -2.408894e-05, 
    0.001112563, -2.065036e-07, -5.395024e-05, 0.001035154, 0.06958757, 
    0.07692499, 0.1023552, 0.04972898, 0.02883369, 0.03569467, 6.240092e-06, 
    1.506534e-07, 5.783137e-07, 0.0002652071, 8.551014e-05, 0.01383959, 
    5.675549e-06, -1.167817e-06, 1.00746e-07,
  6.50325e-06, 9.225371e-07, 3.679342e-06, -2.747726e-06, 0.003389988, 
    0.04021754, 0.02004735, 0.05300532, 0.04548389, 0.02962749, 0.0001011698, 
    0.0001695495, 0.08038194, 0.12361, 0.07628266, 0.1570406, 0.07664014, 
    0.0005542688, 0.0001470858, 6.612718e-05, 2.577861e-07, 3.433334e-06, 
    0.009777733, 0.00553272, -7.759389e-05, -8.910828e-05, -1.898171e-07, 
    5.080828e-06, 7.852592e-06,
  0.0208649, 0.03988057, 0.06383794, 5.513876e-06, 0.0006021436, 0.05205107, 
    0.1017593, 0.03446909, 0.1638884, 0.09313195, 0.03238139, 0.06239303, 
    0.2111396, 0.08261951, 0.09322909, 0.00902076, 0.001553648, 0.01762251, 
    6.775503e-06, 0.002321529, 0.00249264, 0.02674687, 0.1088787, 0.2389272, 
    0.06914351, 0.003153142, 0.004573421, 0.000257282, 0.003236692,
  0.1189014, 0.04987295, 0.06125795, 0.001720706, 0.03450854, 0.09025095, 
    0.1694425, 0.2309113, 0.2363095, 0.08414754, 0.03030421, 0.07144726, 
    0.2422968, 0.1574161, 0.1132583, 0.1268782, 0.09938595, 0.01822998, 
    0.01627273, 0.01725978, 0.0923265, 0.2416812, 0.2988535, 0.1581729, 
    0.0836554, 0.04531259, 0.0234727, 0.1867659, 0.1395183,
  0.0140658, -3.005905e-05, -2.479716e-05, 0.002484657, 0.00900449, 
    0.09561074, 0.1347462, 0.2063214, 0.1496195, 0.1776706, 0.1317053, 
    0.0782106, 0.125173, 0.04106287, 0.03897807, 0.03517354, 0.03663334, 
    0.04654825, 0.04796204, 0.003819985, 0.01661303, 0.1184811, 0.1267785, 
    0.1570993, 0.03817994, 0.01197582, 9.533454e-06, 0.00832592, 0.04277227,
  0.05709082, 0.06550375, 0.01001704, 0.003682119, -9.901884e-07, 
    -2.110875e-05, 0.05435975, 0.08981103, 0.3466141, 0.1427711, 0.2310623, 
    0.1242696, 0.108199, 0.1058133, 0.1442203, 0.0791278, 0.07319439, 
    0.03662084, 0.02774451, 0.01169893, 0.03509789, 0.1168909, 0.0557398, 
    0.135643, 0.1192501, 0.08483408, 0.01427337, 0.0007305689, 0.008223883,
  0.08883219, 0.111747, 0.06244, 0.06083605, 0.05074231, 0.05528293, 
    0.04356778, 0.1882424, 0.2122506, 0.1427489, 0.1353329, 0.1866513, 
    0.2390946, 0.1970918, 0.1328334, 0.2131465, 0.2212433, 0.1597832, 
    0.04866315, 0.006883563, 0.007569137, 0.1334396, 0.07552405, 0.08517853, 
    0.1021005, 0.116512, 0.06804332, 0.118395, 0.06819608,
  0.1052721, 0.03080566, 0.09027086, 0.1209184, 0.1104131, 0.07377887, 
    0.06042077, 0.02337465, 0.04463383, 0.1322731, 0.2033057, 0.2508583, 
    0.130033, 0.1133241, 0.1678011, 0.20659, 0.2133784, 0.2600958, 0.1795958, 
    0.02977492, 0.1270489, 0.1131343, 0.1313556, 0.1055773, 0.138063, 
    0.1865572, 0.2189023, 0.1458233, 0.186596,
  0.1525928, 0.01980259, 0.02339035, 0.0630601, 0.07425123, 0.08693282, 
    0.09802177, 0.0289325, 0.005952849, 0.01463972, 0.07340755, 0.09731482, 
    0.07844044, 0.1193948, 0.1027786, 0.04108592, 0.03108756, 0.04136868, 
    0.05218707, 0.0696753, 0.06193073, 0.08561048, 0.08802579, 0.07299184, 
    0.09997306, 0.04212286, 0.0502551, 0.149299, 0.1328984,
  0.03627687, 0.04352205, 0.01122228, 0.01256802, 0.0113771, 0.03056626, 
    0.02610497, 0.01252818, 0.01992284, -0.0003995643, 0.04403416, 
    0.06197111, 0.01200873, 0.02637793, 0.0001346067, -0.0002182673, 
    0.0005475788, -0.0002413607, 0.01701226, 0.05207748, 0.08803864, 
    0.01199102, 0.0001099697, 0.0003010555, 0.007410829, -1.787525e-05, 
    -3.482686e-06, 0.000932203, 0.03738983,
  0.005101427, 0.006170345, 0.002873736, -0.0003095476, -1.452392e-08, 
    -7.321695e-06, -0.0009794408, 0.003966039, 0.001346419, -0.0002330681, 
    0.0006880323, -1.81311e-05, -9.362279e-05, 0.001365749, -1.836201e-07, 0, 
    0, 0, 0, 0, -0.0002445847, 0.002235288, -5.149301e-06, -4.697303e-05, 
    -6.127326e-06, 0, 0, -2.686357e-05, -0.0006897886,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, -0.000207011, 0.0002847069, 0, 0, -1.952933e-05, 
    -1.065325e-06, 0, -7.49324e-05, 5.526057e-06, 0.009606269, 0.001132104, 
    -1.734719e-05, 0, -0.0001810837, 0.002453235, 0.0007527581, 4.192508e-05, 
    -5.694092e-05, 0.001192906, 0.0004618434, 0, -1.690839e-05, 0, 0,
  0.01918785, 0.02440211, 0.02489228, 0.02704698, 0.01387623, 0.01414828, 
    0.005677442, 0.01708907, 0.004416754, 0.002665421, 0.006203004, 
    0.02122856, 0.03317077, 0.03057763, 0.02803567, 0.009149161, 0.01096385, 
    0.008822633, 0.01226392, 0.001125386, 0.004753313, 0.01353509, 
    0.05223329, 0.02054876, 0.004692578, 0.005303041, 0.009192417, 
    0.00669074, 0.0002207189,
  0.1812336, 0.1607883, 0.1392677, 0.08703392, 0.0904445, 0.0994458, 
    0.04512223, 0.0637292, 0.02150591, 0.02065232, 0.03449914, 0.07864599, 
    0.07742157, 0.02910453, 0.04202192, 0.07601181, 0.1156458, 0.1383469, 
    0.1118508, 0.1320118, 0.09873316, 0.118915, 0.1188025, 0.03802615, 
    0.06512456, 0.06374689, 0.08951533, 0.1690214, 0.1469931,
  0.1487703, 0.08958329, 0.08410607, 0.08354159, 0.07970731, 0.1013334, 
    0.07693079, 0.09340353, 0.06749208, 0.03970537, 0.07093022, 0.06423866, 
    0.0631834, 0.07547529, 0.04717014, 0.1346391, 0.1363659, 0.1030257, 
    0.1288904, 0.1224245, 0.1805641, 0.2384673, 0.1360001, 0.1103498, 
    0.1042604, 0.1532692, 0.1729096, 0.1663494, 0.1774546,
  0.01832039, 0.008791882, 0.0006923647, 0.002930682, 0.01405212, 0.03521011, 
    0.0003143586, 0.0004792812, 0.01401142, 0.04522121, 0.1079053, 0.1232202, 
    0.05267657, 0.05111029, 0.1116454, 0.1454486, 0.08245847, 0.1050613, 
    0.1798034, 0.1976319, 0.05339517, 0.02579765, 0.05729472, 0.01911764, 
    0.06804883, 0.0583817, 0.1118989, 0.03821305, 0.01231557,
  2.90299e-07, 3.082301e-07, 3.499046e-07, 6.814874e-08, 0.0006691797, 
    -0.0008356005, -7.259349e-07, -1.283415e-06, 0.00778123, 0.00115585, 
    0.003369269, -1.85971e-06, -4.457464e-05, 8.17511e-06, 0.06080177, 
    0.08143008, 0.05887813, 0.03865362, 0.02378196, 0.01924367, 
    -2.003994e-06, 4.118057e-08, 3.258068e-08, 0.0005652234, 0.0003280249, 
    0.007107735, 2.082084e-06, -8.30818e-06, -8.092994e-08,
  2.423142e-06, 6.861188e-08, 2.543788e-06, -6.64121e-05, 0.01466132, 
    0.03314694, 0.01679222, 0.04620869, 0.03718717, 0.05474501, 8.830284e-06, 
    -0.0001264617, 0.07492079, 0.107884, 0.06331456, 0.1288501, 0.06548344, 
    0.0006801619, 0.0001126197, 9.674687e-05, 4.215339e-08, 4.743103e-07, 
    0.003422592, 0.002142409, -4.865189e-05, -2.622112e-05, -2.564148e-08, 
    9.407126e-06, 3.727205e-06,
  0.01672837, 0.02719884, 0.03093651, 0.0005451423, 0.0005973718, 0.04917635, 
    0.07668614, 0.02584258, 0.1225392, 0.0982236, 0.02269655, 0.04784717, 
    0.1978765, 0.05895859, 0.08013573, 0.009149849, 0.001744081, 0.01753357, 
    4.294462e-06, 0.0009597876, -2.642448e-05, 0.01202125, 0.09663912, 
    0.1912678, 0.05825118, 0.00880952, 0.004106802, 5.045014e-05, 0.002127069,
  0.09387533, 0.06140851, 0.06247677, -4.39289e-05, 0.02738424, 0.0610679, 
    0.133069, 0.1099588, 0.1883475, 0.0606681, 0.02636638, 0.05614214, 
    0.2100305, 0.1445804, 0.1022926, 0.09548175, 0.09845583, 0.01187118, 
    0.01580816, 0.01462494, 0.08665292, 0.2147659, 0.2483104, 0.113405, 
    0.07077063, 0.03113387, 0.01606234, 0.1543158, 0.1174005,
  0.01829275, 0.003378053, -7.954943e-05, 0.0006171247, 0.01504813, 
    0.1005575, 0.1299718, 0.1698145, 0.1385529, 0.1569247, 0.1094161, 
    0.06886172, 0.09256238, 0.03939084, 0.03134544, 0.01868121, 0.01213305, 
    0.01071448, 0.04651356, 0.0009009992, 0.012232, 0.09588651, 0.09555002, 
    0.1397244, 0.03200977, 0.008745351, 0.001011999, 0.01001779, 0.04736115,
  0.04609993, 0.05900349, 0.007019787, 0.001368918, -3.231994e-05, 
    -8.310237e-06, 0.04912073, 0.09458978, 0.3230389, 0.1267525, 0.2205329, 
    0.1194794, 0.09693523, 0.1027984, 0.1394181, 0.07735024, 0.06589733, 
    0.04112777, 0.03918332, 0.01618391, 0.01787238, 0.08379146, 0.03648042, 
    0.1157718, 0.1200776, 0.05844766, 0.004994385, 0.0004883436, 0.00239152,
  0.09083226, 0.09408938, 0.06556951, 0.09069696, 0.05345805, 0.05341958, 
    0.07280828, 0.1883305, 0.1913793, 0.1662534, 0.1406888, 0.1753123, 
    0.2147302, 0.1795089, 0.1308031, 0.1839562, 0.1887053, 0.140967, 
    0.04769599, 0.03916828, 0.05743204, 0.107977, 0.05545265, 0.06971703, 
    0.08787487, 0.1038346, 0.05972181, 0.08851997, 0.07940159,
  0.08638166, 0.1654109, 0.1179513, 0.09668457, 0.143278, 0.05988332, 
    0.07154624, 0.06434083, 0.1444775, 0.2142046, 0.2384472, 0.3051997, 
    0.1217437, 0.1220182, 0.1676924, 0.2143505, 0.2096897, 0.261437, 
    0.1708775, 0.05787669, 0.1351864, 0.08495945, 0.105006, 0.1250663, 
    0.1645462, 0.1967463, 0.2040124, 0.1383354, 0.178366,
  0.2183426, 0.07425743, 0.1184465, 0.1017885, 0.1228332, 0.137757, 
    0.1389435, 0.07865472, 0.09698468, 0.08099101, 0.1885398, 0.1646795, 
    0.1096594, 0.1880522, 0.1344001, 0.1011709, 0.08344047, 0.1436737, 
    0.1147294, 0.1141197, 0.08116041, 0.08945794, 0.09500017, 0.1351811, 
    0.159264, 0.08931592, 0.1084974, 0.186603, 0.214183,
  0.144173, 0.1772797, 0.1643892, 0.09858765, 0.09324212, 0.09321848, 
    0.07516292, 0.03478792, 0.06514, 0.05117733, 0.1207773, 0.1196385, 
    0.05949602, 0.01664493, 0.04703112, 0.04246524, 0.06735852, 0.09951174, 
    0.1441997, 0.1510589, 0.1626913, 0.0743606, 0.02505952, -0.009581244, 
    0.06293936, 0.0002478668, -9.73711e-05, 0.1234128, 0.1425415,
  0.03721701, 0.06636182, 0.06985556, 0.03690727, 0.0212581, 0.02941937, 
    0.05742958, 0.1135611, 0.1190063, 0.1174356, 0.1170789, 0.07586376, 
    0.02586408, 0.003303163, 0.00313542, -0.0006168921, 0.0002926251, 
    -0.0004185706, 0.013247, 0.02008156, 0.04134339, 0.0721948, 0.04810932, 
    0.02546102, 0.01305771, -0.0001531513, -0.0002691008, 0.0003756092, 
    0.01827938,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.533132e-05, 0, 0, 0, 
    0, 0, -2.927595e-05, 0, 0, 0, 0, 0,
  0, -5.881756e-05, 0.0002241578, 0.0003140645, -6.751414e-06, -0.00020585, 
    0.01519093, 0, 0, -0.0003926768, -2.43698e-05, -4.731964e-05, 
    -0.0003807917, 0.003711261, 0.03277481, 0.01730724, 0.01700931, 
    0.01103192, 0.005495731, 0.008602384, 0.01327905, 0.01286139, 0.02253468, 
    0.01790217, 0.01026744, -6.33511e-05, -0.0001472494, -0.0001387222, 0,
  0.0453824, 0.05816558, 0.1191872, 0.1281506, 0.1228695, 0.09133465, 
    0.1043549, 0.1032153, 0.1032571, 0.03610573, 0.04774814, 0.06650448, 
    0.09113738, 0.1001154, 0.1173966, 0.04730873, 0.02197963, 0.04563685, 
    0.06792538, 0.04935752, 0.09384993, 0.1259859, 0.1255494, 0.06850763, 
    0.04129253, 0.0165406, 0.03046117, 0.02145774, 0.02970869,
  0.196516, 0.1857888, 0.1995453, 0.1695275, 0.1238845, 0.1555567, 0.1354295, 
    0.1274387, 0.07499687, 0.1067335, 0.08858731, 0.1643058, 0.131813, 
    0.09057839, 0.1636637, 0.1460313, 0.1730819, 0.1764046, 0.1862659, 
    0.1896858, 0.1866349, 0.1924412, 0.1543301, 0.06020169, 0.08752155, 
    0.1537017, 0.1542251, 0.2151673, 0.1752843,
  0.1296301, 0.07676627, 0.0692738, 0.08818374, 0.09485441, 0.1083786, 
    0.07587943, 0.09501792, 0.08156133, 0.06306505, 0.1057502, 0.09763359, 
    0.07674622, 0.1203658, 0.09312626, 0.1458188, 0.1477873, 0.1004499, 
    0.1429563, 0.1238935, 0.1716727, 0.2597536, 0.160458, 0.1381303, 
    0.1170833, 0.1667661, 0.159771, 0.1569758, 0.1637862,
  0.01149145, 0.002614508, 0.002034019, 0.002531636, 0.01151244, 0.01351761, 
    0.002616016, 0.001673951, 0.01401536, 0.05796338, 0.09024751, 0.1193787, 
    0.05687108, 0.05234591, 0.1167208, 0.142544, 0.07409377, 0.09963384, 
    0.1631002, 0.1931836, 0.02376538, 0.01680169, 0.05034895, 0.03657833, 
    0.07512948, 0.0605592, 0.09012097, 0.02478925, 0.009249024,
  5.891859e-08, 3.373819e-07, 1.483133e-07, 2.039963e-06, 0.001158018, 
    -0.001027518, 0.00115492, -8.017501e-05, 0.01199315, 0.01020482, 
    0.007604872, 4.138432e-06, -1.780766e-05, 2.734055e-06, 0.05946584, 
    0.07818052, 0.03056345, 0.018831, 0.02057209, 0.01768802, 4.499521e-07, 
    5.028446e-08, 1.783099e-07, 0.002869421, 0.0003270694, 0.0008714129, 
    4.297771e-07, -1.48329e-05, -1.731909e-07,
  1.814447e-06, 2.795472e-08, 4.21145e-06, 0.0009957843, 0.01910406, 
    0.03148644, 0.01665791, 0.03684887, 0.03612916, 0.03952315, 0.0001139054, 
    0.0007956877, 0.06218767, 0.08472715, 0.05267653, 0.1238744, 0.05523413, 
    0.000690292, 9.498583e-05, 7.695475e-07, 6.137632e-09, 1.005651e-07, 
    0.009240428, -0.000141391, 1.629807e-06, -4.825676e-07, -3.818756e-07, 
    1.307968e-05, 3.673606e-06,
  0.01406062, 0.02471435, 0.02002692, 0.003877831, 0.001336623, 0.04148633, 
    0.05827225, 0.01757809, 0.08805411, 0.08577451, 0.01463825, 0.03321735, 
    0.1706745, 0.04439025, 0.06320184, 0.006453898, 0.001178166, 0.01840185, 
    5.94511e-06, 1.934772e-05, 4.234901e-06, 0.000744588, 0.06286174, 
    0.1576962, 0.04678513, 0.03447643, 0.004356534, 0.0004841328, 0.00304014,
  0.06463302, 0.05495944, 0.08008482, -9.248452e-05, 0.01915262, 0.04088319, 
    0.1089963, 0.04982185, 0.1334913, 0.04545787, 0.01598531, 0.03475473, 
    0.1823209, 0.1229771, 0.09850397, 0.06739832, 0.09198629, 0.006826807, 
    0.01614863, 0.01909796, 0.0873963, 0.185737, 0.1965381, 0.0738814, 
    0.06720062, 0.02299964, 0.01590437, 0.1310104, 0.09276915,
  0.01830816, 0.002702333, -3.012124e-05, 0.0003031539, 0.01203161, 
    0.1016924, 0.1257309, 0.1395473, 0.1298941, 0.1468241, 0.0899797, 
    0.0548032, 0.06607955, 0.02522732, 0.02657983, 0.01211485, 0.00390848, 
    0.000245941, 0.04271589, 1.602322e-05, 0.01043798, 0.09178897, 
    0.05232255, 0.1131516, 0.02590171, 0.004776814, 0.0002336112, 
    0.007664031, 0.06284229,
  0.03366467, 0.05361081, 0.01082481, 0.0005119971, -1.186769e-05, 
    -1.926699e-05, 0.03701147, 0.07866365, 0.2902488, 0.1090905, 0.1897373, 
    0.1068169, 0.1052079, 0.08873288, 0.1360708, 0.05402379, 0.03651313, 
    0.02079432, 0.0194483, 0.01231874, 0.00367928, 0.05179093, 0.02550557, 
    0.07867772, 0.1233081, 0.05225149, 0.0005853171, 2.812946e-05, 
    -0.0002737479,
  0.08028736, 0.08978821, 0.05364609, 0.06787521, 0.04768862, 0.05681552, 
    0.11969, 0.1527981, 0.1685779, 0.1429183, 0.1423929, 0.1622069, 
    0.2078926, 0.1688935, 0.1398527, 0.1769366, 0.1574035, 0.1149838, 
    0.03774705, 0.03802687, 0.06109608, 0.1122308, 0.04682774, 0.05597206, 
    0.08076458, 0.09741775, 0.04783255, 0.07727707, 0.06979071,
  0.06215931, 0.1578308, 0.1184646, 0.08067385, 0.1351018, 0.0573195, 
    0.0589854, 0.1115737, 0.191986, 0.2384004, 0.1952625, 0.2883627, 
    0.1030734, 0.1217878, 0.1477029, 0.202145, 0.2246118, 0.2434419, 
    0.1518203, 0.08804233, 0.1349333, 0.06720993, 0.09620976, 0.1177781, 
    0.1546715, 0.190045, 0.1767387, 0.1203838, 0.1530853,
  0.2105161, 0.07982469, 0.1209878, 0.1230618, 0.1212411, 0.1212887, 
    0.1279436, 0.09093048, 0.1191484, 0.1529251, 0.2319167, 0.1974446, 
    0.158759, 0.1803732, 0.1286252, 0.1503597, 0.1157411, 0.221942, 
    0.1585272, 0.1235247, 0.08362662, 0.09357475, 0.1120395, 0.1527506, 
    0.1840342, 0.1180101, 0.1142354, 0.2053677, 0.201851,
  0.232279, 0.2012092, 0.2242967, 0.1060261, 0.1386327, 0.1624779, 
    0.08669462, 0.05893811, 0.1065817, 0.08896678, 0.106379, 0.0929362, 
    0.06422028, 0.05848018, 0.1292616, 0.2198426, 0.1618799, 0.1898717, 
    0.1825928, 0.2069818, 0.2204645, 0.1595164, 0.1246157, 0.05806859, 
    0.0936747, 0.005925831, 0.0005556724, 0.1720767, 0.1883246,
  0.1378148, 0.1601564, 0.0740351, 0.05154834, 0.09585751, 0.2055056, 
    0.2509934, 0.2555715, 0.2382369, 0.2027241, 0.256364, 0.2442382, 
    0.1956242, 0.08753627, 0.1318535, 0.09486183, 0.02301695, 0.009255362, 
    0.02445216, 0.07416078, 0.09044812, 0.09928419, 0.09913296, 0.07154249, 
    0.0534872, 0.003927827, 0.001949843, 0.03840449, 0.1593965,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.439364e-05, 
    -8.82418e-05, 0.0002727489, 7.280989e-06, -1.783056e-06, 0, 7.348985e-05, 
    0.0001687828, 0.0001073174, 0, 0, 0, 0,
  0.001049044, 0.01588891, 0.02069155, 0.008016451, -0.0007861581, 
    -0.002482464, 0.04657708, -0.0005278005, -0.0002613995, -0.001147085, 
    -8.065866e-06, -0.0002728429, 0.0002585777, 0.0279938, 0.04196087, 
    0.03853448, 0.03139282, 0.0132445, 0.03514363, 0.06110639, 0.05989176, 
    0.06939229, 0.1022107, 0.05579712, 0.04152951, 0.0110872, 0.02287417, 
    0.005600124, 0.0001973257,
  0.10075, 0.1293887, 0.1569221, 0.1348637, 0.1379645, 0.1185926, 0.1561479, 
    0.1350762, 0.1495635, 0.1405488, 0.1398538, 0.1495523, 0.1432895, 
    0.1901575, 0.2481519, 0.1081524, 0.1175471, 0.09755411, 0.1377761, 
    0.1533808, 0.1981517, 0.1893235, 0.1918553, 0.1426866, 0.1182797, 
    0.04609243, 0.05701748, 0.09125677, 0.09239803,
  0.2283109, 0.2005151, 0.2288954, 0.1876059, 0.1521426, 0.18254, 0.1501969, 
    0.1302609, 0.1169999, 0.1714703, 0.1620104, 0.2126626, 0.2064411, 
    0.2022814, 0.2121038, 0.21444, 0.2157187, 0.2137836, 0.241694, 0.2385559, 
    0.2287983, 0.2319201, 0.1898249, 0.09798928, 0.1217624, 0.1591616, 
    0.1719379, 0.2426858, 0.190575,
  0.1166807, 0.06026437, 0.06257162, 0.08529052, 0.09182294, 0.09568076, 
    0.06873828, 0.1017522, 0.100439, 0.07186449, 0.1010665, 0.1064187, 
    0.08445124, 0.1169795, 0.1067857, 0.1432454, 0.1339358, 0.1132611, 
    0.1198851, 0.1475351, 0.1660615, 0.2565691, 0.1807502, 0.1488017, 
    0.1160667, 0.1491968, 0.1471554, 0.1369287, 0.1363663,
  0.007685991, 1.173607e-06, 0.006440544, 0.003661713, 0.008491365, 
    0.01130432, 0.001551754, 0.002631112, 0.01196786, 0.03189208, 0.08207176, 
    0.1193665, 0.05992796, 0.05697829, 0.08265882, 0.1544542, 0.0490619, 
    0.08745565, 0.1562201, 0.1880079, 0.008407553, 0.01909175, 0.03047215, 
    0.0387495, 0.0659835, 0.06024159, 0.06546865, 0.02135311, 0.00768935,
  2.727987e-08, 2.127765e-07, 9.268596e-09, 2.846484e-05, 0.0006386629, 
    0.03777464, 0.009558499, 0.004278568, 0.002524219, 0.003692607, 
    0.00453987, 2.979901e-07, -1.991999e-05, -2.151868e-06, 0.06182718, 
    0.07690368, 0.01877518, 0.005326339, 0.016574, 0.0326349, 5.949017e-07, 
    4.347249e-09, 7.849053e-08, 0.008880824, 0.0003366611, 2.587813e-05, 
    9.296577e-07, -3.123075e-06, -9.385892e-05,
  3.151456e-05, 1.069643e-06, 4.763321e-06, 0.006283119, 0.02128329, 
    0.02981011, 0.01981983, 0.03663205, 0.0439401, 0.0337175, 0.0008258459, 
    0.01340167, 0.05583803, 0.08090291, 0.05668063, 0.1141613, 0.04233812, 
    0.001664396, 0.002614661, 1.527382e-08, -2.131091e-08, 1.461594e-07, 
    0.01259663, 0.0002235946, -1.367211e-05, -3.628823e-06, 2.39188e-07, 
    4.287024e-06, 1.777422e-06,
  0.0143385, 0.03509092, 0.01786902, 0.009102635, 0.001417423, 0.03833665, 
    0.03169505, 0.01102921, 0.05481939, 0.06584211, 0.01667793, 0.03278141, 
    0.1490996, 0.05084881, 0.04490078, 0.005763458, 0.006146525, 0.02185578, 
    -6.482597e-05, -6.620781e-06, 1.070589e-06, -7.1959e-05, 0.05564813, 
    0.1398936, 0.04931599, 0.05083708, 0.01585535, 0.002634061, 0.002630553,
  0.04557325, 0.04422817, 0.07937432, -3.521214e-05, 0.01004603, 0.03064289, 
    0.09430913, 0.02615219, 0.1014985, 0.03284366, 0.008439644, 0.02357603, 
    0.1764006, 0.1056697, 0.08445007, 0.05593396, 0.09462674, 0.005059693, 
    0.02233699, 0.01717941, 0.09782553, 0.1782806, 0.1549204, 0.0574083, 
    0.07110619, 0.02509613, 0.01571029, 0.1385399, 0.07014849,
  0.01257536, 0.002427965, -3.28203e-06, -6.602244e-06, 0.003493513, 
    0.1034563, 0.1089021, 0.1090071, 0.09070469, 0.1401591, 0.07914576, 
    0.04405701, 0.04833785, 0.01833567, 0.02739539, 0.01145508, 0.002211061, 
    -2.033684e-05, 0.03232912, 1.280344e-05, 0.005636205, 0.08861644, 
    0.03298313, 0.09390196, 0.01523407, 0.0009157209, 0.0002648481, 
    0.004257743, 0.04914875,
  0.01941199, 0.04917044, 0.01191035, 0.0009959781, -2.676999e-05, 
    -2.927587e-06, 0.02931552, 0.06977125, 0.2860192, 0.1066498, 0.1667338, 
    0.1177273, 0.1008907, 0.04839913, 0.1215233, 0.05061141, 0.04381418, 
    0.004579681, 0.0008034632, 0.007466443, 0.001042301, 0.03024207, 
    0.01900819, 0.04418693, 0.1211657, 0.02322797, 0.0009356607, 
    1.067834e-06, 0.0003886429,
  0.07466318, 0.08202123, 0.03985706, 0.0632979, 0.05480697, 0.05816295, 
    0.1509114, 0.1307937, 0.1512871, 0.1333072, 0.1397653, 0.1403526, 
    0.1947104, 0.157876, 0.1412713, 0.162168, 0.1594218, 0.09154904, 
    0.01758157, 0.02589203, 0.04729993, 0.1239861, 0.03911907, 0.04756311, 
    0.08491785, 0.08768986, 0.03803798, 0.06536518, 0.04947091,
  0.06427762, 0.1368709, 0.1059248, 0.07815698, 0.1050064, 0.04538948, 
    0.05289787, 0.1052558, 0.1932919, 0.2355166, 0.1738649, 0.2669805, 
    0.08760331, 0.1128049, 0.13503, 0.1895186, 0.2307091, 0.2535011, 
    0.1477847, 0.06539717, 0.1375932, 0.05506095, 0.09353821, 0.1014141, 
    0.148524, 0.1857553, 0.1690862, 0.1236616, 0.1593789,
  0.1945221, 0.06153221, 0.1086663, 0.1149405, 0.1004589, 0.1028819, 
    0.1139103, 0.1098979, 0.1818732, 0.1692125, 0.2161945, 0.2112923, 
    0.1644709, 0.1684379, 0.1180031, 0.1461822, 0.1841038, 0.2508066, 
    0.1634412, 0.1103373, 0.08121296, 0.08273071, 0.09878211, 0.1684598, 
    0.1740596, 0.1663672, 0.1236354, 0.2364996, 0.2002717,
  0.2566319, 0.1843139, 0.2203754, 0.1007559, 0.1412945, 0.1719826, 
    0.1102093, 0.08590297, 0.09713686, 0.09628323, 0.1417757, 0.09353728, 
    0.08231565, 0.05869982, 0.1222397, 0.2006067, 0.1869504, 0.2584149, 
    0.183863, 0.1973792, 0.226457, 0.1624317, 0.128028, 0.0855087, 
    0.07380917, 0.04393611, 0.01691703, 0.195043, 0.2160864,
  0.128282, 0.144839, 0.0680118, 0.09682187, 0.1391722, 0.2643203, 0.2843822, 
    0.2842866, 0.22747, 0.196399, 0.2364355, 0.2448429, 0.2449996, 0.1618875, 
    0.2095357, 0.171773, 0.08741651, 0.06329992, 0.09549229, 0.1150659, 
    0.1104325, 0.1242022, 0.1087265, 0.06211307, 0.1215142, 0.02160159, 
    0.03085437, 0.07316318, 0.1583448,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9.157618e-09, -6.694824e-08, 
    -5.577335e-05, -0.0001025184, -0.0001690417, 0.008750577, 0.001309512, 
    0.001564824, 3.266035e-06, 0.003725671, 0.05222247, 0.03698675, 
    0.001952862, 0.001651777, 0.005839238, 0,
  0.02129914, 0.0445413, 0.07335045, 0.03096221, 0.000205867, 0.01201172, 
    0.06770802, 0.0003543109, 0.001185307, 0.00303275, 0.003139404, 
    -0.000625131, 0.01367128, 0.1155659, 0.2071911, 0.1256876, 0.13986, 
    0.08787212, 0.1651862, 0.1525163, 0.1219788, 0.1728572, 0.1891718, 
    0.1079507, 0.1061306, 0.02940326, 0.08228981, 0.1038149, 0.02492889,
  0.1640575, 0.212647, 0.2188775, 0.1782677, 0.1565895, 0.1369383, 0.159021, 
    0.1451069, 0.1820656, 0.2000391, 0.2019767, 0.2069708, 0.2353819, 
    0.2600591, 0.2895248, 0.1985908, 0.180482, 0.186277, 0.2127637, 
    0.2436397, 0.2732679, 0.2257981, 0.2429208, 0.1960772, 0.2032527, 
    0.1039744, 0.1250173, 0.1523017, 0.1587952,
  0.2604707, 0.218397, 0.2446873, 0.1819296, 0.1744196, 0.1889046, 0.1523984, 
    0.1330932, 0.1423499, 0.1761053, 0.1870812, 0.2070484, 0.2079301, 
    0.2225847, 0.2062004, 0.2146689, 0.2595635, 0.2503805, 0.2348618, 
    0.2521072, 0.2667367, 0.2313026, 0.2109801, 0.143973, 0.1373262, 
    0.1842892, 0.219236, 0.2676977, 0.2250939,
  0.1108413, 0.05845527, 0.0647594, 0.08294617, 0.08582673, 0.0791651, 
    0.0671159, 0.1003047, 0.1016567, 0.07606902, 0.1117954, 0.09683039, 
    0.08119369, 0.117884, 0.1096002, 0.1446493, 0.1203943, 0.1119168, 
    0.1290842, 0.1628612, 0.165761, 0.2282612, 0.1909304, 0.1655388, 
    0.09761798, 0.1424427, 0.1410807, 0.1249545, 0.1150096,
  0.005326481, -9.884026e-06, 0.01188456, 0.004664488, 0.01100374, 
    0.01664245, 0.005164925, 0.003539294, 0.008051623, 0.01914548, 
    0.06550838, 0.124364, 0.06333508, 0.06865489, 0.06071768, 0.1580724, 
    0.03360611, 0.07988776, 0.1459991, 0.1703941, 0.009378735, 0.01647059, 
    0.02484553, 0.02537775, 0.05660055, 0.0635342, 0.05311897, 0.02606156, 
    0.003800892,
  9.807265e-09, 7.688585e-08, 1.612163e-09, 0.0002344974, 0.001547144, 
    0.04688881, 0.01245441, 0.0009290863, 0.0126498, 0.001495789, 
    0.003824475, 5.879315e-07, -0.0001464817, -9.648508e-05, 0.06878053, 
    0.07860255, 0.01018722, 0.002272015, 0.01805262, 0.03656897, 
    4.175345e-07, 0, 7.044288e-09, 0.01394267, 0.0003600827, 4.356974e-06, 
    1.269371e-06, 0.000328497, -0.0003290576,
  6.536652e-05, 1.529523e-06, 4.075508e-06, 0.008773422, 0.01958774, 
    0.04825522, 0.02278242, 0.03287425, 0.04881533, 0.02992435, 0.01888038, 
    0.01490677, 0.05058324, 0.08110399, 0.04800683, 0.1022333, 0.05831083, 
    0.004520162, 0.0003896578, 4.3275e-08, -9.545179e-09, 4.007782e-07, 
    0.007084787, 0.002730732, 5.84017e-05, -3.155755e-05, 5.207114e-07, 
    3.073422e-07, 9.818971e-07,
  0.003457096, 0.03661257, 0.01599523, 0.01261342, 0.003668947, 0.03687991, 
    0.02725399, 0.008467495, 0.03202375, 0.06112545, 0.02677727, 0.04322991, 
    0.144717, 0.0428293, 0.03519405, 0.007443742, 0.009368355, 0.01623028, 
    -8.442321e-05, 3.751909e-05, 1.573997e-05, -1.634402e-06, 0.04755302, 
    0.1451625, 0.06833091, 0.07732356, 0.02875304, 0.01705638, 0.0005807584,
  0.0347439, 0.03983825, 0.06223668, -9.533364e-05, 0.002270212, 0.02412639, 
    0.08777934, 0.01984279, 0.07159862, 0.01840064, 0.005739372, 0.02007736, 
    0.1586312, 0.1010946, 0.0818394, 0.05481774, 0.1004945, 0.01500216, 
    0.03201317, 0.02292298, 0.1102636, 0.1756197, 0.1320306, 0.05073122, 
    0.0745051, 0.02218351, 0.01823247, 0.1439761, 0.04922515,
  0.04131656, 0.0017103, -7.103152e-07, 0.000645323, 0.002726186, 0.09073441, 
    0.111288, 0.08620413, 0.0923098, 0.1438293, 0.0664202, 0.03363671, 
    0.03531647, 0.01398982, 0.02506655, 0.01299417, 0.0001460607, 
    1.506027e-05, 0.00671219, 2.276833e-06, 0.003407312, 0.08674594, 
    0.02317022, 0.07643376, 0.00915698, 0.00489044, 0.001837378, 0.006935806, 
    0.04020422,
  0.01006278, 0.05271256, 0.01450139, 0.005476239, -9.721142e-05, 
    0.0007835812, 0.03309697, 0.08708283, 0.2822585, 0.09871237, 0.145493, 
    0.1182555, 0.1053408, 0.04679967, 0.1358889, 0.03423416, 0.03440748, 
    0.0001085407, -1.097807e-05, 0.002997693, 0.002437142, 0.02348703, 
    0.01748496, 0.02781349, 0.1204502, 0.008472994, 0.0001375525, 
    -7.093436e-06, 0.0001166348,
  0.06740093, 0.07673761, 0.03300529, 0.0683932, 0.05878893, 0.03702781, 
    0.1562178, 0.1158958, 0.1409722, 0.1488547, 0.1254712, 0.1127793, 
    0.1751308, 0.1489355, 0.1265427, 0.1712381, 0.1625442, 0.05205843, 
    0.002559377, 0.01836123, 0.04164726, 0.1155488, 0.03315638, 0.0380274, 
    0.0863782, 0.08117694, 0.05261842, 0.05935285, 0.04334211,
  0.06379506, 0.118262, 0.1072953, 0.07084589, 0.09233394, 0.04060256, 
    0.04229433, 0.09286586, 0.1935657, 0.2180704, 0.1717377, 0.2464608, 
    0.07602537, 0.1171925, 0.1385628, 0.1730375, 0.2286845, 0.2577354, 
    0.17096, 0.0525067, 0.1361888, 0.04899322, 0.08880711, 0.08733913, 
    0.1411154, 0.1922895, 0.1545973, 0.1320225, 0.1694009,
  0.1683299, 0.04262168, 0.09515207, 0.1122286, 0.09882967, 0.0942799, 
    0.09893144, 0.0930407, 0.1875581, 0.1686738, 0.2015089, 0.2098381, 
    0.1611944, 0.1572755, 0.107131, 0.1434928, 0.1862562, 0.270494, 
    0.1552689, 0.08894982, 0.07281487, 0.07092328, 0.08878018, 0.1656188, 
    0.1672439, 0.2057408, 0.1307093, 0.2577755, 0.2111006,
  0.2519172, 0.168457, 0.2193039, 0.08110087, 0.1427581, 0.1699404, 
    0.1078098, 0.1251045, 0.07783913, 0.09739001, 0.1552747, 0.09450214, 
    0.07884756, 0.03716063, 0.1082528, 0.1658464, 0.1702152, 0.2374035, 
    0.1796252, 0.1833752, 0.2110209, 0.1531352, 0.1355769, 0.09819183, 
    0.04743879, 0.1466659, 0.08315911, 0.1773267, 0.2440168,
  0.1208402, 0.1261977, 0.06471946, 0.1297736, 0.1768298, 0.285394, 
    0.2712857, 0.2669772, 0.2087665, 0.1741053, 0.1891232, 0.2326374, 
    0.2455967, 0.1862724, 0.2192494, 0.1842403, 0.0954484, 0.07220551, 
    0.1236611, 0.1221563, 0.117722, 0.1244802, 0.104837, 0.05477544, 
    0.1035352, 0.05186414, 0.08475622, 0.07601308, 0.1498452,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.003427406, 0.01918685, 0.02625854, 
    0.04833312, 0.01492764, 0.01784475, 0.004682666, 0.004650822, 
    0.001582552, 0.01410729, 0.1106602, 0.120233, 0.03554815, 0.03928156, 
    0.01010505, 0,
  0.04744544, 0.1554267, 0.1367793, 0.08688159, 0.009326582, 0.03620252, 
    0.09108499, 0.01870036, 0.006391956, 0.01689873, 0.007647778, 
    -0.002274456, 0.06150845, 0.2473687, 0.2142124, 0.1520118, 0.1629101, 
    0.1878073, 0.2016896, 0.2222956, 0.2444451, 0.2740478, 0.2229304, 
    0.1603774, 0.2007168, 0.1078063, 0.151557, 0.1222104, 0.04712905,
  0.1962938, 0.267028, 0.2761231, 0.2654516, 0.244268, 0.1752873, 0.1841713, 
    0.1742371, 0.2086612, 0.2900464, 0.2507991, 0.263919, 0.262317, 
    0.2609819, 0.2851969, 0.2005326, 0.1912121, 0.2083944, 0.2207654, 
    0.2197676, 0.2652311, 0.2239443, 0.2325867, 0.2053274, 0.2397897, 
    0.1945113, 0.2119181, 0.1732002, 0.2039997,
  0.2636239, 0.2097575, 0.2462402, 0.1705109, 0.1739197, 0.1750648, 
    0.1591008, 0.1434765, 0.1533936, 0.1781904, 0.2075086, 0.2077321, 
    0.1949016, 0.2141651, 0.2025587, 0.2082171, 0.2573629, 0.2529139, 
    0.2578204, 0.2367807, 0.2277495, 0.2348105, 0.2137414, 0.1645433, 
    0.1544812, 0.1784648, 0.2488685, 0.2851644, 0.2549941,
  0.09653812, 0.07382119, 0.05855655, 0.07613599, 0.08499125, 0.07612823, 
    0.06915444, 0.08934073, 0.09044575, 0.07658879, 0.1170818, 0.0867932, 
    0.08198623, 0.1179149, 0.110126, 0.1258301, 0.1344998, 0.1094875, 
    0.1195187, 0.1646751, 0.1579611, 0.1930014, 0.1793948, 0.1945893, 
    0.08165331, 0.1404597, 0.125556, 0.1137922, 0.1062172,
  0.003413785, 9.269629e-05, 0.01429547, 0.005871884, 0.01262975, 0.02161508, 
    0.005108002, 0.003539755, 0.009726723, 0.01715056, 0.05196343, 0.1079635, 
    0.06849671, 0.05790246, 0.04749652, 0.1541762, 0.04448768, 0.06725474, 
    0.1434472, 0.1710979, 0.01653038, 0.01767689, 0.0208106, 0.0204784, 
    0.05318819, 0.05940104, 0.03834351, 0.03062331, 0.001088451,
  -8.060756e-09, 3.914461e-08, -9.461821e-10, 3.552778e-06, 0.006512217, 
    0.04107044, 0.0064126, 2.27836e-05, 0.01588773, 0.006476462, 0.01119166, 
    -1.939896e-06, -0.0003470945, 0.0001114896, 0.07167944, 0.07439329, 
    0.01385496, 0.00202746, 0.009151366, 0.04243026, 1.568718e-08, 
    1.062621e-13, -4.071511e-10, 0.03402491, 0.000312885, 4.434635e-06, 
    2.518216e-06, 0.001372141, 0.005388546,
  1.974955e-05, -4.988407e-07, 2.965354e-05, 0.009908656, 0.01814768, 
    0.06251109, 0.02303665, 0.02905128, 0.04946265, 0.03255317, 0.03262328, 
    0.01341895, 0.04526621, 0.08413807, 0.05379485, 0.1125523, 0.08124465, 
    0.007545423, 0.0005027674, 9.471648e-08, 1.030643e-08, 6.056084e-07, 
    0.0003859581, 0.00332774, 4.471173e-05, 0.001313606, -5.34727e-07, 
    7.119553e-08, 4.779085e-07,
  0.001502428, 0.04580343, 0.0167571, 0.02224239, 0.003707462, 0.03053983, 
    0.0240189, 0.006927163, 0.02570052, 0.06351051, 0.0242861, 0.04135346, 
    0.1243895, 0.04566279, 0.03342531, 0.007560718, 0.004234074, 0.01425808, 
    0.004414769, 0.000324108, 4.401957e-05, -2.216405e-06, 0.0479249, 
    0.1495622, 0.09872435, 0.08238495, 0.03901044, 0.002713646, 0.0003550353,
  0.03188706, 0.04671968, 0.04620546, 0.001496159, 0.00164439, 0.01551976, 
    0.08856563, 0.02180966, 0.04810062, 0.0206017, 0.005189962, 0.01663557, 
    0.1517941, 0.09878407, 0.06743269, 0.05624712, 0.1044705, 0.03692075, 
    0.04243048, 0.02899768, 0.1104002, 0.1723464, 0.1177258, 0.05525623, 
    0.06145686, 0.03047649, 0.02487233, 0.1384213, 0.04799464,
  0.05369797, 0.008279272, -6.541164e-07, 1.368448e-05, 0.0002362451, 
    0.07169477, 0.1247151, 0.09000936, 0.09416562, 0.137995, 0.05878627, 
    0.02869292, 0.03029402, 0.00820672, 0.01484592, 0.01681034, 2.869188e-05, 
    1.498817e-06, 0.02074938, -5.658697e-06, 0.006162343, 0.08984084, 
    0.01596923, 0.06241717, 0.007186914, 0.01914814, 0.01377039, 0.003184773, 
    0.03344229,
  0.005900461, 0.06226392, 0.01951686, 0.01545888, -0.0002215696, 
    0.006011008, 0.0195435, 0.09745291, 0.2722369, 0.07507603, 0.1304239, 
    0.1216475, 0.1111526, 0.04505643, 0.1317395, 0.02371506, 0.01629468, 
    4.691212e-05, 0.0003076806, 0.001645594, 0.007972173, 0.02972949, 
    0.01486228, 0.0189243, 0.100833, 0.00858382, -8.577124e-07, 1.362016e-07, 
    0.00085385,
  0.0638314, 0.07484135, 0.02709161, 0.07006533, 0.0530203, 0.01852836, 
    0.1537166, 0.1028142, 0.1351568, 0.1701122, 0.1156286, 0.09717345, 
    0.1562441, 0.149467, 0.1157192, 0.1810511, 0.1448675, 0.03130023, 
    0.004480116, 0.009408658, 0.05071842, 0.09696113, 0.03357064, 0.03288537, 
    0.09187831, 0.06958748, 0.03562401, 0.06160329, 0.03363999,
  0.05185831, 0.09469669, 0.108802, 0.06463888, 0.08592145, 0.03357072, 
    0.04405441, 0.09903419, 0.186735, 0.2145888, 0.1749732, 0.2167451, 
    0.07335459, 0.1203715, 0.1383516, 0.1709699, 0.2105357, 0.2441058, 
    0.1399196, 0.04800291, 0.138938, 0.04695486, 0.08631986, 0.07425819, 
    0.1394311, 0.1885677, 0.1408898, 0.1175939, 0.1558073,
  0.1608363, 0.03544682, 0.07438341, 0.1029521, 0.09401948, 0.08864897, 
    0.09505377, 0.0792046, 0.1789685, 0.1840928, 0.1934087, 0.1982753, 
    0.1556118, 0.1280526, 0.0857537, 0.1480678, 0.1933412, 0.299178, 
    0.1466328, 0.08240582, 0.06643574, 0.05805599, 0.09233103, 0.1779329, 
    0.1761049, 0.2414788, 0.1563026, 0.2575231, 0.2037476,
  0.2475516, 0.1681351, 0.2211449, 0.07523225, 0.1337001, 0.1801528, 
    0.1104028, 0.1393462, 0.06337851, 0.1011881, 0.1459413, 0.09508403, 
    0.0873017, 0.0329328, 0.1131425, 0.1404224, 0.1509114, 0.2188124, 
    0.177361, 0.1818351, 0.1931161, 0.1362602, 0.1373234, 0.1094971, 
    0.04562412, 0.2171277, 0.1361428, 0.17266, 0.2375309,
  0.1211432, 0.1279135, 0.05948556, 0.163807, 0.1859566, 0.3087847, 
    0.3073098, 0.2667111, 0.1927617, 0.168796, 0.1833732, 0.2272759, 
    0.2291875, 0.1859691, 0.2175367, 0.1823893, 0.09468018, 0.0780937, 
    0.1451289, 0.1336432, 0.1289914, 0.122648, 0.1042777, 0.05899908, 
    0.09245335, 0.07717481, 0.09961901, 0.07300454, 0.1614805,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01957734, 0.05339067, 0.1027235, 
    0.1105623, 0.09353364, 0.06032145, 0.03135996, 0.009888103, 0.008965865, 
    0.07528188, 0.2039551, 0.2418415, 0.160809, 0.09813417, 0.03245788, 
    0.0001993931,
  0.08699787, 0.2513617, 0.2941843, 0.2180031, 0.0380582, 0.07256581, 
    0.1594979, 0.05117589, 0.02251754, 0.05067247, 0.04415363, 0.03327441, 
    0.1510613, 0.2855705, 0.2226509, 0.1422199, 0.1795634, 0.2523272, 
    0.2610077, 0.3267585, 0.3439788, 0.3125626, 0.2264184, 0.281042, 
    0.2600639, 0.1516228, 0.1835988, 0.1621578, 0.102231,
  0.2151287, 0.3219078, 0.2847305, 0.2842907, 0.3024635, 0.227027, 0.2315203, 
    0.2089641, 0.2441271, 0.3414122, 0.2712601, 0.2682524, 0.2493814, 
    0.2474822, 0.2726561, 0.2178204, 0.21456, 0.2235013, 0.2293395, 
    0.1995194, 0.2739439, 0.2547491, 0.2681023, 0.2325256, 0.2723869, 
    0.2420268, 0.2632541, 0.2137985, 0.226296,
  0.249124, 0.1996295, 0.2363057, 0.1624294, 0.1693243, 0.1617754, 0.1641588, 
    0.1541716, 0.1464656, 0.1990071, 0.2086636, 0.1960063, 0.1626608, 
    0.203933, 0.1958469, 0.1536821, 0.2553135, 0.2426815, 0.2353028, 
    0.2314541, 0.2505935, 0.2335992, 0.1800674, 0.1632318, 0.141702, 
    0.2138214, 0.2562372, 0.3036312, 0.2485634,
  0.09029854, 0.07893422, 0.05811946, 0.07271644, 0.08438671, 0.07814474, 
    0.07107021, 0.0905164, 0.07333551, 0.05689306, 0.1085378, 0.09029212, 
    0.0897436, 0.1023657, 0.09983756, 0.1112145, 0.120839, 0.1118263, 
    0.1005119, 0.1657001, 0.1534422, 0.1747819, 0.1795772, 0.2146724, 
    0.07630204, 0.1232374, 0.1178845, 0.102234, 0.1026717,
  0.005741696, 0.000638128, 0.01436098, 0.009153281, 0.02060972, 0.02204055, 
    0.004807215, 0.004986329, 0.01832587, 0.01931956, 0.04086564, 0.09948285, 
    0.05611781, 0.0408665, 0.03526095, 0.1539805, 0.03674188, 0.0562925, 
    0.1309343, 0.1789969, 0.03232932, 0.01517118, 0.02013926, 0.02802913, 
    0.04602655, 0.05856593, 0.04046813, 0.03000147, 0.002974856,
  -2.652946e-09, 2.864929e-09, -5.178586e-10, 1.262981e-05, 0.02923048, 
    0.04363438, 0.006375057, 1.537075e-05, 0.009950031, 0.007282892, 
    0.01494902, 2.61832e-07, 0.001363244, 0.003365621, 0.04037287, 
    0.07290297, 0.02892759, 0.001333505, 0.005998847, 0.04729705, 
    2.036664e-09, 3.022316e-08, 4.098291e-09, 0.03698684, 0.0002749814, 
    5.845949e-06, 3.137432e-07, 0.000409819, 0.008316849,
  1.199634e-05, 1.324964e-07, 3.712259e-05, 0.01180607, 0.01840873, 
    0.0611081, 0.02570897, 0.03559704, 0.0426389, 0.03132079, 0.03881971, 
    0.01450523, 0.05488415, 0.08248031, 0.05726361, 0.1326709, 0.09318005, 
    0.00435982, 0.0005649471, -1.038178e-06, 9.600555e-08, 1.501634e-06, 
    8.401894e-06, 0.0009285482, 3.522313e-05, 2.159676e-05, -6.97643e-09, 
    2.217006e-07, 5.018848e-07,
  0.008043179, 0.03774877, 0.02272068, 0.02895267, 0.004294347, 0.01545628, 
    0.02615662, 0.005009906, 0.02411886, 0.06443853, 0.02851265, 0.05376676, 
    0.114648, 0.08938768, 0.03468695, 0.008901122, 0.004894529, 0.009994647, 
    0.02391934, 0.0002587552, 2.735515e-05, 1.067979e-05, 0.05518369, 
    0.1410307, 0.1104441, 0.06537441, 0.04925435, 0.006073391, 0.002708133,
  0.03632467, 0.03942063, 0.03848013, 0.03159361, 0.004140864, 0.009410287, 
    0.1012083, 0.02214669, 0.03571795, 0.02799615, 0.005785954, 0.01941125, 
    0.1462301, 0.1106486, 0.07230937, 0.05911924, 0.09270493, 0.03897611, 
    0.0625003, 0.03436748, 0.121265, 0.1749621, 0.1137363, 0.07156032, 
    0.07075813, 0.0326547, 0.04208594, 0.1269333, 0.04715568,
  0.08129042, 0.02973686, -3.987802e-05, 2.151813e-06, -3.523137e-07, 
    0.04829698, 0.1689973, 0.1369745, 0.1222998, 0.1551117, 0.06132729, 
    0.02522938, 0.03203922, 0.004976673, 0.01113668, 0.01262789, 
    9.318835e-05, 3.281466e-05, 0.02879275, -2.341192e-05, 0.01121696, 
    0.09776668, 0.01353122, 0.05763097, 0.006201462, 0.01875127, 0.004270105, 
    5.514998e-05, 0.02019713,
  0.003766789, 0.05497219, 0.0064724, 0.008816903, 0.000113884, 0.001570444, 
    0.02483147, 0.09665823, 0.2684526, 0.06216275, 0.1253687, 0.1311439, 
    0.1077381, 0.05155789, 0.1374353, 0.01348336, 0.007196776, 0.0001194377, 
    1.478322e-05, 0.0005608493, 0.0122664, 0.02172984, 0.00944712, 
    0.01638396, 0.0932323, 0.01140442, 2.89943e-06, 8.207709e-08, 0.000843714,
  0.06713006, 0.07631458, 0.02591264, 0.07528546, 0.04039978, 0.01696823, 
    0.164513, 0.09375581, 0.1215603, 0.1763578, 0.1059304, 0.08401697, 
    0.1439992, 0.1433375, 0.1107224, 0.1705655, 0.1283772, 0.03443501, 
    0.002489821, 0.004420727, 0.06116607, 0.08458745, 0.03801523, 0.0334082, 
    0.09190697, 0.06647673, 0.04355589, 0.04265668, 0.03002816,
  0.02895798, 0.1100341, 0.118647, 0.06470273, 0.09329478, 0.0374819, 
    0.05955678, 0.1026255, 0.1807108, 0.2135874, 0.1560274, 0.1956311, 
    0.08062717, 0.1270519, 0.1451108, 0.1657971, 0.2182331, 0.2448295, 
    0.1401717, 0.04889141, 0.1453543, 0.05198281, 0.08661496, 0.07069295, 
    0.142199, 0.1856577, 0.1437963, 0.112512, 0.1228495,
  0.1713292, 0.05936938, 0.0590095, 0.1018691, 0.09786251, 0.08844238, 
    0.1002376, 0.08766686, 0.1797414, 0.1966745, 0.1789214, 0.2015871, 
    0.1590213, 0.1121714, 0.0741666, 0.166686, 0.2101722, 0.3371561, 
    0.1464765, 0.08737165, 0.06756385, 0.06062144, 0.09917694, 0.1861697, 
    0.1708939, 0.2458779, 0.1870434, 0.2990197, 0.2263758,
  0.2746735, 0.177095, 0.25713, 0.0831501, 0.1305842, 0.2256193, 0.1380712, 
    0.1543785, 0.06116566, 0.1187705, 0.1404508, 0.1205378, 0.1024887, 
    0.0610132, 0.1012025, 0.1253655, 0.1379051, 0.1965253, 0.1699769, 
    0.1788421, 0.1920608, 0.1449199, 0.1455692, 0.1294531, 0.04643923, 
    0.2166475, 0.2593017, 0.1768477, 0.225728,
  0.1451894, 0.1465662, 0.0647079, 0.1638421, 0.1801556, 0.314093, 0.2811657, 
    0.2252948, 0.1748557, 0.1463231, 0.2082946, 0.2323214, 0.2299144, 
    0.194231, 0.2166689, 0.1667732, 0.08666192, 0.07574239, 0.159303, 
    0.153639, 0.1434457, 0.1239489, 0.11028, 0.06188318, 0.08697413, 
    0.07912996, 0.08718811, 0.0880857, 0.2144677,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0002076328, -0.0001904485, 
    -0.0001732641, -0.0001560798, -0.0001388954, -0.0001217111, 
    -0.0001045267, 5.756757e-05, 4.038322e-05, 2.319887e-05, 6.014522e-06, 
    -1.116983e-05, -2.835418e-05, -4.553852e-05, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3.384607e-07, 0.07229615, 0.1539227, 
    0.1875242, 0.1541281, 0.1414418, 0.1283234, 0.06527811, 0.04284469, 
    0.04360433, 0.128022, 0.2540832, 0.3059874, 0.231399, 0.2057099, 
    0.04675732, 0.001767912,
  0.09915364, 0.2930616, 0.3110733, 0.3331235, 0.06959631, 0.1096855, 
    0.2278472, 0.08628528, 0.07361934, 0.083391, 0.09155999, 0.1037614, 
    0.2017808, 0.2756905, 0.193603, 0.1217174, 0.1766403, 0.2632951, 
    0.2730659, 0.3219894, 0.3725983, 0.3135026, 0.2562424, 0.2921426, 
    0.2806134, 0.1849516, 0.1866467, 0.2331477, 0.1540878,
  0.2164353, 0.3482307, 0.2702564, 0.287707, 0.3066658, 0.2396927, 0.2436365, 
    0.2410612, 0.2474353, 0.3409863, 0.2829734, 0.2561132, 0.2495628, 
    0.2434659, 0.2609321, 0.2085688, 0.2248258, 0.248277, 0.2611818, 
    0.1984639, 0.2479465, 0.2330364, 0.2648684, 0.2214895, 0.2756464, 
    0.2447999, 0.2583765, 0.2161842, 0.2088137,
  0.2446016, 0.1902419, 0.2201106, 0.1383809, 0.1559595, 0.1488183, 
    0.1756199, 0.1716556, 0.14235, 0.1880543, 0.2008711, 0.1962913, 
    0.1609572, 0.2058439, 0.1916529, 0.1896798, 0.248228, 0.212892, 
    0.2175129, 0.2576547, 0.209067, 0.2399213, 0.179629, 0.1553962, 0.130155, 
    0.1818093, 0.2470453, 0.294474, 0.2536161,
  0.0789335, 0.08844125, 0.06996025, 0.09398192, 0.09856407, 0.07675778, 
    0.06902581, 0.08561771, 0.08546933, 0.06059103, 0.1206015, 0.08886675, 
    0.08797892, 0.09153953, 0.1079842, 0.106513, 0.1119411, 0.09429238, 
    0.09592193, 0.1513716, 0.1384418, 0.1639936, 0.1833616, 0.2313785, 
    0.07247715, 0.1104151, 0.1162867, 0.0964165, 0.1040549,
  0.00530152, 0.001515644, 0.02076058, 0.01776746, 0.03051688, 0.02200395, 
    0.005460567, 0.01032276, 0.02605681, 0.02921421, 0.02845064, 0.09386513, 
    0.05891557, 0.03465453, 0.03086941, 0.1650759, 0.02713296, 0.05653788, 
    0.1208788, 0.195232, 0.04951189, 0.01790236, 0.0205138, 0.02490526, 
    0.03910583, 0.07297628, 0.04254516, 0.02832807, 0.009975545,
  1.311991e-07, 1.906832e-08, 1.646186e-08, 0.0001875227, 0.0517914, 
    0.05255828, 0.00148358, 0.000343549, 0.006630346, 0.005043788, 
    0.01731364, -0.0001124531, 0.003974246, 0.004192703, 0.03024866, 
    0.05898518, 0.04544663, 0.003378624, 0.006174483, 0.05183859, 
    2.093554e-08, 9.985101e-08, 8.843639e-08, 0.02818511, 0.0003376948, 
    9.647786e-06, 9.780416e-07, 0.0008580352, 0.01386274,
  5.202396e-06, 4.123097e-07, 2.039202e-06, 0.02416762, 0.03432383, 
    0.05555359, 0.03274995, 0.04102373, 0.05183141, 0.03338071, 0.03946124, 
    0.03643697, 0.06772263, 0.103903, 0.07960109, 0.1431413, 0.1156922, 
    0.01020294, 0.002278366, -3.356443e-06, 4.138776e-07, 2.265893e-06, 
    0.0004680688, 0.001792711, 4.382551e-05, -9.765516e-06, 3.092569e-07, 
    1.128894e-06, 2.389686e-06,
  0.02998986, 0.0422594, 0.03784789, 0.03184456, 0.002319591, 0.01267525, 
    0.03566662, 0.006303741, 0.03223846, 0.06997856, 0.05033507, 0.06673206, 
    0.1296456, 0.1235006, 0.0376181, 0.008833401, 0.004595785, 0.005970701, 
    0.02033658, 0.001042431, 0.006768947, 0.0003436997, 0.04832897, 
    0.1651854, 0.1242765, 0.0607171, 0.059837, 0.01773041, 0.007466604,
  0.04169026, 0.02637631, 0.01708851, 0.1896613, 0.003668722, 0.01721375, 
    0.1079642, 0.02743021, 0.04275331, 0.04142696, 0.01504666, 0.02432685, 
    0.1722786, 0.1254268, 0.08577613, 0.06699289, 0.08597314, 0.04981662, 
    0.07802719, 0.03547608, 0.1293224, 0.1880862, 0.1237586, 0.08646222, 
    0.09179329, 0.05088919, 0.06012294, 0.1527437, 0.05841351,
  0.05179107, 0.03160699, 0.0001398245, 3.196059e-06, 4.387257e-06, 
    0.01231142, 0.1864378, 0.1859739, 0.1908754, 0.1887382, 0.07709645, 
    0.02799399, 0.04608109, 0.006127952, 0.01588848, 0.007964571, 
    0.0007170443, 0.0004034989, 0.03095925, 2.852881e-05, 0.01182535, 
    0.1132806, 0.01930494, 0.05535042, 0.007133943, 0.02148158, 0.002517312, 
    0.0001247779, 0.01647816,
  0.003394112, 0.05585711, 0.005719048, 0.004839433, -0.0001831529, 
    0.0001390233, 0.02536994, 0.1135574, 0.2453628, 0.06171125, 0.1294683, 
    0.1562158, 0.1054406, 0.0545066, 0.1424367, 0.01047645, 0.007436451, 
    0.0002625968, 4.026569e-06, 0.0001776682, 0.01517771, 0.02006051, 
    0.009879477, 0.01840012, 0.08430872, 0.01186589, 2.864589e-06, 
    7.68243e-08, 0.002030685,
  0.06827747, 0.07122043, 0.02815474, 0.08087282, 0.02536823, 0.01052112, 
    0.1562467, 0.08504938, 0.1049865, 0.1595193, 0.1026096, 0.07305096, 
    0.1412161, 0.1435853, 0.107755, 0.1742739, 0.1159538, 0.03591204, 
    0.01080819, 0.004526891, 0.05959388, 0.07241111, 0.04432123, 0.04870041, 
    0.09048758, 0.06686839, 0.04296567, 0.03348689, 0.03477351,
  0.03098314, 0.09447421, 0.1366811, 0.072673, 0.08728127, 0.03546359, 
    0.0617708, 0.106914, 0.1857054, 0.2184886, 0.1563167, 0.1991485, 
    0.09714106, 0.1384727, 0.155463, 0.1712878, 0.2118765, 0.2263965, 
    0.1541726, 0.04751728, 0.1509194, 0.05908357, 0.09019765, 0.07283682, 
    0.1512996, 0.1846527, 0.1480792, 0.1112234, 0.1263721,
  0.1706285, 0.05433755, 0.06448653, 0.09831741, 0.1158708, 0.119986, 
    0.1094096, 0.104217, 0.1836056, 0.1979571, 0.1712593, 0.2151505, 
    0.1604165, 0.1062428, 0.09484109, 0.1680702, 0.2230815, 0.3586902, 
    0.1316059, 0.09390757, 0.1009349, 0.05405535, 0.1083424, 0.1836778, 
    0.1736551, 0.2703768, 0.2293557, 0.3028042, 0.218068,
  0.2339213, 0.1691618, 0.2476031, 0.08947465, 0.1634133, 0.2479726, 
    0.1753391, 0.1576996, 0.05459663, 0.1284186, 0.1259191, 0.1596714, 
    0.1135594, 0.09153943, 0.0907122, 0.1247037, 0.137796, 0.1916284, 
    0.1575373, 0.1795433, 0.1916351, 0.1397793, 0.1636349, 0.1289703, 
    0.02653265, 0.2140478, 0.3008373, 0.1675196, 0.2401617,
  0.1303367, 0.1604551, 0.1033194, 0.1989861, 0.2159798, 0.3147539, 
    0.3034173, 0.2522606, 0.1986734, 0.2029441, 0.1943441, 0.2078679, 
    0.2341606, 0.2131628, 0.2291146, 0.1656245, 0.105496, 0.1128514, 
    0.1706546, 0.1816334, 0.1537162, 0.1302605, 0.1231185, 0.06995168, 
    0.08211315, 0.08037927, 0.09086021, 0.1412484, 0.1796092,
  0, 0, 0, 0, 0, 0, 0, -0.0001520815, -0.0001005284, -4.89754e-05, 
    2.577652e-06, 5.41307e-05, 0.0001056838, 0.0001572368, -0.0007332514, 
    -0.000716067, -0.0006988827, -0.0006816983, -0.000664514, -0.0006473296, 
    -0.0006301453, 0.0002302703, 0.0001615329, 9.279548e-05, 2.405809e-05, 
    -4.467931e-05, -0.0001134167, -0.0001821541, 0,
  -0.002399456, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0.000627482, 0.0001893941, 
    0.0001545213, 0.1405375, 0.2029918, 0.227357, 0.2210037, 0.1965712, 
    0.2233836, 0.136943, 0.08480222, 0.09730329, 0.1787517, 0.2503303, 
    0.291209, 0.2824224, 0.3323669, 0.1139661, 0.01997199,
  0.09516176, 0.2806457, 0.3234039, 0.3775795, 0.1182854, 0.1225247, 
    0.2988472, 0.1122137, 0.08191728, 0.1383883, 0.1310664, 0.1564349, 
    0.2331283, 0.3000558, 0.1882955, 0.1181603, 0.1735862, 0.2685413, 
    0.3189738, 0.3666337, 0.3511944, 0.3513002, 0.2447375, 0.3094628, 
    0.2851561, 0.1786165, 0.1676475, 0.2128959, 0.1402577,
  0.2414749, 0.375118, 0.289039, 0.305314, 0.3161747, 0.2370827, 0.2407729, 
    0.2253928, 0.2478506, 0.3433802, 0.2936331, 0.2443113, 0.2405672, 
    0.2101984, 0.2497453, 0.1923372, 0.2216592, 0.2616267, 0.2754572, 
    0.1772071, 0.2202812, 0.2115871, 0.2609883, 0.2318321, 0.2925238, 
    0.2203868, 0.2569766, 0.2069237, 0.2025501,
  0.2623154, 0.1938601, 0.2219876, 0.1286767, 0.1570385, 0.1466203, 
    0.1740892, 0.1564496, 0.1270679, 0.1636551, 0.2032535, 0.1924637, 
    0.1707099, 0.2011596, 0.1728975, 0.1943327, 0.2398937, 0.2028841, 
    0.217549, 0.2018247, 0.1977774, 0.2342965, 0.1950128, 0.1485894, 
    0.1363213, 0.1833112, 0.224553, 0.2845939, 0.2640847,
  0.07810917, 0.0968326, 0.08297592, 0.1100086, 0.1107249, 0.08174314, 
    0.06826517, 0.08722188, 0.08153638, 0.06127432, 0.1525511, 0.1106622, 
    0.08958354, 0.09985524, 0.1320304, 0.1037623, 0.103955, 0.08287756, 
    0.09328847, 0.1254548, 0.1218593, 0.1434198, 0.1815727, 0.2375274, 
    0.0743636, 0.1108246, 0.11345, 0.0939322, 0.08732741,
  0.004756622, 0.001662398, 0.03095433, 0.02723506, 0.03879293, 0.03440012, 
    0.006729418, 0.0193026, 0.03152465, 0.02901073, 0.0297158, 0.07300168, 
    0.05175187, 0.03963945, 0.03535159, 0.1643302, 0.0372155, 0.05698349, 
    0.12509, 0.2028961, 0.08299183, 0.01997897, 0.02142772, 0.01541615, 
    0.03838108, 0.09808885, 0.06494686, 0.03409427, 0.005801992,
  1.876541e-07, 7.621502e-08, 9.062598e-08, -5.44769e-05, 0.08764791, 
    0.05938022, 0.001002059, 0.01977401, 0.004384797, 0.007783421, 
    0.02387924, 0.001010866, 0.001904252, 0.008257267, 0.03086663, 
    0.05847103, 0.05682627, 0.008675565, 0.01382298, 0.0477429, 3.052188e-07, 
    2.655891e-07, 1.228714e-07, 0.004098387, 0.003878761, 5.043011e-05, 
    1.121915e-05, 0.001041993, 0.01856709,
  4.364768e-06, 5.245856e-07, 1.238949e-05, 0.02679794, 0.04816601, 
    0.06132578, 0.0267153, 0.04153338, 0.07459322, 0.04675483, 0.0384112, 
    0.03770329, 0.08903047, 0.1237892, 0.09073343, 0.162718, 0.1322963, 
    0.01023621, 0.003513715, 2.761763e-07, 8.164433e-08, 1.176858e-06, 
    0.0007266115, 0.004804695, 5.399224e-05, -1.284913e-05, -2.470763e-06, 
    0.0001403037, -7.072982e-06,
  0.04030081, 0.0574836, 0.08288451, 0.02939295, 0.001726972, 0.01422824, 
    0.03982369, 0.006093375, 0.04878668, 0.07427765, 0.04187608, 0.07062184, 
    0.1588704, 0.1185089, 0.04755088, 0.007759098, 0.004961884, 0.007617434, 
    0.01480426, 0.003447108, 0.009258867, 0.001778439, 0.05269961, 0.2162371, 
    0.1257773, 0.06658798, 0.0747372, 0.01883359, 0.01227321,
  0.0461197, 0.01974023, 0.01131047, 0.3056267, 0.002709573, 0.0375502, 
    0.1127601, 0.03036832, 0.05192721, 0.04114672, 0.02375423, 0.02554074, 
    0.1878272, 0.1329695, 0.08595432, 0.06271225, 0.0989193, 0.05755639, 
    0.06986725, 0.03743589, 0.1301007, 0.18966, 0.1492935, 0.1036524, 
    0.110292, 0.07221585, 0.07948047, 0.1779157, 0.06267731,
  0.03342248, 0.01842947, 4.029964e-07, 7.190432e-07, 4.640372e-06, 
    0.0004949067, 0.2178678, 0.1548152, 0.2444963, 0.2255315, 0.08279324, 
    0.03671934, 0.05540176, 0.006063418, 0.02309419, 0.005392903, 
    0.001878966, 6.187945e-05, 0.01660098, 0.0003377495, 0.01482427, 
    0.1267563, 0.02152036, 0.05001873, 0.007227309, 0.01994887, 0.002785702, 
    0.0001835609, 0.0274439,
  0.001046569, 0.05688038, 0.001563534, 0.0006228289, -8.811346e-05, 
    -0.0001628503, 0.01931211, 0.1130558, 0.2334724, 0.06159882, 0.1378455, 
    0.1270047, 0.1266108, 0.06292997, 0.1580731, 0.0081891, 0.01565091, 
    0.0007256138, 1.537084e-06, 1.044362e-05, 0.007853069, 0.01948761, 
    0.01194968, 0.03416166, 0.09329168, 0.01558991, 1.534564e-05, 
    2.005191e-07, 0.0001513067,
  0.07814825, 0.05501318, 0.03337304, 0.08850075, 0.01901294, 0.006953508, 
    0.1339814, 0.0848223, 0.0843745, 0.122262, 0.09939294, 0.07627784, 
    0.1475263, 0.1457767, 0.1057696, 0.1950401, 0.1019197, 0.0377733, 
    0.01581833, 0.003800458, 0.04293005, 0.07307095, 0.05443802, 0.07874348, 
    0.1078517, 0.07588057, 0.05274332, 0.02728066, 0.03269562,
  0.04673333, 0.09655873, 0.1491975, 0.07527044, 0.09747791, 0.04115627, 
    0.05567599, 0.1193414, 0.1850593, 0.2169434, 0.1576388, 0.1771926, 
    0.09480982, 0.1552452, 0.1930866, 0.1747955, 0.213702, 0.2126934, 
    0.1771263, 0.04432802, 0.1454425, 0.08470723, 0.1039915, 0.07637874, 
    0.1576545, 0.1805036, 0.1552133, 0.09201179, 0.1332447,
  0.157221, 0.04875446, 0.05607307, 0.1352534, 0.1397705, 0.1676967, 
    0.09818941, 0.09917564, 0.1785273, 0.1887808, 0.1515812, 0.2309079, 
    0.195062, 0.1247351, 0.151464, 0.1487316, 0.269385, 0.3936819, 0.1484723, 
    0.09843963, 0.0890775, 0.04837371, 0.1127021, 0.2361815, 0.2311837, 
    0.2748567, 0.214549, 0.263961, 0.2008351,
  0.2317775, 0.1755223, 0.2768641, 0.07324916, 0.1282574, 0.2191809, 
    0.1376487, 0.1441468, 0.05474504, 0.1528854, 0.1235557, 0.1824593, 
    0.09315777, 0.08580164, 0.0946338, 0.1090656, 0.1305397, 0.1727096, 
    0.1558177, 0.1713648, 0.1810513, 0.1312888, 0.1874228, 0.1403486, 
    0.02396564, 0.2166482, 0.3086347, 0.1717887, 0.1902447,
  0.1048561, 0.1374608, 0.08397399, 0.2158551, 0.2283541, 0.2736352, 
    0.2038537, 0.1806745, 0.1566739, 0.2181274, 0.1716987, 0.1489419, 
    0.1939663, 0.2199948, 0.2559079, 0.1966382, 0.1871141, 0.1781597, 
    0.1966428, 0.2633973, 0.2209997, 0.1540319, 0.132652, 0.07439505, 
    0.07219002, 0.08583944, 0.09563753, 0.09675012, 0.1676486,
  1.073616e-06, 3.451996e-07, -3.832167e-07, -1.111633e-06, -1.840049e-06, 
    -2.568466e-06, -3.296882e-06, -0.000396291, -0.0002619551, -0.0001276191, 
    6.716796e-06, 0.0001410527, 0.0002753887, 0.0004097246, -0.00146676, 
    -0.001413742, -0.001360723, -0.001307705, -0.001254686, -0.001201667, 
    -0.001148649, 0.0006195023, 0.0004328762, 0.0002462501, 5.962398e-05, 
    -0.0001270021, -0.0003136282, -0.0005002543, 1.656349e-06,
  -0.001885479, 0, 0, 0, 0, -0.001188064, -0.0006400249, -4.095932e-05, 
    -2.86697e-07, 0.0007820179, 0.007757294, 0.00128632, 0.001778025, 
    0.2138546, 0.2525131, 0.2411417, 0.236584, 0.2507591, 0.245698, 
    0.2309809, 0.1774597, 0.1279112, 0.2143135, 0.2501971, 0.2682345, 
    0.2831326, 0.3384607, 0.2567548, 0.02554368,
  0.09940236, 0.2806365, 0.3290215, 0.3760012, 0.1768969, 0.137624, 
    0.3271847, 0.1554583, 0.1228925, 0.1784145, 0.1790813, 0.1985606, 
    0.247659, 0.3215277, 0.1908071, 0.128393, 0.1941564, 0.3359739, 
    0.3130789, 0.3806522, 0.3487926, 0.3718315, 0.264428, 0.3067146, 
    0.2827775, 0.1558134, 0.1618003, 0.2023593, 0.1047048,
  0.2553449, 0.3749503, 0.3406177, 0.3244691, 0.3320907, 0.2334655, 
    0.2518884, 0.2448423, 0.2530573, 0.3327615, 0.3064686, 0.2430409, 
    0.2692682, 0.2274164, 0.2648521, 0.1943707, 0.1886279, 0.2880988, 
    0.2564662, 0.1714637, 0.2280726, 0.2065185, 0.2811767, 0.2395983, 
    0.2866477, 0.2029706, 0.2458957, 0.1701772, 0.1769534,
  0.2543844, 0.1894121, 0.2111821, 0.130827, 0.1646151, 0.1432139, 0.1613183, 
    0.1661026, 0.136619, 0.1862327, 0.2222997, 0.2134947, 0.1754533, 
    0.1955461, 0.1695216, 0.1512786, 0.225881, 0.1951326, 0.2034649, 
    0.1982821, 0.1725518, 0.2654159, 0.1837202, 0.1455812, 0.1395846, 
    0.1705115, 0.207655, 0.277792, 0.261455,
  0.08220888, 0.1044309, 0.08504143, 0.1190399, 0.1069547, 0.08207636, 
    0.06173727, 0.08197526, 0.09726001, 0.07716495, 0.1748946, 0.1312928, 
    0.09832656, 0.1045785, 0.1219757, 0.09828756, 0.1047459, 0.08382498, 
    0.07959475, 0.1002196, 0.128047, 0.1367864, 0.174908, 0.2377575, 
    0.07373713, 0.1051242, 0.1275113, 0.09324706, 0.09166192,
  0.004543365, 0.0024976, 0.04019395, 0.03442019, 0.04900768, 0.03640497, 
    0.007695418, 0.02074838, 0.0384121, 0.03627258, 0.05701844, 0.06159585, 
    0.04425879, 0.04592316, 0.04568618, 0.1521677, 0.05415474, 0.06007, 
    0.1315835, 0.2117113, 0.09223556, 0.01790575, 0.02216224, 0.003664106, 
    0.03840266, 0.1239281, 0.06931461, 0.03681312, 0.01122174,
  2.622109e-07, 4.385736e-08, -2.076441e-07, -8.230085e-05, 0.08500407, 
    0.03811005, 0.000369396, 0.04179081, 0.002812999, 0.02304691, 0.01876877, 
    0.002203395, 0.003209499, 0.00662136, 0.03125249, 0.04272424, 0.05565199, 
    0.01885508, 0.04712031, 0.05776727, 3.427225e-07, 9.71623e-08, 
    1.709007e-08, 4.164725e-05, 0.006783021, 0.0001927688, 6.013189e-05, 
    0.005130157, 0.002715573,
  -7.569913e-06, -1.458663e-05, 2.772605e-05, 0.028278, 0.05553442, 
    0.05562782, 0.02086566, 0.03888592, 0.07768245, 0.03378256, 0.03604624, 
    0.03330004, 0.08661956, 0.1114926, 0.08190967, 0.1542293, 0.1318385, 
    0.01988102, 0.005467666, -4.613107e-08, 2.034076e-06, 5.332748e-07, 
    0.0006117102, 0.007153138, 8.273607e-05, 5.655877e-06, 4.616262e-05, 
    0.001178744, 5.506779e-05,
  0.03937594, 0.06758819, 0.08801721, 0.02744455, 0.001720335, 0.0119712, 
    0.02988616, 0.006026092, 0.05149886, 0.07675256, 0.04013542, 0.05750147, 
    0.1378488, 0.1025594, 0.03647721, 0.008623788, 0.004010383, 0.006961239, 
    0.01939629, 0.004946487, 0.0115525, 0.0178183, 0.04338906, 0.2526004, 
    0.1400207, 0.06737245, 0.06783436, 0.01192421, 0.01863574,
  0.0402518, 0.01441364, 0.008908042, 0.2237403, 0.002809216, 0.02307322, 
    0.1085847, 0.02523722, 0.01927096, 0.03032629, 0.01561965, 0.01666633, 
    0.149012, 0.1101203, 0.064195, 0.04466423, 0.07535578, 0.06480028, 
    0.06680884, 0.04533199, 0.1230325, 0.1605797, 0.1505154, 0.1019402, 
    0.1002439, 0.0800985, 0.07287451, 0.1457312, 0.07691991,
  0.03155439, 0.003364034, -7.445082e-08, 1.047824e-07, 1.108012e-05, 
    -7.548445e-06, 0.192451, 0.1060853, 0.2427722, 0.1744068, 0.06288169, 
    0.02677085, 0.03820089, 0.00804057, 0.02657458, 0.008477157, 
    0.0009353888, -0.0001833248, 0.002278549, 0.0005462253, 0.008626241, 
    0.1115624, 0.01784503, 0.03593173, 0.0065973, 0.01490534, 0.0001134899, 
    0.000157766, 0.03148615,
  0.000582176, 0.02899704, 6.184913e-05, 2.569938e-05, -2.919525e-05, 
    -2.982694e-05, 0.01579935, 0.1416861, 0.2370194, 0.05939293, 0.1272276, 
    0.09896646, 0.1381652, 0.06021081, 0.17018, 0.01921365, 0.01669563, 
    0.001188872, 7.878045e-08, 8.241483e-07, 0.003827856, 0.01469639, 
    0.01411458, 0.04985968, 0.09079722, 0.01676439, 3.182025e-05, 
    5.976748e-07, -7.2829e-05,
  0.104435, 0.05827417, 0.04527321, 0.09245973, 0.01677668, 0.007660961, 
    0.1022632, 0.08121994, 0.05481988, 0.1023617, 0.1074265, 0.08139954, 
    0.1375629, 0.1606385, 0.1101592, 0.202026, 0.1127392, 0.05017687, 
    0.02027817, 0.004635331, 0.03064056, 0.07702274, 0.05724027, 0.07656287, 
    0.107622, 0.08305145, 0.07600735, 0.02684152, 0.05373296,
  0.04987571, 0.09248815, 0.1501538, 0.08165363, 0.07969486, 0.03614869, 
    0.07367686, 0.130635, 0.1760533, 0.2273399, 0.1604161, 0.18167, 
    0.1212618, 0.156911, 0.2179781, 0.1807683, 0.2158052, 0.2294219, 
    0.2019155, 0.06483738, 0.1477218, 0.109924, 0.114666, 0.08718729, 
    0.1767945, 0.2109959, 0.1640676, 0.09296552, 0.1473996,
  0.1687658, 0.05698774, 0.05330845, 0.1337739, 0.1583489, 0.1332495, 
    0.1006197, 0.1519331, 0.2033398, 0.2130608, 0.1733449, 0.2761471, 
    0.1994706, 0.172315, 0.1312318, 0.1418497, 0.2622942, 0.4015745, 
    0.1573697, 0.1035576, 0.09832101, 0.064014, 0.1265167, 0.2438417, 
    0.2262338, 0.2737256, 0.2510804, 0.3055101, 0.2333849,
  0.2863089, 0.1764677, 0.2821629, 0.1134579, 0.1799037, 0.2415227, 
    0.2176344, 0.1261326, 0.05082284, 0.1308073, 0.12658, 0.2174087, 
    0.2121534, 0.1339357, 0.08605658, 0.1822167, 0.1805651, 0.1495105, 
    0.1561221, 0.1633772, 0.1891843, 0.1320058, 0.153796, 0.1359402, 
    0.03377733, 0.2125798, 0.3078461, 0.1713992, 0.206536,
  0.2467178, 0.149712, 0.09893916, 0.2275235, 0.2601919, 0.2592954, 
    0.2112578, 0.1674842, 0.1841043, 0.2573501, 0.1465877, 0.1453796, 
    0.1949628, 0.3482991, 0.2629239, 0.2041599, 0.2654932, 0.3350136, 
    0.2615465, 0.2763431, 0.2791483, 0.1973719, 0.1770471, 0.1061403, 
    0.0694892, 0.08651394, 0.09127951, 0.1861719, 0.3271025,
  0.001102697, 0.0006314904, 0.0001602839, -0.0003109227, -0.0007821292, 
    -0.001253336, -0.001724542, -0.0008706916, -0.0005506236, -0.0002305557, 
    8.951226e-05, 0.0004095802, 0.0007296482, 0.001049716, 0.0003496778, 
    0.0003369878, 0.0003242978, 0.0003116078, 0.0002989178, 0.0002862278, 
    0.0002735378, -0.001661488, -0.001497659, -0.001333831, -0.001170002, 
    -0.001006173, -0.0008423447, -0.0006785161, 0.001479662,
  0.02886408, -0.00110208, -3.412964e-06, 0, -0.0004833642, 0.004137062, 
    0.006563833, -0.003181461, 0.0008520506, 0.01532496, 0.01388039, 
    0.000774711, 0.006686518, 0.2397414, 0.2689336, 0.2337568, 0.21539, 
    0.2829637, 0.2633848, 0.2728951, 0.2807566, 0.20494, 0.2135196, 
    0.2503512, 0.2404281, 0.2153329, 0.3349659, 0.2763996, 0.05745925,
  0.09823687, 0.311952, 0.3646562, 0.3627278, 0.2582774, 0.1719217, 
    0.3803124, 0.2955314, 0.2048396, 0.2022478, 0.2036028, 0.2298777, 
    0.2426437, 0.3468256, 0.2020003, 0.1253182, 0.1857999, 0.3208202, 
    0.3464205, 0.405629, 0.3525767, 0.3884647, 0.3236974, 0.2879684, 
    0.2734287, 0.1275942, 0.1412254, 0.2087988, 0.08621819,
  0.2762009, 0.3611242, 0.3445421, 0.3226625, 0.3419547, 0.2360346, 
    0.2950505, 0.2571689, 0.2825001, 0.374425, 0.2906935, 0.2417978, 
    0.2882564, 0.1921286, 0.2409845, 0.1619475, 0.2453206, 0.2664298, 
    0.2700131, 0.1826712, 0.2459972, 0.2595679, 0.2724577, 0.2167768, 
    0.263618, 0.233452, 0.2755682, 0.1790642, 0.201205,
  0.2570302, 0.1943877, 0.2608548, 0.1519873, 0.1907425, 0.1509238, 
    0.1845303, 0.1719927, 0.1606205, 0.198682, 0.2258141, 0.2203456, 
    0.1940128, 0.1835752, 0.169199, 0.1811035, 0.2117497, 0.2162242, 
    0.1955887, 0.1786487, 0.1530911, 0.2393818, 0.17257, 0.1513564, 
    0.1484535, 0.1672223, 0.211221, 0.2565099, 0.2747683,
  0.09980989, 0.1260164, 0.09319177, 0.1245853, 0.1153568, 0.09397326, 
    0.07096858, 0.0858012, 0.1036117, 0.09617665, 0.1715046, 0.1352473, 
    0.1132472, 0.1197714, 0.1230641, 0.1055453, 0.1149073, 0.08320718, 
    0.07799161, 0.08414948, 0.1395764, 0.1280011, 0.1746663, 0.2356725, 
    0.07668894, 0.1107252, 0.1490998, 0.09978505, 0.1107373,
  0.009646239, 0.004051952, 0.04908285, 0.04088812, 0.04414976, 0.04427921, 
    0.01967392, 0.02448382, 0.04513015, 0.05125561, 0.06135954, 0.07721559, 
    0.03979708, 0.05193303, 0.06172014, 0.1550084, 0.05676644, 0.06674422, 
    0.1518385, 0.2206851, 0.1100118, 0.02728416, 0.03198294, 0.002125345, 
    0.04498291, 0.1345459, 0.07894328, 0.04312278, 0.02123417,
  1.354128e-07, -4.732363e-07, -1.476404e-05, 0.00535422, 0.06525682, 
    0.03051826, 0.0006664506, 0.0563339, 0.001753133, 0.02462189, 0.00957683, 
    0.0008647652, 0.01186511, 0.01309705, 0.03219328, 0.03130422, 0.05783222, 
    0.02453229, 0.08681503, 0.0818578, 1.514241e-07, -6.692785e-08, 
    -6.813864e-07, 1.83094e-05, 0.01238961, 0.0001477928, 0.009693959, 
    0.007635626, 0.003121558,
  1.390455e-07, -2.850104e-05, 7.021031e-05, 0.03055304, 0.05642496, 
    0.05732073, 0.01885112, 0.04093605, 0.07493786, 0.02605926, 0.04238902, 
    0.03860429, 0.08908817, 0.09035441, 0.07043362, 0.1404812, 0.142915, 
    0.03047225, 0.008649504, 4.233234e-05, 2.812458e-06, 2.844628e-07, 
    0.0001313762, 0.009313041, 0.0003939566, 0.0002297747, 0.003612216, 
    0.001326449, 8.254978e-07,
  0.0205661, 0.04312524, 0.07217599, 0.02469978, 0.001780349, 0.01202381, 
    0.02299024, 0.005419947, 0.03704923, 0.06512773, 0.03700832, 0.04456367, 
    0.1181671, 0.1031196, 0.03107549, 0.009273682, 0.004596585, 0.00226798, 
    0.01121855, 0.007702276, 0.0007645618, 0.002758994, 0.02606336, 
    0.2499114, 0.1615971, 0.07019773, 0.0742996, 0.005455143, 0.008663866,
  0.03377933, 0.01338207, 0.007641723, 0.1376987, 0.006177548, 0.01112046, 
    0.1084288, 0.02334589, 0.007825398, 0.02671252, 0.01313046, 0.01589379, 
    0.1307085, 0.087014, 0.05483328, 0.04119457, 0.05761297, 0.06157835, 
    0.06900521, 0.05748844, 0.1095468, 0.1230856, 0.1228787, 0.09727547, 
    0.08629889, 0.074733, 0.06328402, 0.122217, 0.05129224,
  0.0171023, 0.0001101783, -2.134694e-08, 2.939735e-08, 7.688962e-06, 
    1.458554e-06, 0.1799278, 0.1034232, 0.2009524, 0.1627412, 0.05533079, 
    0.01748304, 0.02673754, 0.008011243, 0.02644291, 0.009949999, 
    0.001529292, 2.666571e-05, 7.772946e-05, 0.0007933461, 0.003469112, 
    0.1069253, 0.01607139, 0.01562905, 0.009608733, 0.002725321, 
    4.968057e-05, 4.591353e-05, 0.01270208,
  0.0005745117, 0.003962611, 1.036417e-05, 3.450314e-06, -3.908869e-05, 
    -1.751528e-06, 0.01253784, 0.1757237, 0.2563137, 0.05625075, 0.1092232, 
    0.09690212, 0.1348849, 0.06127237, 0.1519284, 0.02014943, 0.01632605, 
    0.003838907, 4.478638e-07, 5.334808e-07, 9.783626e-05, 0.01202889, 
    0.01609348, 0.03767677, 0.07966457, 0.01334852, 0.0001120004, 
    3.11043e-07, 2.03226e-05,
  0.1106458, 0.06012327, 0.05293804, 0.09883122, 0.006798273, 0.003595081, 
    0.07595704, 0.0734093, 0.03256037, 0.09973543, 0.1110255, 0.08319497, 
    0.1476571, 0.1463677, 0.1173093, 0.1872557, 0.1214287, 0.05965415, 
    0.01396828, 0.008780839, 0.02276561, 0.07942197, 0.06538414, 0.07332741, 
    0.106315, 0.08706642, 0.06369451, 0.02720429, 0.05465341,
  0.04926331, 0.09207933, 0.1523919, 0.07211935, 0.07174484, 0.0464414, 
    0.05632707, 0.1178475, 0.1830275, 0.2114093, 0.1744412, 0.210703, 
    0.1230466, 0.1587578, 0.2095855, 0.2049747, 0.2395606, 0.2468928, 
    0.2087057, 0.08226757, 0.1649303, 0.1264435, 0.1327902, 0.09711345, 
    0.1797818, 0.2379941, 0.1558277, 0.1196769, 0.1670397,
  0.1651497, 0.06766623, 0.0784495, 0.1428505, 0.1649694, 0.1425546, 
    0.1118939, 0.139032, 0.2433148, 0.2366079, 0.1888802, 0.3158838, 
    0.2333187, 0.2059788, 0.1393665, 0.1526044, 0.2628476, 0.439156, 
    0.1900814, 0.1131354, 0.1142052, 0.09629367, 0.1450312, 0.2484633, 
    0.1908341, 0.2788397, 0.2598821, 0.2953184, 0.2192834,
  0.2488392, 0.1620289, 0.2494819, 0.08875987, 0.203603, 0.2493408, 
    0.1763372, 0.1244521, 0.09351321, 0.1494057, 0.09626506, 0.194909, 
    0.1396679, 0.1213342, 0.1473727, 0.1757702, 0.165039, 0.1433239, 
    0.1424415, 0.1605485, 0.188594, 0.1245217, 0.193021, 0.1984888, 
    0.03750742, 0.1879321, 0.2939898, 0.1500298, 0.2410396,
  0.2093433, 0.2110491, 0.1692535, 0.2315708, 0.2145741, 0.2426608, 
    0.2068862, 0.1916458, 0.1608169, 0.183235, 0.1147902, 0.09596936, 
    0.1892469, 0.2396058, 0.2503429, 0.2307456, 0.2230172, 0.2709738, 
    0.2782393, 0.2776349, 0.2178046, 0.1827092, 0.2077589, 0.1278137, 
    0.0888145, 0.1122108, 0.1413511, 0.169015, 0.280649,
  0.02229615, 0.01872572, 0.0151553, 0.01158488, 0.008014461, 0.004444039, 
    0.0008736185, 0.0005508244, 0.00121712, 0.001883415, 0.002549711, 
    0.003216006, 0.003882302, 0.004548597, 0.007115309, 0.01055621, 
    0.0139971, 0.017438, 0.0208789, 0.0243198, 0.02776069, 0.04325485, 
    0.04271808, 0.04218131, 0.04164454, 0.04110777, 0.04057099, 0.04003422, 
    0.02515248,
  0.06581829, 0.005058833, -5.244686e-06, -0.0001014923, 0.009027805, 
    0.02322088, 0.0345391, 0.03584521, 0.007723213, 0.02882788, 0.0121361, 
    0.02212896, 0.01282944, 0.2516128, 0.2750846, 0.2401304, 0.2186826, 
    0.2847738, 0.2780157, 0.2731688, 0.3145744, 0.2674514, 0.1934617, 
    0.2441025, 0.2219325, 0.2032826, 0.3136546, 0.2610307, 0.1226692,
  0.1012288, 0.2833502, 0.3798004, 0.3749551, 0.3009212, 0.1892095, 
    0.4293288, 0.4215917, 0.3009977, 0.2086471, 0.2344824, 0.2631609, 
    0.2390266, 0.3981673, 0.2322895, 0.1617782, 0.208415, 0.2924258, 
    0.3538206, 0.4053291, 0.3628311, 0.3360126, 0.314697, 0.3525562, 
    0.2483004, 0.08258387, 0.1467731, 0.1813215, 0.06365997,
  0.317007, 0.4388932, 0.4128437, 0.3142305, 0.3800298, 0.3391646, 0.3334227, 
    0.2608963, 0.2949865, 0.3423353, 0.2817055, 0.2527655, 0.2716635, 
    0.2341187, 0.2959911, 0.2436257, 0.2562864, 0.2744783, 0.2671062, 
    0.2367672, 0.2963539, 0.238586, 0.2792451, 0.2005086, 0.2893498, 
    0.2517257, 0.2730208, 0.1773978, 0.2057403,
  0.2715959, 0.2315484, 0.2805378, 0.1759716, 0.2181139, 0.1502701, 
    0.1891183, 0.1777636, 0.1811559, 0.2032827, 0.2378556, 0.2102159, 
    0.2077491, 0.1739142, 0.1779347, 0.1971909, 0.2488113, 0.2187777, 
    0.2008058, 0.1914722, 0.1649431, 0.2466626, 0.1970824, 0.1496727, 
    0.1498827, 0.160947, 0.2034567, 0.2550105, 0.2645377,
  0.1373785, 0.1444697, 0.1201141, 0.1395016, 0.1331029, 0.1050939, 
    0.09568903, 0.09572767, 0.1224731, 0.1072526, 0.1959249, 0.1414174, 
    0.140774, 0.1352335, 0.1448001, 0.1062069, 0.1438294, 0.08487443, 
    0.09338792, 0.08262329, 0.1686685, 0.1282304, 0.1809656, 0.2478776, 
    0.08803238, 0.1220744, 0.1656544, 0.1073211, 0.1390156,
  0.02424335, 0.00771239, 0.06962154, 0.04647714, 0.04025852, 0.05230182, 
    0.02742204, 0.03784838, 0.05565998, 0.05025681, 0.06169958, 0.07239499, 
    0.05241989, 0.06173921, 0.08613394, 0.1774707, 0.06020057, 0.07904667, 
    0.1760681, 0.2219256, 0.1223303, 0.02701668, 0.05582115, 0.0026777, 
    0.06176626, 0.160288, 0.08946056, 0.04890341, 0.03256553,
  6.652789e-08, -8.086387e-06, 0.0009561553, 0.01132859, 0.07238061, 
    0.02106275, 0.00118763, 0.08324717, 0.005847793, 0.02737137, 0.006742984, 
    -0.000215842, 0.01358557, 0.01777012, 0.05697339, 0.01412454, 0.06003049, 
    0.03651824, 0.1060562, 0.113264, 0.0001446964, -6.566834e-06, 
    1.489108e-05, 1.800517e-05, 0.02678114, 0.001112226, 0.03741344, 
    0.01483593, 0.01127605,
  1.704827e-07, -1.085576e-05, 0.0002202879, 0.08275411, 0.06592903, 
    0.06672081, 0.02264555, 0.04422982, 0.077521, 0.02085268, 0.05035763, 
    0.04872532, 0.102293, 0.08662229, 0.0619842, 0.128332, 0.1538457, 
    0.03569141, 0.01790682, -2.071016e-05, 1.631518e-06, 3.475887e-08, 
    7.986347e-06, 0.01139694, 0.001021963, 0.01087235, 0.008867711, 
    0.001580436, 4.393532e-07,
  0.009296214, 0.046406, 0.07435331, 0.02167203, 0.002379763, 0.01071503, 
    0.01749014, 0.005387233, 0.03024854, 0.06295963, 0.04020598, 0.03407343, 
    0.1051688, 0.09568672, 0.02951393, 0.0130776, 0.008865397, 0.006835727, 
    0.008168534, 0.003582048, 0.000169985, 0.001754582, 0.03199419, 
    0.2807709, 0.1892045, 0.06321475, 0.07958905, 0.000597264, 0.004952291,
  0.03022708, 0.006088242, 0.005424568, 0.06395307, 0.003850287, 0.009030494, 
    0.1019848, 0.02275681, 0.005978962, 0.02196337, 0.01341436, 0.01974496, 
    0.1191908, 0.07340196, 0.05062822, 0.03957524, 0.05461459, 0.05885946, 
    0.07047844, 0.06133579, 0.1019296, 0.1038726, 0.1149754, 0.09259987, 
    0.08090171, 0.08071554, 0.0532865, 0.1084794, 0.0422219,
  0.002230498, 2.890083e-05, -1.244706e-09, 2.974511e-08, 1.792257e-06, 
    -4.226304e-07, 0.1581628, 0.108911, 0.1978735, 0.1577687, 0.05894142, 
    0.0162349, 0.02450257, 0.01384809, 0.02644584, 0.02239247, 0.001069715, 
    0.0001935314, 1.175986e-06, 0.0008123321, 0.001424819, 0.09814086, 
    0.01491423, 0.01287247, 0.01649763, 0.004595951, 1.203693e-05, 
    7.933212e-06, 0.01259836,
  0.0005603239, 0.0001347973, 3.285257e-06, 1.329672e-06, -2.506302e-05, 
    -2.554992e-07, 0.009816841, 0.1856931, 0.2632958, 0.06547974, 0.1052821, 
    0.1029753, 0.1092018, 0.06210998, 0.1191671, 0.01654842, 0.01510281, 
    0.01219039, 4.019156e-07, 2.186808e-07, -0.0001389035, 0.01298152, 
    0.02329817, 0.0378588, 0.07841485, 0.01320567, 0.0003496825, 
    1.127586e-05, 0.0004614256,
  0.09974658, 0.05766266, 0.05714011, 0.09641329, 0.001094888, 0.0004147149, 
    0.06132272, 0.05974552, 0.02396475, 0.09839261, 0.0994812, 0.06775969, 
    0.1419852, 0.1288904, 0.1005475, 0.1831496, 0.1441397, 0.0948262, 
    0.008286227, 0.02024354, 0.01380703, 0.07104541, 0.07560433, 0.06702881, 
    0.0969633, 0.1047968, 0.06684345, 0.03617719, 0.05539157,
  0.06656916, 0.1305155, 0.2059752, 0.07257447, 0.08406461, 0.02981666, 
    0.05433568, 0.1185404, 0.1823592, 0.2021481, 0.1824032, 0.2155509, 
    0.1380822, 0.1897213, 0.2268084, 0.2017127, 0.24968, 0.2579289, 
    0.2233005, 0.1016848, 0.1664597, 0.1305684, 0.1355493, 0.1158897, 
    0.2019785, 0.2550879, 0.1612529, 0.1474443, 0.1943953,
  0.1746361, 0.08034822, 0.09631061, 0.168279, 0.1984944, 0.1730545, 
    0.1109736, 0.1290447, 0.21529, 0.2333165, 0.2514961, 0.33213, 0.2969475, 
    0.1984186, 0.1652717, 0.2027707, 0.3065054, 0.4866659, 0.1957092, 
    0.1195121, 0.1285322, 0.1068002, 0.164304, 0.2806078, 0.2145881, 
    0.2792681, 0.2615418, 0.3157389, 0.2278021,
  0.2903611, 0.2331122, 0.2651592, 0.1201772, 0.1921141, 0.2577505, 
    0.2364667, 0.1576968, 0.1892861, 0.2196087, 0.09688155, 0.1929111, 
    0.1163063, 0.1177556, 0.1455839, 0.1689001, 0.1433922, 0.1385894, 
    0.1539773, 0.1639777, 0.198068, 0.1412685, 0.1752223, 0.2424413, 
    0.0765293, 0.1734727, 0.2725388, 0.1867299, 0.292999,
  0.2188802, 0.2174258, 0.1175306, 0.240475, 0.2343079, 0.3234921, 0.227101, 
    0.1740538, 0.1790977, 0.1788973, 0.1265823, 0.1848705, 0.2663559, 
    0.275908, 0.2852454, 0.2727811, 0.2848451, 0.2881988, 0.3545557, 
    0.3009441, 0.2702033, 0.1984243, 0.2008009, 0.1297484, 0.1504158, 
    0.1434899, 0.190757, 0.1736346, 0.2530115,
  0.07222524, 0.06773897, 0.0632527, 0.05876643, 0.05428017, 0.0497939, 
    0.04530763, 0.04859346, 0.04946177, 0.05033009, 0.0511984, 0.05206672, 
    0.05293503, 0.05380335, 0.04499644, 0.04908443, 0.05317242, 0.05726041, 
    0.0613484, 0.06543639, 0.06952438, 0.0795265, 0.07905646, 0.07858643, 
    0.07811639, 0.07764636, 0.07717633, 0.0767063, 0.07581425,
  0.1017247, 0.04196965, -0.001940764, 0.002687033, 0.01350909, 0.02857641, 
    0.05530962, 0.06309059, 0.07640148, 0.02978136, 0.02279422, 0.04823711, 
    0.06905402, 0.2440904, 0.2926803, 0.2057662, 0.1755347, 0.2836533, 
    0.2840324, 0.2954451, 0.340913, 0.3092428, 0.182207, 0.2287468, 0.215189, 
    0.1769473, 0.330172, 0.2586307, 0.1716149,
  0.103006, 0.2456002, 0.4203206, 0.3726941, 0.2955783, 0.1927092, 0.4852412, 
    0.4820959, 0.3204661, 0.2274733, 0.2376498, 0.2773437, 0.2221556, 
    0.3987752, 0.198215, 0.1615473, 0.2219877, 0.3006354, 0.3442107, 
    0.3489072, 0.3262556, 0.3039494, 0.2804157, 0.345589, 0.2252673, 
    0.06281511, 0.1367227, 0.139236, 0.06396725,
  0.3045572, 0.4204365, 0.3634132, 0.2956215, 0.3704189, 0.3126347, 
    0.3285786, 0.2417591, 0.2923986, 0.3514897, 0.3450606, 0.2559502, 
    0.320345, 0.2653073, 0.3500964, 0.268928, 0.2424663, 0.2984764, 0.303901, 
    0.2268157, 0.2662174, 0.291, 0.2739501, 0.242529, 0.3052205, 0.2320168, 
    0.2893939, 0.2308421, 0.2250693,
  0.2842637, 0.2530896, 0.312331, 0.1995664, 0.2251198, 0.1852858, 0.2010872, 
    0.2064948, 0.1854929, 0.2235428, 0.2688202, 0.2415236, 0.2111865, 
    0.1850135, 0.2120999, 0.2159508, 0.2719158, 0.2387671, 0.2305284, 
    0.2076482, 0.1872745, 0.2665446, 0.2160445, 0.1580663, 0.1510628, 
    0.1775808, 0.2173751, 0.2791499, 0.2893023,
  0.1324903, 0.1584581, 0.1312073, 0.1595871, 0.1365551, 0.1292682, 
    0.1381978, 0.1238476, 0.160451, 0.1331449, 0.2171079, 0.1495404, 
    0.1350804, 0.1548613, 0.1846909, 0.1155725, 0.152444, 0.1124246, 
    0.1060744, 0.09215, 0.1859796, 0.1345875, 0.1877066, 0.2715192, 
    0.09400555, 0.1401314, 0.1730192, 0.1179417, 0.1606383,
  0.02494902, 0.01385349, 0.07176692, 0.0472888, 0.04018718, 0.06382233, 
    0.04655043, 0.04214806, 0.06464277, 0.0690854, 0.05562884, 0.0601982, 
    0.06507308, 0.0726236, 0.09386197, 0.1723729, 0.0653716, 0.09011945, 
    0.1974193, 0.2037665, 0.1430446, 0.04284098, 0.06429061, 0.002617572, 
    0.08736494, 0.1323718, 0.09667499, 0.05326127, 0.04983244,
  6.417181e-08, 7.557124e-06, 0.0261463, 0.03644976, 0.07787628, 0.0182745, 
    0.003938888, 0.1192967, 0.03031322, 0.03284702, 0.01228597, 0.01076858, 
    0.004571231, 0.03038565, 0.07601558, 0.01427649, 0.05250784, 0.06556049, 
    0.1143267, 0.1298553, 0.001281863, 0.0003087325, 0.0007262624, 
    0.000353598, 0.08062348, 0.00364542, 0.06775522, 0.04295635, 0.01620192,
  6.114279e-07, 2.748171e-05, 0.0003215105, 0.1045661, 0.0810921, 0.06782598, 
    0.02663752, 0.04819148, 0.08154126, 0.02028284, 0.07830915, 0.06394968, 
    0.1116667, 0.09357829, 0.05783358, 0.1206669, 0.1449316, 0.04296118, 
    0.02853981, 0.004152756, 8.490464e-05, 1.102753e-07, 1.609344e-06, 
    0.01337931, 0.002582419, 0.0893976, 0.02192758, 0.0009092465, 2.542613e-05,
  0.003727925, 0.06830995, 0.08134381, 0.01965854, 0.005262647, 0.01128582, 
    0.01547883, 0.006238736, 0.03143428, 0.06552009, 0.04508018, 0.02728844, 
    0.1074274, 0.08531339, 0.02885706, 0.01576759, 0.0148683, 0.01366418, 
    0.01021826, 0.002258913, 2.874937e-05, 0.0002624823, 0.02897182, 
    0.3092821, 0.2003774, 0.05013495, 0.08041003, 0.001024839, 0.003758899,
  0.0282441, 0.003983001, 0.004079468, 0.02426569, 0.0005704603, 0.008826579, 
    0.09073711, 0.02415477, 0.006672326, 0.01835369, 0.01292335, 0.02325253, 
    0.1107826, 0.08014753, 0.05246519, 0.04758481, 0.06277102, 0.06274686, 
    0.08042046, 0.07962396, 0.1054744, 0.09206907, 0.1248953, 0.09839818, 
    0.07628654, 0.07536545, 0.04757006, 0.1068422, 0.03512298,
  0.0001186747, 2.273436e-06, 4.312668e-10, 3.463137e-08, 3.566693e-07, 
    -4.509616e-07, 0.122232, 0.1099418, 0.2230704, 0.1530751, 0.06416655, 
    0.01883756, 0.02550531, 0.0206475, 0.03460027, 0.03573063, 0.002322592, 
    6.682841e-05, 3.720177e-07, 0.002996295, 0.0007412087, 0.09131203, 
    0.01508251, 0.01345037, 0.02191208, 0.02250296, 4.092032e-05, 
    2.337068e-06, 0.008397431,
  0.000603632, 9.414912e-06, 1.715928e-06, 6.829987e-07, -1.31366e-05, 
    7.265476e-08, 0.00773913, 0.1869484, 0.2669984, 0.07216169, 0.1020449, 
    0.1110905, 0.09555087, 0.07516657, 0.1088153, 0.02033138, 0.01993416, 
    0.01907391, 3.516718e-07, 1.988348e-07, -1.252672e-05, 0.01546745, 
    0.03862083, 0.04095686, 0.08534379, 0.01707972, 0.003437486, 
    8.668144e-05, 0.001128317,
  0.06622873, 0.06528173, 0.05469413, 0.0972633, -0.0002336634, 3.312544e-06, 
    0.04777945, 0.03237662, 0.01041595, 0.0641636, 0.09332102, 0.06853935, 
    0.1421608, 0.12445, 0.0957467, 0.1770572, 0.1321713, 0.08253238, 
    0.01218143, 0.04460334, 0.01195847, 0.05611617, 0.06885605, 0.05946705, 
    0.09603409, 0.1160765, 0.06562644, 0.032789, 0.05349691,
  0.06265762, 0.1502796, 0.2178356, 0.07791495, 0.04797487, 0.03225104, 
    0.04249652, 0.1144286, 0.1778826, 0.2028543, 0.1897743, 0.2139477, 
    0.1266119, 0.1877405, 0.2322925, 0.2206415, 0.2888531, 0.2536328, 
    0.222003, 0.1627446, 0.1786331, 0.1129207, 0.1366495, 0.1302723, 
    0.2192604, 0.2326286, 0.1867369, 0.1603608, 0.169101,
  0.1764166, 0.1097483, 0.1140219, 0.1961746, 0.2115085, 0.1774021, 
    0.1552108, 0.1514849, 0.272275, 0.2309062, 0.2610056, 0.3572615, 
    0.2449515, 0.2178317, 0.2161077, 0.2291409, 0.3239279, 0.5225832, 
    0.1913074, 0.1268965, 0.1374258, 0.1114165, 0.1640356, 0.2846883, 
    0.1821351, 0.2734559, 0.2595143, 0.3562345, 0.2487585,
  0.2801251, 0.2371659, 0.3024187, 0.1012259, 0.2066973, 0.2397479, 
    0.2501355, 0.1695158, 0.1588733, 0.1727401, 0.1240906, 0.2261037, 
    0.09836055, 0.1477283, 0.1285229, 0.2556827, 0.1518826, 0.1376699, 
    0.1855081, 0.2071872, 0.2084673, 0.1748001, 0.161705, 0.1937655, 
    0.04842274, 0.1571191, 0.2607968, 0.2022439, 0.34883,
  0.2669924, 0.2618147, 0.1441814, 0.2649422, 0.3064666, 0.2741555, 
    0.2050572, 0.2090896, 0.17363, 0.1619189, 0.1635766, 0.1393124, 0.239813, 
    0.2735195, 0.2779117, 0.2613906, 0.2264236, 0.2471113, 0.2964079, 
    0.3744055, 0.3093832, 0.2891317, 0.2117085, 0.1833661, 0.06966868, 
    0.1540207, 0.1697373, 0.1647951, 0.3274015,
  0.1152714, 0.1120449, 0.1088184, 0.1055919, 0.1023654, 0.09913897, 
    0.09591249, 0.08669867, 0.08714453, 0.0875904, 0.08803626, 0.08848213, 
    0.08892798, 0.08937385, 0.0851181, 0.08981436, 0.09451061, 0.09920687, 
    0.1039031, 0.1085994, 0.1132957, 0.1290386, 0.127123, 0.1252073, 
    0.1232917, 0.121376, 0.1194604, 0.1175448, 0.1178526,
  0.1259371, 0.1177407, 0.01877048, 0.00345206, 0.01686813, 0.04018854, 
    0.08394457, 0.08337203, 0.06590895, 0.02408003, 0.04274565, 0.07494841, 
    0.1344742, 0.2340181, 0.2801989, 0.1834259, 0.1911383, 0.259862, 
    0.2791485, 0.2937824, 0.3570481, 0.3266982, 0.1770863, 0.2188845, 
    0.1913712, 0.1597172, 0.3255135, 0.2485339, 0.2149828,
  0.1204227, 0.2714889, 0.4207385, 0.3386552, 0.3056831, 0.1910563, 
    0.5162026, 0.4843023, 0.3012491, 0.228296, 0.2446244, 0.3022086, 
    0.2201591, 0.3781432, 0.1767078, 0.1116167, 0.2053553, 0.276573, 
    0.3205891, 0.3225462, 0.3382947, 0.2678002, 0.2631271, 0.2995478, 
    0.2070452, 0.07933189, 0.1418302, 0.1726669, 0.07055453,
  0.2717943, 0.4344704, 0.33118, 0.2924555, 0.3833877, 0.2633184, 0.3103906, 
    0.2655295, 0.2954969, 0.3558237, 0.3323144, 0.2896508, 0.3224524, 
    0.2218028, 0.2947392, 0.2288893, 0.2708987, 0.2868392, 0.3395089, 
    0.2383128, 0.282153, 0.3031025, 0.280664, 0.288381, 0.2928848, 0.218379, 
    0.2760534, 0.2466706, 0.2451336,
  0.3022171, 0.2460127, 0.3102184, 0.2317355, 0.2478203, 0.2069921, 
    0.2143695, 0.2327339, 0.2327703, 0.2657738, 0.2654282, 0.2573352, 
    0.255466, 0.2264557, 0.232634, 0.2169925, 0.2852853, 0.2651818, 
    0.2758614, 0.243678, 0.2319566, 0.2832067, 0.233212, 0.1740522, 
    0.1635734, 0.2072777, 0.2332769, 0.2886704, 0.3210754,
  0.1473623, 0.1748307, 0.1539914, 0.1896233, 0.1529706, 0.1554582, 
    0.1692019, 0.1528924, 0.1914796, 0.1720885, 0.2262983, 0.18653, 
    0.1451797, 0.1548643, 0.2073957, 0.1221074, 0.1354796, 0.1264622, 
    0.12904, 0.1324181, 0.1938656, 0.1398076, 0.212193, 0.2924386, 0.1151571, 
    0.1617146, 0.1840113, 0.1508255, 0.1857912,
  0.04058171, 0.0279935, 0.06160565, 0.05905757, 0.04993994, 0.07347344, 
    0.07234428, 0.07676886, 0.08689735, 0.09703591, 0.0375086, 0.03329803, 
    0.060529, 0.07432789, 0.09053347, 0.1451372, 0.07319564, 0.1105247, 
    0.1906008, 0.1907149, 0.1616336, 0.05841946, 0.06401724, 0.002779895, 
    0.1155392, 0.1140623, 0.1077278, 0.06513309, 0.05071407,
  -3.212863e-06, -1.412918e-06, 0.09860037, 0.05802104, 0.07823163, 
    0.02773899, 0.03696012, 0.0976128, 0.04430107, 0.04135774, 0.007056464, 
    0.02325504, 0.006130975, 0.01745129, 0.07603683, 0.01963396, 0.07098986, 
    0.08716442, 0.1095118, 0.1239646, 0.02359895, 0.006847861, 0.002489708, 
    0.001749028, 0.1040801, 0.01785487, 0.04932561, 0.06598439, 0.01543923,
  -1.716636e-06, 0.0003942976, 0.00132166, 0.1279134, 0.08271576, 0.06009635, 
    0.02891263, 0.06009474, 0.08568478, 0.02246047, 0.09967975, 0.08818468, 
    0.1249525, 0.08899929, 0.04973964, 0.09783618, 0.1354662, 0.0393704, 
    0.03637414, 0.02111219, 0.0002435993, -1.09581e-06, 4.356143e-07, 
    0.01310465, 0.006569131, 0.01073365, 0.02749958, 0.003852041, 0.002450331,
  0.003044965, 0.07120471, 0.1136941, 0.02480043, 0.01274982, 0.01335756, 
    0.0136359, 0.007257813, 0.03970167, 0.07709449, 0.04027995, 0.02227753, 
    0.09507655, 0.06834217, 0.02424153, 0.01705914, 0.01790934, 0.01811975, 
    0.01520757, 0.003123285, 0.0001374917, 0.0004692307, 0.02330351, 
    0.3117648, 0.206815, 0.04136508, 0.06834381, 0.00384866, 0.002123767,
  0.02694746, 0.002626004, 0.002297312, 0.005440676, 0.0001075742, 
    0.008561796, 0.0790104, 0.02488832, 0.00877736, 0.01651892, 0.0121656, 
    0.02255229, 0.1045443, 0.07326559, 0.05510718, 0.05261571, 0.06979388, 
    0.06799953, 0.08107706, 0.0864292, 0.1099663, 0.08584581, 0.1338282, 
    0.1032098, 0.0728559, 0.08164834, 0.05719271, 0.1049957, 0.03263396,
  2.127757e-05, 7.872832e-07, 2.551106e-09, 3.785409e-08, 1.193626e-07, 
    -2.624219e-06, 0.1024794, 0.1027493, 0.2327644, 0.1425414, 0.06493, 
    0.01934451, 0.03023699, 0.02756225, 0.03102201, 0.04288216, 0.02018083, 
    0.002668998, 1.729538e-06, 0.00595597, 0.0001868064, 0.08716181, 
    0.01300871, 0.01183317, 0.03018146, 0.02786408, 0.002657068, 
    7.640458e-07, 0.004585802,
  0.000558704, 4.40596e-06, 7.675431e-07, 4.296051e-07, -3.943188e-06, 
    7.650784e-08, 0.004122983, 0.1506315, 0.2702563, 0.06583814, 0.1084997, 
    0.1248495, 0.0800475, 0.07092213, 0.09934168, 0.02939516, 0.03243237, 
    0.01991428, 0.0003046344, 1.583028e-07, 3.758957e-06, 0.02335139, 
    0.03817901, 0.05035613, 0.08451601, 0.02444721, 0.03709564, 0.0008706558, 
    0.002626187,
  0.05595091, 0.05563781, 0.05368201, 0.09840091, -0.0001349709, 7.03599e-07, 
    0.03409012, 0.01308058, 0.004800297, 0.04244995, 0.09233655, 0.06443566, 
    0.1470719, 0.1196232, 0.09016972, 0.2037969, 0.1210449, 0.09043136, 
    0.009987179, 0.05050194, 0.003475757, 0.05122252, 0.06892563, 0.04620461, 
    0.09510418, 0.1398126, 0.09254833, 0.04471561, 0.04256245,
  0.04601803, 0.1926322, 0.2113846, 0.08329622, 0.04370679, 0.03083229, 
    0.01940499, 0.114019, 0.186052, 0.1896687, 0.1750139, 0.2177605, 
    0.1171982, 0.1818611, 0.2265567, 0.2511466, 0.2669979, 0.2520233, 
    0.1928335, 0.1361765, 0.1999031, 0.1117285, 0.1310681, 0.14673, 
    0.2036631, 0.2327309, 0.1933424, 0.1745016, 0.1384328,
  0.1915839, 0.1243409, 0.12341, 0.1946181, 0.2178161, 0.2145632, 0.1382981, 
    0.1393023, 0.2909395, 0.2522669, 0.2891332, 0.3627516, 0.2480655, 
    0.2496192, 0.2239189, 0.2017619, 0.3480794, 0.5245484, 0.2258183, 
    0.1454063, 0.1273485, 0.09460021, 0.1373575, 0.2847005, 0.1707531, 
    0.243601, 0.2749722, 0.3607174, 0.2382024,
  0.3439461, 0.2101605, 0.3313381, 0.101425, 0.2203103, 0.2427977, 0.2089619, 
    0.1951965, 0.09614165, 0.119112, 0.1492722, 0.1873351, 0.134544, 
    0.1251781, 0.06471317, 0.1495975, 0.1338979, 0.1479794, 0.151533, 
    0.1876806, 0.1656359, 0.173789, 0.1665239, 0.1310092, 0.04078816, 
    0.1890893, 0.2549656, 0.2090589, 0.3110623,
  0.2241543, 0.2247296, 0.1409832, 0.2277882, 0.2098027, 0.2175601, 
    0.1648978, 0.1763285, 0.1309777, 0.1048448, 0.1217352, 0.09393747, 
    0.152426, 0.2487415, 0.2739004, 0.2466964, 0.2236328, 0.2039521, 
    0.2251793, 0.2756717, 0.2217648, 0.2414497, 0.3279068, 0.1789322, 
    0.07695271, 0.1157537, 0.1781394, 0.2044684, 0.3099363,
  0.1255099, 0.1244332, 0.1233566, 0.12228, 0.1212033, 0.1201267, 0.1190501, 
    0.1273159, 0.1293328, 0.1313497, 0.1333666, 0.1353836, 0.1374005, 
    0.1394174, 0.1338656, 0.1352563, 0.1366471, 0.1380378, 0.1394286, 
    0.1408193, 0.1422101, 0.1385111, 0.1361801, 0.133849, 0.131518, 0.129187, 
    0.126856, 0.1245249, 0.1263712,
  0.1567555, 0.1483307, 0.1017282, 0.009757032, 0.02534306, 0.05509933, 
    0.1084683, 0.09772044, 0.05279203, 0.02373246, 0.05230467, 0.09218056, 
    0.183873, 0.1969057, 0.2856402, 0.2020163, 0.1912928, 0.2342243, 
    0.2908754, 0.3015611, 0.3763896, 0.334296, 0.2102918, 0.1963359, 
    0.1863747, 0.1584408, 0.3174681, 0.2369267, 0.2595317,
  0.1397197, 0.2632169, 0.3597602, 0.3276955, 0.3084334, 0.207954, 0.4963048, 
    0.5008801, 0.2922658, 0.2424275, 0.2546914, 0.2889295, 0.2324465, 0.3782, 
    0.2234281, 0.1341934, 0.1623344, 0.2881502, 0.3848834, 0.3143516, 
    0.3330786, 0.2715628, 0.2786666, 0.3310673, 0.1897583, 0.09414502, 
    0.1635469, 0.1798094, 0.08907685,
  0.3411208, 0.4742833, 0.3636842, 0.3175904, 0.3858845, 0.3031228, 
    0.3230857, 0.2921452, 0.3445394, 0.391827, 0.3859219, 0.2885636, 
    0.3390106, 0.2619176, 0.2607708, 0.2359142, 0.2566973, 0.2599353, 
    0.3491775, 0.2594229, 0.3221639, 0.306588, 0.372705, 0.3444753, 0.292923, 
    0.2448439, 0.2932318, 0.2874702, 0.3026459,
  0.3377506, 0.2913305, 0.3302496, 0.2390213, 0.2807324, 0.2217337, 0.24949, 
    0.2680628, 0.2521523, 0.2949414, 0.2846595, 0.2745332, 0.248533, 
    0.2347209, 0.278589, 0.2733817, 0.3066975, 0.2946196, 0.3343144, 
    0.2861085, 0.2795167, 0.3207313, 0.2527448, 0.198139, 0.1708204, 
    0.2480915, 0.2699591, 0.3177162, 0.3517555,
  0.152475, 0.1812292, 0.197275, 0.2072673, 0.2020844, 0.2161719, 0.1765329, 
    0.1836963, 0.2260132, 0.1764104, 0.226101, 0.191172, 0.1510089, 
    0.1763907, 0.2067352, 0.1334091, 0.152413, 0.1366607, 0.1763427, 
    0.1778488, 0.2085182, 0.1707535, 0.2444087, 0.3215324, 0.1304701, 
    0.1723835, 0.2107429, 0.1572763, 0.1993693,
  0.1079719, 0.05581063, 0.04035181, 0.07503322, 0.07613334, 0.1215483, 
    0.07978006, 0.09916096, 0.1340588, 0.1282707, 0.01142167, 0.02636626, 
    0.06646544, 0.07003728, 0.09279069, 0.1549979, 0.09354028, 0.1432976, 
    0.1709978, 0.1579211, 0.1735659, 0.07054023, 0.09782517, 0.004734544, 
    0.1258472, 0.1218076, 0.1036993, 0.05421409, 0.06201907,
  0.002529843, 9.961872e-08, 0.01603224, 0.06282018, 0.08460165, 0.03662888, 
    0.09083959, 0.1020041, 0.08048337, 0.04781827, 0.002073405, 0.02662122, 
    0.02757869, 0.01130767, 0.09073924, 0.02593142, 0.130219, 0.1090783, 
    0.1232288, 0.1098098, 0.09795853, 0.06260587, 0.018396, 0.003756572, 
    0.09856349, 0.09348426, 0.04030576, 0.06051372, 0.04665386,
  9.688399e-08, -1.587703e-05, 0.004894386, 0.1496903, 0.08291062, 
    0.06022957, 0.02658634, 0.06676796, 0.08359512, 0.02595384, 0.08911818, 
    0.098378, 0.1466624, 0.07760758, 0.04143203, 0.077521, 0.1074231, 
    0.03911611, 0.02928435, 0.0330218, 0.003724511, 0.0002792249, 
    6.392244e-07, 0.02019819, 0.00607996, 0.0009203121, 0.02779424, 
    0.01387571, 0.01892816,
  0.005264095, 0.08710522, 0.1060189, 0.01802103, 0.02001375, 0.01712718, 
    0.01317337, 0.009538609, 0.04888281, 0.09839886, 0.02847466, 0.01765541, 
    0.08328153, 0.04915484, 0.02167437, 0.01928879, 0.01962726, 0.01715089, 
    0.01606823, 0.006441544, 0.001185834, 0.002286351, 0.01820908, 0.2990781, 
    0.2060136, 0.03146838, 0.05832759, 0.01121608, 0.000704214,
  0.0260358, 0.001626852, 0.001113996, 0.001214506, 3.384137e-05, 0.01094917, 
    0.07093167, 0.02543452, 0.02090048, 0.0163568, 0.01458876, 0.02125388, 
    0.08776811, 0.06337818, 0.04787273, 0.05052866, 0.07415626, 0.08401573, 
    0.08314429, 0.08748321, 0.1031702, 0.08258761, 0.1244581, 0.1050731, 
    0.06328575, 0.08557821, 0.0786094, 0.1023625, 0.03484948,
  1.472696e-06, 3.71937e-07, 1.737869e-09, 4.253608e-08, 7.261385e-08, 
    -6.263433e-05, 0.086531, 0.09164254, 0.2362866, 0.1387356, 0.05851496, 
    0.02043402, 0.026441, 0.02566108, 0.02641847, 0.03285101, 0.06073698, 
    0.01218796, 2.289957e-05, 0.008074942, 0.0004726514, 0.07831346, 
    0.01272247, 0.01163094, 0.03109693, 0.0422942, 0.02739655, 2.893618e-06, 
    0.002866783,
  0.0004121693, 1.681083e-06, 2.870069e-07, 2.956048e-07, -8.439513e-08, 
    5.344735e-08, 0.002279094, 0.1116282, 0.2705557, 0.06403509, 0.1121162, 
    0.1506504, 0.06604674, 0.05543438, 0.09914924, 0.03885959, 0.0495868, 
    0.05463782, 0.01690006, 1.121075e-07, 3.242405e-06, 0.02445478, 
    0.01857056, 0.05412539, 0.07885865, 0.04082536, 0.09075371, 0.01415971, 
    0.003566457,
  0.03917028, 0.04133445, 0.04620707, 0.09853276, -2.824735e-05, 
    3.919465e-07, 0.02110359, 0.006681844, 0.002706714, 0.0350959, 
    0.09550583, 0.0624418, 0.1515282, 0.1297664, 0.1148523, 0.2070303, 
    0.1427537, 0.1149271, 0.02031941, 0.0491644, 0.00130995, 0.04467133, 
    0.0707928, 0.04846651, 0.1124414, 0.1795362, 0.1689255, 0.09051184, 
    0.03934824,
  0.05113733, 0.1718275, 0.2193041, 0.08123907, 0.02770072, 0.02349392, 
    0.009809452, 0.1306353, 0.180558, 0.1671733, 0.1681685, 0.2029484, 
    0.09163073, 0.1879551, 0.2487341, 0.2548456, 0.2891695, 0.3054208, 
    0.2061941, 0.09718958, 0.191697, 0.1282825, 0.1314656, 0.1398764, 
    0.1838735, 0.2531081, 0.2047523, 0.187085, 0.1518631,
  0.206203, 0.1626698, 0.1046389, 0.1880231, 0.2538511, 0.1942464, 0.161512, 
    0.2052118, 0.2763757, 0.221779, 0.3105121, 0.3308317, 0.2640359, 
    0.2708037, 0.2362173, 0.1721121, 0.3840559, 0.5352602, 0.2938403, 
    0.1074374, 0.09145511, 0.05695391, 0.1087475, 0.2322808, 0.200519, 
    0.2056062, 0.3407049, 0.3760518, 0.2583586,
  0.3496624, 0.246967, 0.3428685, 0.1172255, 0.2807266, 0.2337509, 0.1980715, 
    0.1819732, 0.1107989, 0.1229015, 0.1717004, 0.1605963, 0.1111742, 
    0.1422445, 0.05414914, 0.109121, 0.1714629, 0.1528709, 0.1363026, 
    0.1715052, 0.1463931, 0.1779361, 0.2412309, 0.1703475, 0.05550118, 
    0.215731, 0.2413994, 0.2266721, 0.2909086,
  0.3031205, 0.3069035, 0.2394281, 0.225252, 0.2023565, 0.2717945, 0.151761, 
    0.192991, 0.1474276, 0.1592749, 0.1493863, 0.1108896, 0.1460976, 
    0.2426686, 0.2697819, 0.3266393, 0.3196825, 0.2762031, 0.2767482, 
    0.3022693, 0.2566614, 0.25952, 0.2535236, 0.1827846, 0.05638634, 
    0.09899327, 0.1475582, 0.2547486, 0.3551068,
  0.1449172, 0.1426661, 0.140415, 0.1381639, 0.1359129, 0.1336618, 0.1314107, 
    0.1427133, 0.1453551, 0.1479969, 0.1506387, 0.1532805, 0.1559223, 
    0.1585641, 0.1576878, 0.1597432, 0.1617987, 0.1638542, 0.1659097, 
    0.1679652, 0.1700207, 0.1705502, 0.168104, 0.1656578, 0.1632116, 
    0.1607654, 0.1583192, 0.155873, 0.1467181,
  0.1848758, 0.1825048, 0.1598238, 0.04437266, 0.04196434, 0.08978102, 
    0.1144027, 0.09533601, 0.03233343, 0.01965851, 0.06580717, 0.1000832, 
    0.2096821, 0.1621481, 0.2884534, 0.231016, 0.1902036, 0.2118024, 
    0.2820057, 0.3124871, 0.4501704, 0.3589633, 0.2343068, 0.1628395, 
    0.183062, 0.178402, 0.2887352, 0.2245831, 0.2718294,
  0.1975214, 0.2794765, 0.3611781, 0.3118052, 0.3104805, 0.2505952, 
    0.4985298, 0.5249262, 0.280873, 0.2505943, 0.2614306, 0.2952784, 
    0.2494389, 0.3743683, 0.2382878, 0.1847715, 0.2107179, 0.3801528, 
    0.3624139, 0.3711405, 0.3502472, 0.3000081, 0.279002, 0.3310927, 
    0.1849505, 0.11004, 0.1790834, 0.1930711, 0.1110949,
  0.3619712, 0.5059398, 0.3807599, 0.3766284, 0.4447218, 0.3800135, 
    0.3774232, 0.3389661, 0.3983024, 0.4490759, 0.3705238, 0.3009818, 
    0.3680727, 0.3996706, 0.3147283, 0.2719837, 0.249588, 0.2666989, 
    0.3664888, 0.2860633, 0.2998845, 0.3737238, 0.4245816, 0.4009234, 
    0.3928672, 0.2494474, 0.2866764, 0.2996829, 0.3035809,
  0.345416, 0.3121763, 0.3489757, 0.2532392, 0.2718968, 0.2576965, 0.2978421, 
    0.335854, 0.2695436, 0.2411139, 0.3101113, 0.303643, 0.2427668, 0.26863, 
    0.2966035, 0.3501925, 0.3653076, 0.3417413, 0.3818951, 0.3465745, 
    0.3355314, 0.3273649, 0.2708091, 0.2238587, 0.1955267, 0.2596386, 
    0.3413161, 0.3394787, 0.3154941,
  0.1583836, 0.184471, 0.2072637, 0.2049237, 0.2232032, 0.2095582, 0.1961329, 
    0.2171736, 0.2415881, 0.1561951, 0.1996484, 0.17449, 0.1383517, 
    0.1577465, 0.2317419, 0.160431, 0.1685932, 0.1319075, 0.1955498, 
    0.2483032, 0.272447, 0.2513905, 0.2589706, 0.3678864, 0.1452381, 
    0.1558932, 0.1932857, 0.1833466, 0.2139196,
  0.1629295, 0.07161062, 0.02539625, 0.1408075, 0.09840856, 0.158676, 
    0.1277985, 0.1309442, 0.1749146, 0.1726083, 0.008490744, 0.01250984, 
    0.04470414, 0.0821718, 0.1472009, 0.2065703, 0.1535295, 0.165747, 
    0.1974348, 0.187572, 0.1904548, 0.08261202, 0.1183652, 0.009595805, 
    0.09502039, 0.1737182, 0.1248996, 0.08245853, 0.1435874,
  0.07757968, -1.090061e-06, 0.003308511, 0.08397515, 0.1121762, 0.03736014, 
    0.1372238, 0.1975449, 0.0911176, 0.03084267, 0.0003860793, 0.01352298, 
    0.1140264, 0.037747, 0.09323566, 0.03264049, 0.1151158, 0.1184001, 
    0.1225332, 0.1181634, 0.1673611, 0.1218842, 0.05100335, 0.0004990136, 
    0.09902291, 0.05457887, 0.04671957, 0.1115472, 0.1627246,
  0.0001340013, 1.844054e-07, 0.01339854, 0.1643445, 0.07460988, 0.05578753, 
    0.04040051, 0.0805722, 0.07603772, 0.03423981, 0.09804066, 0.1047667, 
    0.1553158, 0.06486739, 0.03883014, 0.07000933, 0.07786973, 0.0371431, 
    0.03030602, 0.03817032, 0.02130392, 0.01953135, 5.760081e-06, 0.03811922, 
    0.01505125, 0.0001667914, 0.04200209, 0.03891993, 0.03881991,
  0.01033185, 0.1025285, 0.1046726, 0.01276508, 0.02843397, 0.02398052, 
    0.01678858, 0.01540775, 0.06210354, 0.1173033, 0.02250735, 0.01460553, 
    0.06947874, 0.03558036, 0.02444565, 0.02383347, 0.0187007, 0.01755996, 
    0.0156226, 0.0171442, 0.01743761, 0.007852179, 0.007724113, 0.2822368, 
    0.1889251, 0.02893328, 0.05259357, 0.01496619, 0.003014786,
  0.02562094, 0.003339536, 0.0005622882, -3.842236e-05, -2.809101e-06, 
    0.01504725, 0.06412813, 0.02920308, 0.01930617, 0.02086018, 0.02390794, 
    0.0221546, 0.07499149, 0.05513926, 0.04457886, 0.0443597, 0.07700181, 
    0.09138501, 0.08840432, 0.08906391, 0.08945432, 0.06915805, 0.1226572, 
    0.1104653, 0.05226807, 0.08486335, 0.08989655, 0.08702752, 0.03290274,
  1.017123e-06, 2.105983e-07, 5.816529e-10, 3.936576e-08, 6.060088e-08, 
    -0.000235601, 0.06701531, 0.08115721, 0.2277396, 0.1300224, 0.05610738, 
    0.02444262, 0.02741383, 0.0274374, 0.02831816, 0.03552784, 0.082779, 
    0.04548194, 0.004316982, 0.01293391, 0.003995431, 0.07261682, 0.01549856, 
    0.01245191, 0.03600492, 0.06723548, 0.06604791, 0.0003612424, 0.001785558,
  0.0002359792, 9.229059e-07, 6.883845e-08, 2.149825e-07, 6.29049e-11, 
    4.043271e-08, 0.001569345, 0.1025024, 0.2699035, 0.06028725, 0.1149404, 
    0.1612593, 0.05767955, 0.04828649, 0.09073398, 0.03741244, 0.0931555, 
    0.1003039, 0.0701412, -3.862023e-07, 2.523898e-06, 0.02461987, 
    0.01317279, 0.05343474, 0.06912593, 0.04515139, 0.106806, 0.05773059, 
    0.006661933,
  0.03196473, 0.02755035, 0.02157499, 0.1003222, -2.75891e-06, 2.900362e-07, 
    0.0179464, 0.004307374, 0.001691968, 0.03081159, 0.1040215, 0.06995282, 
    0.1614286, 0.1467068, 0.1761283, 0.2315273, 0.171236, 0.1634528, 
    0.04937646, 0.03460336, 0.0006729022, 0.03789477, 0.06571053, 0.0404803, 
    0.1396941, 0.1990683, 0.1716986, 0.1139543, 0.04788649,
  0.03607879, 0.1530609, 0.1892979, 0.07519262, 0.02106058, 0.008844109, 
    0.01000274, 0.134558, 0.158373, 0.1391708, 0.1505955, 0.1883128, 
    0.1039362, 0.202483, 0.2712274, 0.2811971, 0.373526, 0.3471957, 
    0.2432178, 0.07942493, 0.1646615, 0.08991101, 0.1266727, 0.1425481, 
    0.1654914, 0.2518989, 0.2333523, 0.2193243, 0.1883955,
  0.2262671, 0.1537787, 0.06705739, 0.2161007, 0.2379201, 0.1624785, 
    0.08706514, 0.2310302, 0.2509878, 0.2065703, 0.2774304, 0.3477985, 
    0.2738514, 0.2919428, 0.2660004, 0.214086, 0.3414115, 0.5413304, 
    0.2753475, 0.06998003, 0.06632622, 0.04084975, 0.08834735, 0.2022258, 
    0.1706475, 0.148688, 0.427512, 0.413198, 0.2853499,
  0.3441744, 0.2651647, 0.333338, 0.1384159, 0.2920369, 0.2416821, 0.2353802, 
    0.1860077, 0.09831061, 0.08997382, 0.1505166, 0.1936067, 0.09103267, 
    0.1529571, 0.09646612, 0.1552899, 0.2366297, 0.1298668, 0.1200638, 
    0.1394098, 0.1758338, 0.1940123, 0.2689704, 0.2175336, 0.05020131, 
    0.2114366, 0.2396771, 0.2513537, 0.3182606,
  0.401549, 0.3484557, 0.2773125, 0.2723879, 0.2726563, 0.2959498, 0.228822, 
    0.2194142, 0.2072726, 0.1946594, 0.1561376, 0.1866952, 0.2269922, 
    0.3045364, 0.3129981, 0.4113488, 0.3628235, 0.4193598, 0.4077237, 
    0.4260794, 0.2996578, 0.2474915, 0.2129316, 0.1677178, 0.0941296, 
    0.08805554, 0.112751, 0.2756173, 0.3999294,
  0.1756151, 0.1719283, 0.1682415, 0.1645547, 0.1608679, 0.1571811, 
    0.1534942, 0.1601699, 0.163068, 0.1659662, 0.1688643, 0.1717624, 
    0.1746605, 0.1775587, 0.1727451, 0.1760493, 0.1793535, 0.1826576, 
    0.1859618, 0.189266, 0.1925702, 0.2061897, 0.2036742, 0.2011587, 
    0.1986433, 0.1961278, 0.1936123, 0.1910968, 0.1785646,
  0.2189726, 0.1882457, 0.1713711, 0.08708274, 0.06280944, 0.104603, 0.1043, 
    0.08610003, 0.02353792, 0.0232601, 0.05594788, 0.09441943, 0.2328893, 
    0.0897872, 0.2753419, 0.2327612, 0.2100749, 0.2049722, 0.3051896, 
    0.3094372, 0.488861, 0.3928792, 0.2250333, 0.1220104, 0.1733824, 
    0.1960952, 0.2539153, 0.2173022, 0.2805482,
  0.2159271, 0.2759194, 0.3716611, 0.2881779, 0.3230519, 0.2896067, 
    0.4251908, 0.5245163, 0.2709755, 0.2589831, 0.2513845, 0.2698545, 
    0.2607336, 0.3449206, 0.2555771, 0.3188717, 0.3403184, 0.3958388, 
    0.3889298, 0.3554115, 0.3395852, 0.3693923, 0.2765935, 0.3419545, 
    0.2038653, 0.1435823, 0.2014814, 0.2089726, 0.1194567,
  0.3699675, 0.5321945, 0.3462879, 0.3765652, 0.4261746, 0.4556423, 
    0.4563886, 0.458296, 0.3788106, 0.4740305, 0.4027639, 0.3757505, 
    0.4151934, 0.4100423, 0.4184284, 0.3343986, 0.2993884, 0.3053927, 
    0.3525429, 0.3061899, 0.3471885, 0.3928745, 0.3351124, 0.4109185, 
    0.436313, 0.2857062, 0.2895839, 0.3786707, 0.303275,
  0.3671076, 0.3426391, 0.3472227, 0.280555, 0.2993383, 0.2857423, 0.3515889, 
    0.3415566, 0.2447403, 0.2512455, 0.3337865, 0.3115118, 0.2268226, 
    0.3165846, 0.3428789, 0.3788971, 0.4202625, 0.3338536, 0.3420225, 
    0.4022059, 0.3581786, 0.3254597, 0.246406, 0.2507174, 0.1962754, 
    0.2427509, 0.3666041, 0.3359959, 0.3429926,
  0.186585, 0.1991068, 0.1668853, 0.1791151, 0.1888609, 0.1721398, 0.2253021, 
    0.2728083, 0.2370891, 0.1368622, 0.1797155, 0.1405987, 0.1128269, 
    0.1444538, 0.2777761, 0.2306272, 0.200974, 0.1459286, 0.1859275, 
    0.2116723, 0.3013782, 0.284541, 0.2216945, 0.4375213, 0.08662543, 
    0.1163358, 0.1669867, 0.1767541, 0.2348825,
  0.2102489, 0.03543054, 0.02159934, 0.09813385, 0.1235444, 0.1684553, 
    0.2143372, 0.1724787, 0.1514907, 0.08209038, 0.00920599, 0.006872537, 
    0.03857509, 0.06732244, 0.1234869, 0.2010261, 0.1334178, 0.1030563, 
    0.1433, 0.153506, 0.1986206, 0.1579919, 0.1384794, 0.007529018, 
    0.1108723, 0.1304239, 0.09597989, 0.1399368, 0.1479813,
  0.2243398, -5.153781e-05, 0.0009359595, 0.03975658, 0.1233893, 0.06474042, 
    0.1317085, 0.2170746, 0.1133958, 0.04434313, 0.0001775212, 0.01265539, 
    0.1542839, 0.1229734, 0.1096776, 0.09305482, 0.09298258, 0.1138423, 
    0.09588407, 0.15985, 0.1688312, 0.1842154, 0.2274923, 1.292279e-05, 
    0.1035329, 0.01300313, 0.05590184, 0.1761115, 0.176368,
  0.03941384, 6.120987e-08, 0.006183764, 0.1399072, 0.07652149, 0.06309909, 
    0.06150818, 0.08999582, 0.09023888, 0.04951435, 0.09708579, 0.1001203, 
    0.1540336, 0.05896585, 0.04259031, 0.0606507, 0.07599201, 0.05975186, 
    0.06049786, 0.05523674, 0.08470138, 0.1905673, -0.000118299, 0.0889563, 
    0.002976077, 8.374456e-06, 0.07469848, 0.0422448, 0.1685514,
  0.03124031, 0.1087783, 0.09677924, 0.01288699, 0.04148911, 0.0474317, 
    0.02697239, 0.02714153, 0.06703255, 0.1028423, 0.02698423, 0.01927073, 
    0.06458806, 0.03207643, 0.03132819, 0.0444925, 0.02328451, 0.02295769, 
    0.01738861, 0.02164499, 0.03039776, 0.02996051, 0.005499589, 0.2483705, 
    0.1630833, 0.02982797, 0.05125827, 0.0195549, 0.01878082,
  0.02133348, 0.00464482, 0.0002705898, -0.0003166624, 6.986946e-07, 
    0.01885008, 0.05948422, 0.03923814, 0.008117518, 0.03169199, 0.02925083, 
    0.02867556, 0.07090727, 0.04848084, 0.04430719, 0.04674544, 0.07690124, 
    0.1097364, 0.108789, 0.1060408, 0.08475901, 0.06352641, 0.1352611, 
    0.1079939, 0.05312175, 0.08473517, 0.1022899, 0.08443989, 0.02483867,
  7.456555e-07, 1.408244e-07, 5.083788e-10, 3.880219e-08, 5.40476e-08, 
    0.002912145, 0.04742147, 0.05823299, 0.2132703, 0.1260405, 0.05419721, 
    0.03458392, 0.03445705, 0.03477738, 0.03664796, 0.05154232, 0.08676497, 
    0.1434179, 0.04101631, 0.01885908, 0.006424457, 0.06946315, 0.01997034, 
    0.01348431, 0.04535193, 0.07731688, 0.1497202, 0.01656005, 0.001003945,
  8.452262e-05, 5.967438e-07, -1.345073e-06, 1.799381e-07, 8.158625e-09, 
    3.281803e-08, 0.0005912908, 0.08640065, 0.2744769, 0.06417156, 0.127785, 
    0.1949797, 0.07160208, 0.0556353, 0.09210258, 0.0453248, 0.08901519, 
    0.1354653, 0.205026, 0.0003097021, 1.849594e-06, 0.02356189, 0.007249536, 
    0.05678333, 0.07616002, 0.04542607, 0.1376164, 0.1720557, 0.004251348,
  0.02860543, 0.01997136, 0.01159585, 0.1002303, 2.754573e-05, 2.197501e-07, 
    0.01531535, 0.0002344725, 0.0004730736, 0.02956143, 0.1110025, 
    0.07791572, 0.1693441, 0.1994586, 0.2007262, 0.2637753, 0.264699, 
    0.255519, 0.1464599, 0.04908773, 0.0001472243, 0.03744979, 0.0562852, 
    0.02728691, 0.1775189, 0.2429622, 0.2177591, 0.1794434, 0.06229281,
  0.03176851, 0.1212458, 0.1400528, 0.05921057, 0.01851002, 0.002659569, 
    0.01384407, 0.1339862, 0.1325471, 0.1075062, 0.1246909, 0.168856, 
    0.1386894, 0.2222729, 0.3191845, 0.3820402, 0.4541058, 0.400759, 
    0.3329754, 0.07959082, 0.1356981, 0.08397071, 0.1233362, 0.1428699, 
    0.1512291, 0.2700667, 0.2312725, 0.2738193, 0.2291782,
  0.2214004, 0.1069351, 0.03166665, 0.144125, 0.218964, 0.112513, 0.06418445, 
    0.1332147, 0.2081769, 0.1852568, 0.2831917, 0.3321058, 0.2525071, 
    0.3014975, 0.290356, 0.2488916, 0.3074343, 0.5262195, 0.2649568, 
    0.05486584, 0.04738504, 0.02549997, 0.07953071, 0.1759875, 0.1679424, 
    0.1410245, 0.4725406, 0.4222963, 0.3425722,
  0.3878547, 0.3682677, 0.3530388, 0.1610884, 0.3698496, 0.2356422, 
    0.2307803, 0.1480049, 0.0877631, 0.09963074, 0.1332711, 0.1959465, 
    0.1224555, 0.1734505, 0.07574747, 0.1745016, 0.2766955, 0.1300613, 
    0.0896427, 0.1240955, 0.2377153, 0.2621526, 0.2447632, 0.2119968, 
    0.05557366, 0.204305, 0.2422617, 0.2840512, 0.4307166,
  0.4019652, 0.3802158, 0.2607674, 0.3164225, 0.3389436, 0.273385, 0.2873341, 
    0.2532161, 0.2246305, 0.2190305, 0.1998813, 0.1872357, 0.2022444, 
    0.3420952, 0.4431491, 0.4862061, 0.4792792, 0.4470503, 0.4140448, 
    0.4907647, 0.3317185, 0.2711296, 0.2221656, 0.2319907, 0.06701408, 
    0.1073273, 0.1410366, 0.3274834, 0.4387226,
  0.2020522, 0.1982561, 0.19446, 0.1906639, 0.1868678, 0.1830717, 0.1792756, 
    0.1806882, 0.1831958, 0.1857033, 0.1882109, 0.1907185, 0.1932261, 
    0.1957337, 0.1814903, 0.1865346, 0.1915788, 0.1966231, 0.2016673, 
    0.2067116, 0.2117558, 0.2381026, 0.2343468, 0.2305911, 0.2268354, 
    0.2230797, 0.2193239, 0.2155682, 0.2050891,
  0.227085, 0.1913392, 0.1941336, 0.1345104, 0.07096787, 0.1330339, 
    0.1317222, 0.09130883, 0.02774674, 0.04081819, 0.05969962, 0.1149607, 
    0.259928, 0.03448752, 0.2571658, 0.2313316, 0.1836293, 0.2203936, 
    0.3234594, 0.3447712, 0.5371015, 0.4328003, 0.1991605, 0.1241918, 
    0.1692192, 0.2130072, 0.2474903, 0.2127722, 0.2920038,
  0.1515571, 0.2354362, 0.3601238, 0.260403, 0.3294241, 0.3220529, 0.3514622, 
    0.5271396, 0.2593899, 0.2822808, 0.2548482, 0.2566257, 0.2803304, 
    0.3311293, 0.3261189, 0.3734178, 0.4631709, 0.4553185, 0.4211126, 
    0.3619551, 0.3770745, 0.3714325, 0.2969305, 0.3410782, 0.206025, 
    0.1762505, 0.246857, 0.2461224, 0.1121138,
  0.4005442, 0.5316422, 0.3422159, 0.345221, 0.3852078, 0.4372958, 0.4987972, 
    0.4011311, 0.3297991, 0.4182776, 0.3801422, 0.3536951, 0.4439973, 
    0.3860174, 0.4499421, 0.4008468, 0.3972628, 0.359741, 0.3739631, 
    0.3306919, 0.3619137, 0.3369952, 0.2897578, 0.3688386, 0.4337083, 
    0.31893, 0.3210676, 0.3650797, 0.3047872,
  0.3651959, 0.3483695, 0.3573647, 0.3320703, 0.3315893, 0.2970812, 
    0.3924341, 0.2994764, 0.2688463, 0.2415436, 0.257945, 0.2777838, 
    0.1940323, 0.3462791, 0.3240567, 0.3981295, 0.4048668, 0.3410608, 
    0.2987477, 0.3976317, 0.308397, 0.3583973, 0.2491811, 0.27486, 0.1503292, 
    0.2646718, 0.3272187, 0.2811702, 0.3366669,
  0.1773773, 0.1602811, 0.1312157, 0.1452947, 0.2127035, 0.1157203, 
    0.2129091, 0.2279855, 0.1647956, 0.07465441, 0.1420735, 0.1291771, 
    0.0710827, 0.1043482, 0.3454089, 0.1678122, 0.1513418, 0.1639816, 
    0.1804843, 0.133289, 0.2616181, 0.2315575, 0.1851231, 0.4680575, 
    0.04846838, 0.0761436, 0.1349892, 0.1678942, 0.2148954,
  0.2305536, 0.03748579, 0.02954516, 0.03698406, 0.117109, 0.1569931, 
    0.1622464, 0.154043, 0.08727881, 0.03726133, 0.004243174, 0.002886424, 
    0.0326841, 0.0317861, 0.07766517, 0.1455368, 0.06616574, 0.04723494, 
    0.09850611, 0.1500842, 0.18121, 0.1485524, 0.1344184, 0.008663789, 
    0.1060433, 0.09932302, 0.08971894, 0.08344731, 0.08675233,
  0.19995, -9.333923e-05, 7.847502e-05, 0.01253695, 0.06172722, 0.04610134, 
    0.07143693, 0.1503974, 0.1596476, 0.03543207, 0.0001463325, 0.008992259, 
    0.03466152, 0.09422714, 0.1103338, 0.07938835, 0.09115406, 0.09721717, 
    0.09913293, 0.1260887, 0.08565642, 0.211002, 0.2914059, 0.001260386, 
    0.1332684, 0.01703971, 0.03219921, 0.0684203, 0.1082234,
  0.1129725, 7.786614e-08, 0.005917856, 0.1195242, 0.06634957, 0.06516668, 
    0.05017856, 0.09764545, 0.08809994, 0.08337938, 0.1076813, 0.07583298, 
    0.1552139, 0.07062413, 0.05285732, 0.06413092, 0.06660321, 0.05809727, 
    0.07699455, 0.0446005, 0.1077875, 0.2943473, 0.15434, 0.06306051, 
    0.000713025, 6.323796e-06, 0.04913456, 0.08322868, 0.3154662,
  0.1051869, 0.03243213, 0.05465742, 0.01817175, 0.04916075, 0.1223305, 
    0.1145279, 0.08587196, 0.04450103, 0.05959501, 0.0706103, 0.08190936, 
    0.09596515, 0.0913351, 0.06511615, 0.1187719, 0.07161339, 0.07553392, 
    0.0600806, 0.06069083, 0.05493847, 0.0924156, 0.02480996, 0.2008159, 
    0.1096375, 0.03399206, 0.0586984, 0.05338803, 0.06067371,
  0.01467476, 0.003743429, 0.0001473763, -0.0002262811, -1.68784e-07, 
    0.01943778, 0.05641573, 0.0443935, 0.002876666, 0.1057331, 0.0321887, 
    0.04318498, 0.07227109, 0.05828315, 0.04735514, 0.04849901, 0.07370857, 
    0.1614623, 0.1902283, 0.1407487, 0.0992404, 0.089063, 0.1538104, 
    0.123334, 0.05367739, 0.08733002, 0.1289369, 0.1045439, 0.01009639,
  5.787538e-07, 1.258586e-07, 5.001822e-10, 4.026905e-08, 5.049885e-08, 
    0.02141199, 0.03828837, 0.04731568, 0.2042615, 0.123529, 0.05566471, 
    0.05917268, 0.04858326, 0.04595566, 0.04087719, 0.05249868, 0.04804705, 
    0.1781773, 0.2619534, 0.04002685, 0.01151991, 0.07272635, 0.03168265, 
    0.01120822, 0.04686795, 0.05735919, 0.2154844, 0.02822254, 0.0004051714,
  5.13793e-05, -4.178783e-07, -0.0001088184, 1.610493e-07, 1.449297e-08, 
    2.807053e-08, 0.0004293901, 0.1022239, 0.2904218, 0.06943094, 0.1451103, 
    0.1896995, 0.1040421, 0.08140979, 0.1275409, 0.091546, 0.1082637, 
    0.2117497, 0.411603, 0.1171734, 1.248161e-06, 0.03658693, 0.003090583, 
    0.06327977, 0.08327831, 0.09452424, 0.1202981, 0.3725945, 0.005643016,
  0.01981432, 0.02026314, 0.005899291, 0.1158994, -6.020497e-05, 
    1.811299e-07, 0.01413463, -8.718522e-05, 0.0001004505, 0.03238375, 
    0.12616, 0.09565365, 0.2680855, 0.2812167, 0.2561204, 0.3279469, 
    0.2935175, 0.4140268, 0.2743193, 0.05638522, -2.697443e-05, 0.04901525, 
    0.04613438, 0.02052568, 0.1957838, 0.2706684, 0.3354897, 0.2790401, 
    0.08105347,
  0.02747086, 0.08774652, 0.1203819, 0.04098323, 0.01628617, 0.001478208, 
    0.01477335, 0.1140887, 0.102154, 0.08502878, 0.1095544, 0.1688237, 
    0.1779629, 0.324515, 0.4339414, 0.5395435, 0.5524139, 0.4226874, 
    0.4068637, 0.06693819, 0.1252201, 0.06493202, 0.1085465, 0.1182252, 
    0.143141, 0.2777263, 0.2504531, 0.2704109, 0.2120248,
  0.1654624, 0.07406588, 0.022651, 0.1129243, 0.2014383, 0.08587154, 
    0.05227865, 0.07820438, 0.1772386, 0.144812, 0.2798663, 0.3284567, 
    0.2513307, 0.3310047, 0.370449, 0.3638606, 0.2817351, 0.5176576, 
    0.243045, 0.04694042, 0.03427158, 0.01724634, 0.08290122, 0.1549695, 
    0.2311321, 0.1250569, 0.4628107, 0.4646038, 0.3263848,
  0.500082, 0.3991217, 0.3211527, 0.2416192, 0.3452215, 0.3041481, 0.2056487, 
    0.1141634, 0.07449674, 0.09061018, 0.09635843, 0.1829715, 0.1229214, 
    0.2182928, 0.1084529, 0.2759132, 0.340378, 0.106371, 0.07687321, 
    0.1145181, 0.2347322, 0.3403485, 0.2517251, 0.2540558, 0.06452543, 
    0.1606754, 0.2705972, 0.3498709, 0.5396267,
  0.3863279, 0.3296807, 0.3085337, 0.3758235, 0.439962, 0.3269188, 0.3740159, 
    0.4052768, 0.3715598, 0.3335582, 0.1880533, 0.2069625, 0.2514389, 
    0.4092031, 0.6092361, 0.5120406, 0.4860396, 0.4088188, 0.3914213, 
    0.4632359, 0.3609343, 0.3325834, 0.2935637, 0.2561962, 0.1137414, 
    0.1223256, 0.2011129, 0.3756963, 0.5045509,
  0.2222029, 0.2180355, 0.213868, 0.2097005, 0.205533, 0.2013656, 0.1971981, 
    0.1847755, 0.1860566, 0.1873378, 0.1886189, 0.1899, 0.1911811, 0.1924623, 
    0.1735647, 0.1771201, 0.1806756, 0.184231, 0.1877865, 0.1913419, 
    0.1948973, 0.2364593, 0.2357902, 0.2351211, 0.234452, 0.2337829, 
    0.2331138, 0.2324447, 0.2255369,
  0.2318976, 0.20593, 0.2041296, 0.1770808, 0.08710694, 0.1389757, 0.1635913, 
    0.1188797, 0.02571031, 0.05084629, 0.07100981, 0.1448398, 0.2797875, 
    0.01033765, 0.2412817, 0.2192418, 0.164359, 0.2306807, 0.3244349, 
    0.3457267, 0.5600145, 0.4491504, 0.185285, 0.1253612, 0.1839701, 
    0.226541, 0.2530909, 0.2315379, 0.2940255,
  0.1150409, 0.1776943, 0.3318291, 0.2057775, 0.3013137, 0.3276521, 
    0.2507239, 0.5002797, 0.2584476, 0.2843648, 0.2577741, 0.24572, 
    0.2771985, 0.3020774, 0.3335632, 0.3774855, 0.4534957, 0.5268111, 
    0.4083546, 0.3620604, 0.3793266, 0.3283314, 0.3204988, 0.3348494, 
    0.2179314, 0.1710221, 0.3715791, 0.3530567, 0.1118997,
  0.4227744, 0.4468877, 0.2976053, 0.2921812, 0.3670556, 0.3691815, 
    0.4638175, 0.2861403, 0.2549517, 0.3710238, 0.3524257, 0.3326377, 
    0.3936197, 0.3899947, 0.4948243, 0.4135475, 0.4309711, 0.4289144, 
    0.3965595, 0.3010465, 0.3405074, 0.3047556, 0.2686276, 0.2989867, 
    0.382225, 0.3469934, 0.4095953, 0.3198383, 0.3175738,
  0.3683175, 0.3454005, 0.3562357, 0.3343993, 0.3606499, 0.3546195, 
    0.3819143, 0.2806859, 0.2711652, 0.2233608, 0.2126241, 0.2387395, 
    0.207096, 0.2650837, 0.2808287, 0.3998586, 0.3699877, 0.3382688, 
    0.2807454, 0.3465034, 0.293286, 0.3348389, 0.22549, 0.2779851, 0.1143247, 
    0.2279786, 0.2892062, 0.2752978, 0.3357968,
  0.1230208, 0.1220128, 0.1173253, 0.1147959, 0.1550204, 0.09070586, 
    0.1597916, 0.1888119, 0.1328451, 0.03888597, 0.1342812, 0.1150672, 
    0.04836656, 0.06928465, 0.4220493, 0.1169663, 0.1180791, 0.1407041, 
    0.1225269, 0.09466945, 0.2065262, 0.1598498, 0.1436092, 0.5064467, 
    0.02921307, 0.06099177, 0.1352877, 0.1732495, 0.2171871,
  0.1115346, 0.04971789, 0.02579673, 0.01069199, 0.08539321, 0.119653, 
    0.08126969, 0.05803956, 0.04066574, 0.02453517, 0.002239369, 0.001895837, 
    0.02656065, 0.02019351, 0.04829146, 0.1166098, 0.04256433, 0.03013219, 
    0.06278329, 0.1411388, 0.1419169, 0.08428565, 0.1027989, 0.009964356, 
    0.09053385, 0.06751683, 0.09902139, 0.04736682, 0.03726119,
  0.06903797, -2.643732e-05, -0.0002286971, 0.001818556, 0.01718314, 
    0.01096686, 0.02064299, 0.06035841, 0.08828911, 0.04189118, 7.614407e-05, 
    0.004432652, 0.01225443, 0.03472328, 0.1344683, 0.05961578, 0.0513024, 
    0.05764169, 0.04648125, 0.05813238, 0.02184546, 0.06116731, 0.1269094, 
    0.004404725, 0.1648035, 0.01891046, 0.01083685, 0.01988943, 0.07300016,
  0.2413595, -1.114066e-08, 0.003626375, 0.0810029, 0.0458153, 0.03133877, 
    0.02094551, 0.03954769, 0.03681686, 0.07236019, 0.05708335, 0.03891102, 
    0.1240317, 0.06270853, 0.04479225, 0.05489062, 0.03049508, 0.01364945, 
    0.02052071, 0.007068495, 0.02216934, 0.1159185, 0.3912805, 0.01428878, 
    0.0001052016, 6.817609e-06, 0.003756528, 0.02922281, 0.1155677,
  0.2646653, 0.007216612, 0.02177667, 0.01468298, 0.03891661, 0.0304889, 
    0.04164326, 0.08260836, 0.02865744, 0.03896442, 0.1084549, 0.2694291, 
    0.07043197, 0.02915983, 0.02622569, 0.02183963, 0.06031713, 0.05509403, 
    0.05845316, 0.04186298, 0.07766441, 0.18641, 0.08118324, 0.1537758, 
    0.05195351, 0.03072511, 0.03828554, 0.04769427, 0.08754696,
  0.006648748, 0.0023174, 0.0001094197, 0.000791127, 7.704489e-09, 
    0.007360272, 0.0550582, 0.007890533, 0.00050239, 0.0353839, 0.03952788, 
    0.1309365, 0.06589463, 0.04360753, 0.03103582, 0.03063481, 0.04565366, 
    0.09198355, 0.1110791, 0.1541727, 0.07893877, 0.06340734, 0.1923542, 
    0.0991944, 0.0400105, 0.04922419, 0.1395835, 0.2475505, 0.003224552,
  4.742644e-07, 1.05846e-07, 4.973604e-10, 2.81411e-08, 4.870416e-08, 
    0.1112578, 0.04215746, 0.04609438, 0.1768959, 0.1129396, 0.1061039, 
    0.01380142, 0.01436411, 0.02173924, 0.01510885, 0.01214112, 0.00659209, 
    0.05776984, 0.4344082, 0.21697, 0.06244193, 0.08512253, 0.005614731, 
    0.002183942, 0.01385459, 0.01202222, 0.08286422, 0.1349855, 0.0002094473,
  6.325227e-05, -6.750404e-06, -0.0001625935, 1.040462e-07, 1.870733e-08, 
    2.490594e-08, -0.0002870777, 0.1008379, 0.2725509, 0.07719474, 0.149485, 
    0.1716643, 0.08968002, 0.1245022, 0.2255363, 0.1227844, 0.03693042, 
    0.1436784, 0.2177272, 0.4121889, 7.547068e-07, 0.02536298, 0.001462256, 
    0.1278904, 0.08089159, 0.1261854, 0.06148015, 0.1483559, 0.00551801,
  0.02084155, 0.02241752, 0.003930295, 0.1417927, -0.0001337505, 
    1.565103e-07, 0.0147492, -0.0001128496, 3.295265e-05, 0.03169931, 
    0.1355687, 0.1197322, 0.27209, 0.3865417, 0.3176287, 0.458232, 0.3639856, 
    0.521542, 0.5187348, 0.05502239, 6.416404e-06, 0.0726623, 0.03672125, 
    0.02414376, 0.2315788, 0.314021, 0.3784858, 0.3965862, 0.1391526,
  0.02022701, 0.06824283, 0.09136475, 0.03251191, 0.01190454, 0.001263119, 
    0.01118854, 0.1093555, 0.07634067, 0.07724065, 0.09764189, 0.1401562, 
    0.3045375, 0.4659565, 0.565253, 0.6078196, 0.5596844, 0.4545367, 
    0.4780833, 0.05884314, 0.1213944, 0.05127485, 0.07881463, 0.11204, 
    0.1305513, 0.2806935, 0.2509321, 0.2802947, 0.1841652,
  0.1333659, 0.04358251, 0.01659291, 0.09090573, 0.1831087, 0.0700046, 
    0.04304905, 0.05701908, 0.1564764, 0.1204781, 0.2693314, 0.3173578, 
    0.2443239, 0.331849, 0.4048839, 0.4650666, 0.2668367, 0.4902537, 
    0.239062, 0.03432437, 0.02339648, 0.008807732, 0.06799289, 0.1605041, 
    0.2945221, 0.1299045, 0.4543206, 0.4045145, 0.2666853,
  0.5796655, 0.3646351, 0.2656029, 0.4225129, 0.3205359, 0.3815983, 
    0.2552876, 0.1123965, 0.0780881, 0.06324042, 0.09317738, 0.1656059, 
    0.1133424, 0.2298936, 0.1628208, 0.3779652, 0.3055276, 0.09394482, 
    0.09927282, 0.08751933, 0.1957222, 0.332417, 0.1900948, 0.2633544, 
    0.121437, 0.1370322, 0.2670244, 0.3218841, 0.565952,
  0.4247237, 0.3167108, 0.3415723, 0.6169518, 0.7210967, 0.5885643, 0.520411, 
    0.5165111, 0.3689713, 0.3458876, 0.2689824, 0.3340209, 0.4308183, 
    0.5982999, 0.6201741, 0.4689631, 0.4261298, 0.348376, 0.3529304, 
    0.4433306, 0.3574031, 0.3059118, 0.2894565, 0.2902655, 0.218786, 
    0.1192451, 0.2165911, 0.4007342, 0.5739911,
  0.1960303, 0.1936831, 0.1913359, 0.1889887, 0.1866415, 0.1842943, 
    0.1819471, 0.1829119, 0.1843536, 0.1857954, 0.1872371, 0.1886788, 
    0.1901206, 0.1915623, 0.1582095, 0.1595874, 0.1609653, 0.1623432, 
    0.1637211, 0.165099, 0.166477, 0.2211275, 0.2206551, 0.2201826, 
    0.2197102, 0.2192378, 0.2187653, 0.2182929, 0.197908,
  0.2712145, 0.2228032, 0.2021052, 0.1819871, 0.09971399, 0.1273939, 
    0.169898, 0.1272908, 0.01995039, 0.05495375, 0.0907402, 0.1054149, 
    0.2975349, 0.002468448, 0.2304579, 0.2466204, 0.205939, 0.2414728, 
    0.3211076, 0.3870682, 0.5806128, 0.4445494, 0.1786453, 0.1307033, 
    0.2121005, 0.2769866, 0.252082, 0.2722076, 0.3168874,
  0.1059075, 0.1447619, 0.2914526, 0.1579772, 0.2627217, 0.3297641, 
    0.1610093, 0.4619549, 0.2633024, 0.2694232, 0.2531731, 0.2308681, 
    0.2238733, 0.2705689, 0.3625725, 0.3725033, 0.4509875, 0.5483339, 
    0.3480063, 0.3895798, 0.3445801, 0.319222, 0.3427928, 0.3560713, 0.23237, 
    0.2546282, 0.4004726, 0.3899887, 0.1202046,
  0.4668847, 0.3606678, 0.2243695, 0.2412482, 0.3680498, 0.3343976, 
    0.4039215, 0.2147211, 0.190858, 0.2874082, 0.3057659, 0.310121, 
    0.3767992, 0.4355215, 0.4498138, 0.3877449, 0.4050289, 0.4162003, 
    0.3579762, 0.305025, 0.2822843, 0.2727906, 0.2587515, 0.240666, 
    0.3245479, 0.4025115, 0.4541136, 0.3392963, 0.336373,
  0.3717072, 0.3154872, 0.3584671, 0.3194613, 0.3511429, 0.3836907, 
    0.4044591, 0.2529811, 0.2568479, 0.2197201, 0.1774888, 0.2040814, 
    0.195354, 0.2190399, 0.2728707, 0.347626, 0.3380966, 0.3103352, 
    0.2953956, 0.3017247, 0.2608694, 0.2825664, 0.1934422, 0.265361, 
    0.0844147, 0.1752785, 0.2690077, 0.2717198, 0.3367205,
  0.1118148, 0.08042071, 0.09657475, 0.07723734, 0.1005005, 0.06403241, 
    0.1307332, 0.157066, 0.09250759, 0.02084755, 0.1081398, 0.08539051, 
    0.0246339, 0.05204242, 0.3863949, 0.09492829, 0.09720831, 0.08887953, 
    0.07991893, 0.08146798, 0.1704099, 0.1412451, 0.1090316, 0.5164458, 
    0.01739928, 0.05014496, 0.1364092, 0.1752678, 0.1928945,
  0.04706437, 0.03051282, 0.01735799, 0.003778643, 0.03340853, 0.06485013, 
    0.03714345, 0.02250247, 0.02043821, 0.01762389, 0.002180225, 
    0.0004843594, 0.02723728, 0.01108493, 0.03098715, 0.1052752, 0.03026342, 
    0.02228278, 0.03831034, 0.1009659, 0.1010166, 0.03301702, 0.04364215, 
    0.02555932, 0.08429798, 0.04834924, 0.07366338, 0.0214948, 0.01813963,
  0.08656146, 0.0001194546, -0.0002112224, 0.0006835089, 0.001809044, 
    0.001737464, 0.005634552, 0.02375053, 0.04386663, 0.009013527, 
    -5.309216e-05, 0.001657535, 0.004472149, 0.007859396, 0.09120779, 
    0.02648713, 0.02841734, 0.02902854, 0.01971208, 0.04171981, 0.004631151, 
    0.02235438, 0.04235152, 0.02730099, 0.151773, 0.02117685, 0.001254601, 
    0.005914018, 0.02322667,
  0.1353863, 3.395488e-07, 0.004150951, 0.06157568, 0.02352401, 0.007836302, 
    0.004965919, 0.01177782, 0.01464632, 0.01837607, 0.03619879, 0.01675351, 
    0.100406, 0.02594631, 0.01541359, 0.03216505, 0.008184841, 0.001449631, 
    0.002601906, 0.0004753479, 0.004847309, 0.03218615, 0.2338717, 
    0.003479138, -2.017843e-06, 5.580668e-06, -0.003981632, 0.008123289, 
    0.04335862,
  0.2450411, 0.001737876, 0.01012394, 0.01268692, 0.01314426, 0.005611905, 
    0.00527623, 0.008694258, 0.02793041, 0.0271286, 0.01685219, 0.05040338, 
    0.05127465, 0.01459076, 0.005902505, 0.004720825, 0.007339965, 
    0.009046652, 0.01950858, 0.0101359, 0.03136458, 0.08347506, 0.4423557, 
    0.1041289, 0.02683337, 0.01157336, 0.01546854, 0.009725307, 0.05871905,
  0.003864494, 0.0009403956, 5.840508e-05, 0.00289524, -5.659017e-06, 
    0.0005800395, 0.04341792, 0.0007993673, -0.001021914, 0.007731182, 
    0.005356111, 0.02255538, 0.04129848, 0.02147639, 0.0107561, 0.01297798, 
    0.01990999, 0.04039573, 0.04905718, 0.04511051, 0.03683456, 0.04446091, 
    0.1943604, 0.08241482, 0.01615282, 0.02238716, 0.06792038, 0.2154434, 
    -0.00166889,
  4.140877e-07, 8.933539e-08, 5.130898e-10, 2.575949e-08, 4.775359e-08, 
    0.07783365, 0.02851644, 0.02750718, 0.1805857, 0.1044308, 0.03312732, 
    0.00484735, 0.001942007, 0.00354957, 0.004172815, 0.0008906708, 
    0.0007095021, 0.01595239, 0.1796402, 0.2766783, 0.0739863, 0.08163597, 
    0.0006348099, -0.001022257, 0.002007449, 0.0008486647, 0.02713362, 
    0.04386212, 5.614449e-05,
  4.72319e-05, -0.0001381498, 0.0001485365, -2.071458e-08, 2.113895e-08, 
    2.27879e-08, -0.0008945243, 0.09149987, 0.2595444, 0.06669443, 0.1554574, 
    0.1654788, 0.1119369, 0.1145759, 0.1059077, 0.03373351, 0.005869508, 
    0.07335431, 0.08179355, 0.2798433, 6.135028e-07, 0.01612275, 
    0.0004732364, 0.07224801, 0.06108416, 0.03897849, 0.03721594, 0.04745519, 
    0.01113949,
  0.01654338, 0.02507774, 0.002534091, 0.163754, -0.0001065289, 1.433636e-07, 
    0.01397741, -7.652132e-05, -3.368884e-05, 0.02723861, 0.1221856, 
    0.149251, 0.2928852, 0.4213111, 0.4925691, 0.4568434, 0.5075901, 
    0.4069107, 0.4468065, 0.05032375, 0.0001247518, 0.07907961, 0.03321986, 
    0.06713814, 0.2620349, 0.3515204, 0.3196321, 0.2746236, 0.1902455,
  0.01902684, 0.05277804, 0.07255714, 0.02220801, 0.008520272, 0.000467337, 
    0.009494177, 0.1048928, 0.06005848, 0.07193831, 0.09588239, 0.1409353, 
    0.4724477, 0.5970683, 0.6400509, 0.5962887, 0.5872267, 0.4897712, 
    0.4542823, 0.05708811, 0.109711, 0.03546095, 0.06858394, 0.1049647, 
    0.1279358, 0.2991824, 0.2733141, 0.2851807, 0.1772908,
  0.202989, 0.03518258, 0.01261936, 0.08130872, 0.1616296, 0.06732554, 
    0.03806963, 0.04421519, 0.1452343, 0.1104755, 0.2584076, 0.3069529, 
    0.2351881, 0.3169989, 0.4078649, 0.4557601, 0.2545947, 0.4584581, 
    0.2247451, 0.0265315, 0.01463479, 0.00317521, 0.0854238, 0.1292683, 
    0.248783, 0.1401997, 0.430903, 0.3685984, 0.2377461,
  0.5680269, 0.3508762, 0.2285161, 0.4900202, 0.2646073, 0.2999637, 
    0.2605529, 0.1041434, 0.05921776, 0.03583163, 0.06971163, 0.1158279, 
    0.06937264, 0.2539765, 0.2426859, 0.446445, 0.2820856, 0.1042002, 
    0.1188709, 0.08746754, 0.1697372, 0.2850796, 0.1393918, 0.2448082, 
    0.376751, 0.1160406, 0.1901373, 0.2915469, 0.6284688,
  0.5412253, 0.3338653, 0.4185804, 0.6629045, 0.7416647, 0.6232457, 0.513626, 
    0.474816, 0.2995111, 0.3109961, 0.3417672, 0.4342243, 0.4771684, 
    0.5428665, 0.5266626, 0.4641415, 0.3907296, 0.3621104, 0.3295116, 
    0.3852783, 0.2872177, 0.2887728, 0.2785394, 0.3288034, 0.278734, 
    0.1318296, 0.2127122, 0.4276146, 0.6660934,
  0.1526051, 0.1496233, 0.1466416, 0.1436599, 0.1406782, 0.1376965, 
    0.1347148, 0.1078391, 0.1124558, 0.1170726, 0.1216893, 0.1263061, 
    0.1309228, 0.1355396, 0.1595904, 0.1587391, 0.1578877, 0.1570364, 
    0.1561851, 0.1553338, 0.1544825, 0.1600145, 0.1592308, 0.1584471, 
    0.1576634, 0.1568796, 0.1560959, 0.1553122, 0.1549904,
  0.2593804, 0.2424669, 0.1543769, 0.158666, 0.09859505, 0.09961139, 
    0.1406862, 0.1254791, 0.006604947, 0.01028827, 0.02986073, 0.09836841, 
    0.3037829, -0.000890751, 0.246523, 0.3212341, 0.2941833, 0.275798, 
    0.3222364, 0.4483649, 0.6087831, 0.458378, 0.154358, 0.08469643, 
    0.2150174, 0.2953164, 0.2954083, 0.2848207, 0.305351,
  0.1222793, 0.1283169, 0.2440322, 0.1085128, 0.2225672, 0.3218609, 
    0.1112654, 0.3845989, 0.250578, 0.240038, 0.2433064, 0.2157857, 
    0.1575574, 0.2239884, 0.4002629, 0.4145927, 0.4696614, 0.5218195, 
    0.2893418, 0.3797633, 0.3079052, 0.3252723, 0.3258109, 0.3539447, 
    0.2254728, 0.313331, 0.4182063, 0.4137946, 0.1724153,
  0.452888, 0.2758091, 0.1743799, 0.1918374, 0.3091733, 0.2908791, 0.3462393, 
    0.1825356, 0.1605967, 0.2277126, 0.2503206, 0.2441865, 0.3709723, 
    0.418059, 0.3562286, 0.3448224, 0.3633146, 0.3706152, 0.3226154, 
    0.2692709, 0.2206807, 0.2476516, 0.2446162, 0.2014677, 0.2746074, 
    0.3962047, 0.4425111, 0.3390992, 0.3176424,
  0.3465206, 0.2730984, 0.337448, 0.3093757, 0.3237483, 0.3869866, 0.3933216, 
    0.2038212, 0.2300185, 0.1837517, 0.1453633, 0.1692978, 0.1487282, 
    0.1771942, 0.2534305, 0.3151886, 0.2739068, 0.2514322, 0.2676087, 
    0.274213, 0.2298059, 0.2690309, 0.1404402, 0.2310524, 0.05530437, 
    0.1165068, 0.2175696, 0.2492166, 0.324997,
  0.0895207, 0.04767463, 0.06841269, 0.04569211, 0.05725493, 0.04505533, 
    0.1024839, 0.1200334, 0.05410617, 0.01223306, 0.08449781, 0.05585266, 
    0.01125802, 0.04031074, 0.33285, 0.08198641, 0.08060827, 0.06209366, 
    0.06020643, 0.0792154, 0.1361081, 0.1221645, 0.08011031, 0.5113007, 
    0.009487596, 0.04235841, 0.1178263, 0.1499831, 0.1610738,
  0.02066326, 0.01248476, 0.01681801, 0.00218979, 0.01485688, 0.03811703, 
    0.02058679, 0.01191507, 0.01054463, 0.004367437, 0.00092458, 
    0.0002562791, 0.03721607, 0.004730149, 0.0181032, 0.08363962, 0.02194032, 
    0.01543661, 0.01907736, 0.05984522, 0.05323761, 0.0102043, 0.01681227, 
    0.01928391, 0.0689566, 0.02595741, 0.04482196, 0.009522114, 0.009113637,
  0.05078364, 0.0004374764, -0.0001673296, 0.0003519724, -0.002078905, 
    0.0007803689, 0.001853671, 0.006851905, 0.02457695, 0.002435157, 
    -0.0001149797, 0.0005432948, 0.001555789, 0.002208899, 0.04522219, 
    0.01280213, 0.01460488, 0.01448117, 0.007694366, 0.03161035, 0.00169004, 
    0.009975947, 0.01780313, 0.01931905, 0.1214215, 0.02420013, 0.0002245477, 
    0.003182065, 0.007908306,
  0.06142203, 8.162427e-07, 0.002001371, 0.04918956, 0.01100018, 0.001504194, 
    0.0005568913, 0.00281361, 0.005854015, 0.003038213, 0.02069767, 
    0.008913401, 0.06472171, 0.007477893, 0.001960936, 0.01005006, 
    0.001715133, 0.0001875657, 0.0005022968, 0.0001598355, 0.002133128, 
    0.01213631, 0.1106472, 0.001400071, -1.343619e-05, 4.926585e-06, 
    -0.001043483, 0.002988832, 0.018836,
  0.08652347, 0.0003050476, 0.006747483, 0.008872547, 0.0029801, 0.001683795, 
    0.001549141, 0.002395488, 0.02775044, 0.01278121, 0.002727173, 
    0.01462946, 0.03527439, 0.005154184, 0.001179578, 0.0009016608, 
    0.001932501, 0.002216633, 0.003766033, 0.001407309, 0.003942471, 
    0.02193583, 0.184015, 0.08596777, 0.02232285, 0.0041769, 0.004872439, 
    0.001304894, 0.0109122,
  0.002957461, 0.0008524956, 2.138923e-05, 0.003513717, -7.228343e-07, 
    1.470304e-05, 0.02457617, 0.000156363, -0.0005917446, 0.003034161, 
    0.001341524, 0.005191827, 0.02456835, 0.01050016, 0.0026457, 0.004004651, 
    0.006524434, 0.01480725, 0.02788736, 0.01914719, 0.01475635, 0.01806884, 
    0.222636, 0.07163266, 0.005139209, 0.008328171, 0.0189881, 0.06979328, 
    -0.001958091,
  3.806611e-07, 7.189937e-08, 5.052389e-10, 2.291263e-08, 4.720732e-08, 
    0.02573367, 0.01577892, 0.009570246, 0.1609038, 0.04981368, 0.01861938, 
    0.0005123048, 0.0002180217, 0.000304317, 0.0006487875, 0.0002882896, 
    0.00028783, 0.006239634, 0.0770538, 0.1676515, 0.02678328, 0.07485895, 
    6.419652e-05, -0.001265549, 0.0001581105, 0.0001157457, 0.009988282, 
    0.01885352, 1.585568e-05,
  2.531703e-05, -7.512423e-05, -8.101456e-05, -7.749856e-07, 2.267748e-08, 
    2.131014e-08, -0.0009212205, 0.08117022, 0.2443707, 0.05201593, 
    0.2079236, 0.1917605, 0.0664337, 0.06321518, 0.0477561, 0.01655839, 
    0.002072242, 0.02917156, 0.03579841, 0.1213216, 5.736474e-07, 
    0.008513291, 0.0002401764, 0.0393726, 0.03567749, 0.008985256, 
    0.007949105, 0.01797958, 0.01968523,
  0.01356042, 0.01408327, 0.0008140368, 0.1719247, 5.597587e-06, 
    1.375115e-07, 0.01554231, -0.000124259, -7.698376e-05, 0.02225172, 
    0.119867, 0.1856279, 0.3172556, 0.4154069, 0.4870601, 0.3914501, 
    0.4014726, 0.2742555, 0.2692535, 0.0450562, 0.0007604154, 0.07554542, 
    0.02859269, 0.08802572, 0.1564604, 0.2718806, 0.2097004, 0.1544202, 
    0.1729749,
  0.07047279, 0.04450035, 0.0552569, 0.01208188, 0.003691933, 0.0003803745, 
    0.007506587, 0.1040551, 0.05037682, 0.07221133, 0.09662832, 0.1327404, 
    0.6119422, 0.6851038, 0.6401515, 0.518496, 0.5682933, 0.4887311, 
    0.4038565, 0.05383667, 0.0838571, 0.01901035, 0.0733563, 0.08997889, 
    0.1256619, 0.3023275, 0.2710364, 0.2223977, 0.1661691,
  0.2060831, 0.0279292, 0.01041522, 0.07327408, 0.1385109, 0.06050389, 
    0.0387433, 0.03603942, 0.130692, 0.1043772, 0.2429626, 0.2773681, 
    0.2135008, 0.2827359, 0.3961442, 0.4289987, 0.238359, 0.4218489, 
    0.2024691, 0.01910806, 0.01179403, 0.001149635, 0.09024909, 0.09910408, 
    0.2292064, 0.1208533, 0.367856, 0.3496063, 0.2246978,
  0.5380289, 0.3035844, 0.1937526, 0.3872178, 0.2754024, 0.2793823, 
    0.2105533, 0.08552148, 0.03581513, 0.02201598, 0.05446918, 0.08047508, 
    0.04191254, 0.2466962, 0.2923138, 0.4092539, 0.2284932, 0.1452357, 
    0.1401258, 0.1179392, 0.1319881, 0.234802, 0.1059411, 0.2396117, 
    0.4662955, 0.1056589, 0.1391436, 0.2692322, 0.6438905,
  0.6304194, 0.3221176, 0.4741116, 0.5835451, 0.6748361, 0.5942059, 
    0.4982316, 0.4534838, 0.3263945, 0.348196, 0.4321632, 0.4268278, 
    0.4210896, 0.4422477, 0.483736, 0.4287091, 0.3503895, 0.3477381, 
    0.3558274, 0.3196138, 0.21661, 0.2385557, 0.2091031, 0.333417, 0.253814, 
    0.1265322, 0.1876204, 0.458022, 0.7291385,
  0.03631271, 0.03447295, 0.03263319, 0.03079343, 0.02895366, 0.0271139, 
    0.02527414, 0.03267104, 0.03941876, 0.04616648, 0.05291419, 0.05966191, 
    0.06640963, 0.07315734, 0.08808207, 0.08894461, 0.08980715, 0.0906697, 
    0.09153224, 0.09239478, 0.09325732, 0.1126938, 0.1069233, 0.1011528, 
    0.09538228, 0.08961178, 0.08384129, 0.07807079, 0.03778452,
  0.2502342, 0.1715394, 0.1198653, 0.05652318, 0.05205386, 0.03548114, 
    0.07683668, 0.09185234, 0.01519724, 0.007857192, 0.006318101, 0.06618195, 
    0.2724968, -0.006138749, 0.2907143, 0.3624699, 0.3606655, 0.3041666, 
    0.2993165, 0.4564767, 0.6662856, 0.4982079, 0.1260008, 0.0479546, 
    0.2332661, 0.3755636, 0.3348264, 0.2581276, 0.2911306,
  0.1592126, 0.1176287, 0.2073043, 0.0638145, 0.183974, 0.3010983, 0.0763985, 
    0.2918673, 0.2287332, 0.1997707, 0.2218945, 0.200166, 0.104364, 
    0.1794976, 0.4272461, 0.3933872, 0.4557029, 0.5080245, 0.2357196, 
    0.3203095, 0.2822854, 0.3144751, 0.310621, 0.3493962, 0.2184204, 
    0.3157045, 0.3996856, 0.4257904, 0.2113855,
  0.4129535, 0.1967865, 0.132104, 0.1462482, 0.2531355, 0.2189514, 0.2851116, 
    0.1532197, 0.1228504, 0.1676321, 0.1919951, 0.1847099, 0.3328312, 
    0.3389778, 0.2767994, 0.2930007, 0.3089154, 0.3009492, 0.2854605, 
    0.2239784, 0.1705278, 0.201304, 0.2125278, 0.1618678, 0.2262108, 
    0.3640338, 0.4014704, 0.2996338, 0.2929723,
  0.2868516, 0.2153747, 0.2893229, 0.2615726, 0.2782137, 0.3341166, 
    0.3638284, 0.1614039, 0.1808864, 0.1489295, 0.1085042, 0.1247999, 
    0.09941062, 0.130828, 0.2142238, 0.2611051, 0.1862796, 0.1836998, 
    0.2005274, 0.2275603, 0.1764405, 0.2231492, 0.09753911, 0.1928544, 
    0.03280206, 0.07684734, 0.1724198, 0.2161517, 0.2755003,
  0.06300636, 0.02521822, 0.04681131, 0.02579329, 0.03324334, 0.02967629, 
    0.07071593, 0.09317891, 0.03470838, 0.007634414, 0.05748545, 0.0368761, 
    0.004457177, 0.03025034, 0.277677, 0.06769028, 0.06266114, 0.04301579, 
    0.04537885, 0.07254178, 0.1054078, 0.08950567, 0.05380335, 0.4821029, 
    0.005135154, 0.03340203, 0.08967914, 0.1024229, 0.1340212,
  0.01152028, 0.009038068, 0.01339602, 0.001391071, 0.007772075, 0.02256617, 
    0.01123282, 0.007438656, 0.004974181, 0.001359359, 0.000299008, 
    0.0003765489, 0.03939652, 0.002262421, 0.01082777, 0.06298064, 
    0.01570326, 0.008851679, 0.009128549, 0.02876183, 0.02802093, 
    0.004561325, 0.007605022, 0.01087375, 0.045045, 0.01389728, 0.02052744, 
    0.00410128, 0.00404975,
  0.03209351, 0.002168824, -0.0001155943, 0.0002183055, -0.002400446, 
    0.0004232792, 0.0009184168, 0.003041376, 0.01269588, 0.001205411, 
    -0.0001356875, 0.0002334895, 0.0008570267, 0.001119308, 0.01767365, 
    0.005946045, 0.00671742, 0.00729729, 0.003563971, 0.01687079, 
    0.0008935747, 0.005628407, 0.00998187, 0.01271821, 0.09690117, 
    0.02547856, 0.000108452, 0.001621822, 0.003984497,
  0.03434382, 1.189823e-05, 0.0008408259, 0.03521903, 0.00493782, 
    0.0002980822, 0.0001580766, 0.0007650955, 0.00175596, 0.0007633749, 
    0.01288304, 0.003698285, 0.03599805, 0.001774841, 0.0005879374, 
    0.002843614, 0.0002723004, 9.349138e-05, 0.0002434036, 7.931706e-05, 
    0.001217013, 0.006429912, 0.06199391, 0.0009714662, -4.069214e-05, 
    -4.241579e-07, -0.0006943071, 0.001462761, 0.01007724,
  0.04328295, 0.0001740641, 0.006048506, 0.006872425, 0.0003845294, 
    0.0009393323, 0.0008095799, 0.001180384, 0.02752268, 0.01224951, 
    0.001020541, 0.007407475, 0.01936802, 0.002447822, 0.0005776124, 
    0.0004391741, 0.0009816291, 0.00104099, 0.001618586, 0.0004925173, 
    0.001485409, 0.01003745, 0.08254386, 0.08606014, 0.02368156, 0.001439637, 
    0.006868204, 0.0006143076, 0.003068753,
  0.00214661, 0.0007535103, 5.321627e-06, 0.002467119, 1.026881e-07, 
    5.454688e-06, 0.01130179, 5.002046e-05, -0.0002325874, 0.001631345, 
    0.0006101175, 0.002271248, 0.01311148, 0.006272985, 0.0008209767, 
    0.00115084, 0.001820602, 0.005045699, 0.01669584, 0.01231441, 
    0.008215212, 0.008021902, 0.2084641, 0.06768295, 0.001743737, 
    0.002601888, 0.007106782, 0.03138936, -0.001848726,
  3.603335e-07, 5.825143e-08, 5.037644e-10, 7.381612e-09, 4.68571e-08, 
    0.0113926, 0.006462111, 0.00265879, 0.121994, 0.01717199, 0.007671633, 
    0.000150763, 8.654495e-05, 5.915199e-05, 4.977675e-05, 0.0001500776, 
    0.0001552273, 0.003300209, 0.04046793, 0.09088373, 0.05282519, 
    0.06322081, 2.859864e-05, -0.0009095627, 2.48409e-05, 4.968106e-05, 
    0.004590769, 0.01016205, 4.18895e-06,
  1.108441e-05, -2.497828e-05, 7.451354e-05, -2.972026e-06, 2.380092e-08, 
    2.024828e-08, -0.0008475721, 0.07645969, 0.2257246, 0.03603044, 
    0.2076523, 0.1247626, 0.03565546, 0.02795757, 0.0259378, 0.004606583, 
    0.001107279, 0.01333161, 0.01940807, 0.0657666, 5.206671e-07, 
    0.004255115, 0.0001219994, 0.02341217, 0.02061772, 0.004001204, 
    0.003437373, 0.00978619, 0.02006521,
  0.01084043, 0.005435772, 1.450149e-05, 0.1799316, -5.880501e-05, 
    1.341541e-07, 0.01507627, -0.0001027946, -7.030385e-05, 0.0161435, 
    0.1175449, 0.2476711, 0.3232742, 0.3782605, 0.4401736, 0.3462889, 
    0.3071986, 0.1806489, 0.1555221, 0.03872644, 0.002305411, 0.05938657, 
    0.02280224, 0.08495864, 0.08971494, 0.1847005, 0.1460056, 0.08803434, 
    0.1312748,
  0.08362257, 0.03966889, 0.03623861, 0.007699089, 0.001667655, 1.5503e-05, 
    0.006640219, 0.09332755, 0.04217271, 0.06695607, 0.08859223, 0.1236898, 
    0.6065943, 0.6096421, 0.5600957, 0.42381, 0.4757904, 0.4329408, 
    0.3438199, 0.04754315, 0.06362005, 0.01012831, 0.06418744, 0.07304597, 
    0.1280029, 0.287187, 0.2232265, 0.1797374, 0.1394564,
  0.1437384, 0.02232346, 0.007257718, 0.06001749, 0.1105588, 0.04769584, 
    0.03712927, 0.03147143, 0.10951, 0.09179602, 0.22725, 0.2284135, 
    0.1932617, 0.2478859, 0.3845006, 0.3884301, 0.2154506, 0.3638768, 
    0.1612855, 0.01636876, 0.007964245, 0.0006121587, 0.08644366, 0.07618169, 
    0.1965978, 0.09334596, 0.2892027, 0.2968633, 0.1936248,
  0.5052397, 0.2338132, 0.1641915, 0.3148369, 0.2736497, 0.2575155, 
    0.1786627, 0.05793346, 0.02041809, 0.0132016, 0.03804008, 0.05963266, 
    0.02630858, 0.2101275, 0.2602449, 0.3448993, 0.1603978, 0.1375818, 
    0.1952953, 0.1159711, 0.107207, 0.1997961, 0.07878148, 0.2483686, 
    0.5486171, 0.09449682, 0.1081231, 0.2743005, 0.6643077,
  0.6081298, 0.2810918, 0.4128258, 0.507491, 0.5926959, 0.567609, 0.4669885, 
    0.4313213, 0.3694473, 0.3458111, 0.3484687, 0.3429599, 0.3459107, 
    0.3955192, 0.426409, 0.3762133, 0.3073521, 0.3090223, 0.2889782, 
    0.2614846, 0.1798833, 0.1834434, 0.1556539, 0.2777033, 0.2278674, 
    0.1022279, 0.1612112, 0.4567026, 0.7160791,
  0.01062638, 0.01064972, 0.01067306, 0.01069641, 0.01071975, 0.0107431, 
    0.01076644, 0.02000875, 0.02367327, 0.02733779, 0.03100232, 0.03466684, 
    0.03833136, 0.04199588, 0.0368106, 0.03823692, 0.03966323, 0.04108955, 
    0.04251586, 0.04394218, 0.04536849, 0.04839421, 0.04328002, 0.03816584, 
    0.03305166, 0.02793748, 0.0228233, 0.01770911, 0.0106077,
  0.2399901, 0.1106699, 0.06061837, 0.008312863, 0.005594532, 0.01664037, 
    0.05101831, 0.07636245, 0.01095495, 0.002412777, 0.01361892, 0.0377378, 
    0.1619044, -0.007328079, 0.2969843, 0.395521, 0.3792614, 0.3383735, 
    0.2691089, 0.4609284, 0.7039312, 0.5911913, 0.1026154, 0.02899289, 
    0.2238417, 0.4870495, 0.3606153, 0.2217541, 0.3037285,
  0.1976889, 0.1060927, 0.170306, 0.04243055, 0.1559329, 0.2765448, 
    0.06112684, 0.2054993, 0.1963516, 0.1782125, 0.2019123, 0.1959852, 
    0.06384066, 0.1564614, 0.4247657, 0.3783723, 0.4151296, 0.4509776, 
    0.1717996, 0.2617987, 0.2590286, 0.2602623, 0.2802658, 0.3461244, 
    0.195275, 0.3074663, 0.3824792, 0.4286552, 0.2226906,
  0.3453699, 0.1381315, 0.09644502, 0.108052, 0.190993, 0.1547567, 0.2255265, 
    0.1237426, 0.09104539, 0.1182691, 0.1419657, 0.1352111, 0.2643914, 
    0.2545047, 0.1948596, 0.2232331, 0.2547791, 0.2439354, 0.2370519, 
    0.1678402, 0.1254798, 0.137628, 0.1617596, 0.1218999, 0.1764458, 
    0.3175796, 0.3396047, 0.2594702, 0.2569758,
  0.2309322, 0.1658626, 0.2269757, 0.2203029, 0.2308413, 0.2604994, 
    0.3064169, 0.1279588, 0.1347005, 0.1292081, 0.07283609, 0.08668704, 
    0.05824773, 0.0862591, 0.1612733, 0.1835116, 0.118309, 0.121118, 
    0.1407755, 0.1557214, 0.1177329, 0.1580661, 0.05787163, 0.1725031, 
    0.01875969, 0.04966914, 0.1200219, 0.1741318, 0.2220468,
  0.0400291, 0.01319152, 0.02931182, 0.01399003, 0.01868675, 0.01685551, 
    0.04244601, 0.06720752, 0.02191216, 0.004211864, 0.03278412, 0.02254552, 
    0.002150604, 0.01775334, 0.2228725, 0.04778557, 0.04173218, 0.02394159, 
    0.03168431, 0.0537043, 0.07356968, 0.05860136, 0.03169274, 0.4441503, 
    0.003133662, 0.0211366, 0.06215826, 0.07017749, 0.09351063,
  0.007984274, 0.006720652, 0.008886509, 0.0009766973, 0.004636727, 
    0.01107222, 0.005876102, 0.005275884, 0.002109, 0.0008314133, 
    6.408428e-05, 0.001508503, 0.03639203, 0.001205575, 0.004554989, 
    0.04365307, 0.008607069, 0.004775358, 0.004419982, 0.0119836, 0.01259728, 
    0.002989075, 0.004900501, 0.006172169, 0.03155285, 0.00706933, 
    0.00754558, 0.002375528, 0.002429487,
  0.02026872, 0.003444561, -5.083734e-05, 0.0001514641, -0.002010641, 
    0.0001625149, 0.0005570255, 0.001898289, 0.005092245, 0.0007579047, 
    -0.0001073695, 8.825307e-05, 0.0005704739, 0.0007198307, 0.007456887, 
    0.003666686, 0.002622596, 0.003143615, 0.001616594, 0.007982023, 
    0.0005733151, 0.003762084, 0.006669321, 0.008653636, 0.07481313, 
    0.02607916, 7.104437e-05, 0.001053168, 0.002602319,
  0.02213325, 7.701962e-07, 0.0004982801, 0.02117824, 0.001866542, 
    0.0001393001, 8.443187e-05, 0.0003826992, 0.00070992, 0.0004340933, 
    0.007388388, 0.001282725, 0.01650381, 0.0006189276, 0.0002891752, 
    0.0008030147, 0.0001326375, 5.908151e-05, 0.0001520131, 4.868842e-05, 
    0.0008092719, 0.004148292, 0.04016792, 0.002009932, -2.326112e-05, 
    -7.344141e-07, -0.0003225043, 0.0008737739, 0.006428838,
  0.02677984, 0.0001493861, 0.004267586, 0.005640794, 0.0001993312, 
    0.0006181874, 0.0005362263, 0.0007188476, 0.02336228, 0.01363223, 
    0.0005830201, 0.004534323, 0.00909799, 0.001040991, 0.0003139865, 
    0.000273842, 0.0006119359, 0.0006477569, 0.001006754, 0.0002816261, 
    0.0008151776, 0.006011456, 0.04949236, 0.07759842, 0.03179272, 
    0.0005583005, 0.00531176, 0.0003958948, 0.001605624,
  0.001593255, 0.001871195, 1.093935e-06, 0.002081865, 8.00431e-08, 
    2.897958e-06, 0.006222993, 2.868739e-05, -7.867056e-05, 0.001045151, 
    0.0003605174, 0.001402406, 0.005495445, 0.003366153, 0.0003148603, 
    0.0003299072, 0.0006430598, 0.001709064, 0.008564447, 0.006464338, 
    0.004441437, 0.003179587, 0.1769855, 0.06465723, 0.0005034191, 
    0.0006402864, 0.003391922, 0.016929, -0.0004892382,
  3.464567e-07, 4.94276e-08, 4.967932e-10, 4.557969e-09, 4.655362e-08, 
    0.006486705, 0.001604171, 0.0008944285, 0.09022538, 0.004516008, 
    0.002731198, 8.450338e-05, 5.368065e-05, 3.573203e-05, 1.859815e-05, 
    9.518578e-05, 0.0001014999, 0.002081882, 0.02573519, 0.05503812, 
    0.04111457, 0.05076395, 1.622292e-05, -0.0006953505, 1.198871e-05, 
    3.022534e-05, 0.002639386, 0.006576623, 2.457183e-06,
  1.359309e-06, -1.404495e-05, 4.166325e-05, -2.677939e-06, 2.464432e-08, 
    1.944853e-08, -0.0007808469, 0.07145862, 0.2073419, 0.02311299, 
    0.1534561, 0.05860237, 0.01811785, 0.007835678, 0.009605884, 0.002468657, 
    0.0007173044, 0.008070547, 0.01286733, 0.04307131, 4.728574e-07, 
    0.004652674, 0.0001230222, 0.011818, 0.009891281, 0.002570194, 
    0.002191981, 0.006471367, 0.0168591,
  0.007264956, 0.002424998, -6.247794e-05, 0.1661727, -4.758218e-05, 
    1.319565e-07, 0.01316551, -7.005642e-05, -6.089662e-05, 0.0107255, 
    0.101895, 0.2223627, 0.2802612, 0.3398606, 0.3573225, 0.2735697, 
    0.2226806, 0.1088312, 0.09912799, 0.03475136, 0.00231523, 0.04428764, 
    0.02070099, 0.08459926, 0.04247046, 0.1182082, 0.09052386, 0.05097491, 
    0.09597533,
  0.08070367, 0.02981109, 0.02183067, 0.004588153, 0.001016267, 2.043804e-06, 
    0.005658744, 0.08180334, 0.03610442, 0.05952427, 0.07725099, 0.1092698, 
    0.5309075, 0.4928922, 0.4427108, 0.3425954, 0.3832427, 0.3341472, 
    0.2621314, 0.0436184, 0.04730331, 0.005623456, 0.05163729, 0.05843407, 
    0.1287308, 0.2543052, 0.1608678, 0.1234568, 0.09970775,
  0.08852841, 0.01683131, 0.003745016, 0.04578929, 0.08239227, 0.03544071, 
    0.03356649, 0.02848548, 0.09037764, 0.07205062, 0.203894, 0.1767652, 
    0.1679274, 0.1982595, 0.3182896, 0.3199539, 0.1883801, 0.3061376, 
    0.1159999, 0.01248749, 0.005164144, 0.0004162932, 0.07775678, 0.05778487, 
    0.1542246, 0.07373098, 0.1905091, 0.1966261, 0.1406735,
  0.4055627, 0.1688459, 0.1333493, 0.2657413, 0.2471255, 0.2211643, 
    0.1454526, 0.05739675, 0.01352209, 0.007368417, 0.02756819, 0.04706575, 
    0.0184785, 0.1929156, 0.2285569, 0.2872754, 0.1047123, 0.1345127, 
    0.2037593, 0.1224022, 0.08867937, 0.1644249, 0.05825089, 0.2236303, 
    0.5016701, 0.08074068, 0.08460831, 0.2710252, 0.6160033,
  0.5470926, 0.2506782, 0.3640893, 0.4563481, 0.5291709, 0.494055, 0.3948248, 
    0.3817741, 0.33659, 0.2932537, 0.2776709, 0.2644094, 0.2842138, 
    0.3243818, 0.3291317, 0.2641703, 0.2474368, 0.2331972, 0.2066477, 
    0.2004258, 0.1246151, 0.1408031, 0.1153195, 0.2418214, 0.2026664, 
    0.09034441, 0.1368583, 0.4369822, 0.6402393,
  0.004458392, 0.004630582, 0.004802772, 0.004974963, 0.005147153, 
    0.005319343, 0.005491533, 0.007182681, 0.009828123, 0.01247356, 
    0.01511901, 0.01776445, 0.02040989, 0.02305533, 0.03141491, 0.03199248, 
    0.03257006, 0.03314764, 0.03372522, 0.0343028, 0.03488038, 0.02307826, 
    0.01968305, 0.01628784, 0.01289263, 0.009497422, 0.006102212, 
    0.002707002, 0.00432064,
  0.1668659, 0.076603, 0.01697333, 0.002713199, 0.001662518, 0.007269546, 
    0.02155758, 0.03234916, -0.000997048, 0.001293797, 0.007154775, 
    0.02286125, 0.1295058, -0.005925428, 0.2668709, 0.3779025, 0.3841428, 
    0.3527828, 0.2372941, 0.513034, 0.7124841, 0.645598, 0.08687682, 
    0.02171622, 0.1980895, 0.5153885, 0.4116956, 0.1859092, 0.2239627,
  0.1989592, 0.08326028, 0.1322385, 0.03316769, 0.1319972, 0.2429572, 
    0.05299596, 0.1510089, 0.1662163, 0.1561729, 0.1976988, 0.2030792, 
    0.04625071, 0.1378754, 0.4278743, 0.3534608, 0.3763151, 0.4185066, 
    0.1354383, 0.2308446, 0.2412881, 0.2093199, 0.2478353, 0.3380641, 
    0.1720848, 0.2841646, 0.3384294, 0.3695487, 0.1996204,
  0.2995915, 0.09874357, 0.07771123, 0.08787395, 0.1567811, 0.1211439, 
    0.1822714, 0.09954701, 0.06973036, 0.08746419, 0.1141048, 0.1046315, 
    0.2139611, 0.206714, 0.1405619, 0.1792123, 0.2136188, 0.202913, 
    0.1915677, 0.1317227, 0.09761868, 0.1014672, 0.1238248, 0.09820081, 
    0.1449609, 0.2942135, 0.2876206, 0.2265354, 0.2245763,
  0.1992891, 0.1404645, 0.1901771, 0.189548, 0.1931653, 0.2105967, 0.2534357, 
    0.09851548, 0.1037332, 0.1102474, 0.05285263, 0.06454425, 0.03931783, 
    0.05644628, 0.123318, 0.127498, 0.07428172, 0.07652416, 0.09892621, 
    0.106029, 0.07996187, 0.110924, 0.03815629, 0.1652839, 0.01202896, 
    0.03345271, 0.08798479, 0.1443925, 0.199022,
  0.02460189, 0.008010937, 0.01884813, 0.008958443, 0.009172853, 0.009988271, 
    0.02724453, 0.04746886, 0.01160077, 0.002381015, 0.01749893, 0.01397557, 
    0.001361534, 0.01039847, 0.1839345, 0.02916622, 0.02615188, 0.01448777, 
    0.01824889, 0.03717818, 0.05340712, 0.03654271, 0.01794921, 0.409245, 
    0.002079252, 0.01181152, 0.0417103, 0.04973427, 0.06388164,
  0.006240954, 0.004437834, 0.006299417, 0.0007504989, 0.003436495, 
    0.006246457, 0.004376794, 0.004162948, 0.001123122, 0.0006129989, 
    -1.041812e-05, 0.003905123, 0.03275047, 0.000843759, 0.001973176, 
    0.02460206, 0.004934005, 0.002721438, 0.002731963, 0.006076953, 
    0.006433082, 0.002370096, 0.00373123, 0.004318358, 0.02448917, 
    0.003978047, 0.004034575, 0.001757246, 0.001668244,
  0.01460952, 0.002533979, -2.48433e-05, 0.0001160341, -0.001586509, 
    7.346761e-05, 0.0003919527, 0.001411457, 0.002127841, 0.0005598722, 
    -6.955124e-05, 0.0001230869, 0.0004310856, 0.0005317081, 0.003650548, 
    0.001998294, 0.001254682, 0.00164302, 0.0009493204, 0.004036952, 
    0.0004215442, 0.002842338, 0.004978071, 0.006578106, 0.06018753, 
    0.02259766, 5.361035e-05, 0.0007899784, 0.001926803,
  0.01626746, 4.177958e-07, 0.0003884841, 0.01139996, 0.0008887896, 
    0.0001022766, 5.736663e-05, 0.0002550763, 0.0003865107, 0.0001241214, 
    0.004609317, 0.0005360115, 0.007921755, 0.0003192386, 0.000183997, 
    0.000377962, 0.0001000893, 4.233907e-05, 0.0001102762, 3.465799e-05, 
    0.0006066583, 0.00306114, 0.0297101, 0.003180529, -9.142587e-06, 
    -2.353393e-06, -0.000185977, 0.0006098535, 0.004712737,
  0.01893284, 0.002152975, 0.002660635, 0.004415996, 0.0001333322, 
    0.0004591264, 0.0004045212, 0.0005058903, 0.0200549, 0.01903691, 
    0.0003943418, 0.003047016, 0.004260115, 0.0005380376, 0.000206031, 
    0.0001971968, 0.0004398286, 0.0004636954, 0.0007273552, 0.0002003178, 
    0.0006618599, 0.004247282, 0.03520194, 0.05947654, 0.03798762, 
    0.0002805818, 0.002523572, 0.0002936103, 0.001100041,
  0.001072411, 0.0009738146, 1.925787e-07, 0.004007592, 8.405863e-08, 
    1.926482e-06, 0.005068813, 2.087142e-05, -9.396639e-05, 0.0007614673, 
    0.0002500429, 0.001020293, 0.002203961, 0.001532294, 0.00015542, 
    0.0001350704, 0.0003469003, 0.000946103, 0.004193062, 0.003356659, 
    0.002317762, 0.001470174, 0.1596534, 0.0584741, 0.000232498, 
    0.0002249363, 0.001840062, 0.01050135, 0.002196878,
  3.361421e-07, 4.541338e-08, 4.950378e-10, 3.515402e-09, 4.625378e-08, 
    0.004389649, 9.709372e-05, 0.0004342385, 0.07138798, 0.001335658, 
    0.001450932, 5.792853e-05, 3.936844e-05, 2.53548e-05, 1.049651e-05, 
    6.905645e-05, 7.543165e-05, 0.001507999, 0.0187163, 0.04009725, 
    0.02947278, 0.04085653, 9.802849e-06, -0.0007980612, 7.562298e-06, 
    2.199732e-05, 0.001806962, 0.004813113, 3.222271e-07,
  4.980208e-07, -1.022626e-05, -1.009701e-05, -1.931932e-06, 2.502228e-08, 
    1.883858e-08, -0.0007314546, 0.06935805, 0.1947483, 0.0154136, 
    0.09800681, 0.02920795, 0.009917911, 0.004355303, 0.00547978, 
    0.001671296, 0.0005314213, 0.005750737, 0.009654498, 0.03211483, 
    4.346772e-07, 0.01497571, 0.0003861617, 0.004153103, 0.004380144, 
    0.001902819, 0.001638974, 0.004845091, 0.01383667,
  0.005400712, 0.00156316, -8.347672e-05, 0.1565681, -3.616792e-05, 
    1.304121e-07, 0.01172731, -4.402273e-05, -5.224541e-05, 0.007572643, 
    0.0893557, 0.1801909, 0.2443054, 0.3056663, 0.2957974, 0.218141, 
    0.1547596, 0.07187178, 0.0643898, 0.03548191, 0.002038864, 0.03584375, 
    0.01742714, 0.05508458, 0.02052311, 0.07172663, 0.04427432, 0.02863532, 
    0.07743499,
  0.07196893, 0.02364088, 0.01554807, 0.002581187, 0.0006750469, 
    1.175896e-06, 0.004000857, 0.07527822, 0.03346849, 0.05362491, 
    0.07101513, 0.09751302, 0.4471278, 0.4015172, 0.3444791, 0.2671453, 
    0.3037011, 0.2601447, 0.1722443, 0.0421578, 0.03593589, 0.003202126, 
    0.04609439, 0.05269078, 0.1367662, 0.2123047, 0.1162623, 0.0803048, 
    0.06365444,
  0.05382044, 0.01320041, 0.002012864, 0.03585847, 0.06594068, 0.02767806, 
    0.03403758, 0.03459333, 0.08206421, 0.05802925, 0.1823249, 0.1462487, 
    0.1451952, 0.1616948, 0.2453455, 0.2379364, 0.1662595, 0.2666253, 
    0.08884446, 0.01162974, 0.003861497, -5.26994e-05, 0.07537553, 
    0.04491761, 0.12434, 0.06744067, 0.133122, 0.1272628, 0.09368212,
  0.2964932, 0.110243, 0.1082952, 0.2420136, 0.2027924, 0.2384, 0.1296142, 
    0.05045505, 0.01035579, 0.008629584, 0.02123198, 0.03928706, 0.01459975, 
    0.1687558, 0.2002581, 0.2319828, 0.06704298, 0.1191953, 0.1875689, 
    0.1686874, 0.07297017, 0.1457685, 0.04324029, 0.2075942, 0.4411571, 
    0.07261275, 0.07456144, 0.2458208, 0.5113329,
  0.4554438, 0.2046472, 0.336286, 0.4021608, 0.4133932, 0.4024451, 0.3477412, 
    0.3242908, 0.2827792, 0.2396222, 0.2292114, 0.22505, 0.2404764, 
    0.2678358, 0.2604191, 0.1913929, 0.1904526, 0.1809254, 0.1542412, 
    0.1465935, 0.09036298, 0.1091586, 0.09507272, 0.2084806, 0.1796053, 
    0.07951877, 0.1249054, 0.4074068, 0.5577056,
  0.003017554, 0.003269679, 0.003521804, 0.003773929, 0.004026054, 
    0.004278179, 0.004530305, 0.005539648, 0.007854698, 0.01016975, 
    0.0124848, 0.01479985, 0.0171149, 0.01942995, 0.02458967, 0.02438657, 
    0.02418348, 0.02398038, 0.02377728, 0.02357419, 0.02337109, 0.01147926, 
    0.009115183, 0.006751104, 0.004387026, 0.002022947, -0.000341132, 
    -0.002705211, 0.002815854,
  0.1405581, 0.02841221, 0.008259493, 0.002781287, 0.001928229, 0.004021202, 
    0.008296233, 0.003169439, -0.0001109211, 3.933635e-06, 0.003754944, 
    0.02049392, 0.1186738, -0.004715995, 0.3094224, 0.3027149, 0.3717005, 
    0.383709, 0.2275818, 0.5441142, 0.623857, 0.6699802, 0.09131324, 
    0.02103303, 0.1442847, 0.4683475, 0.3509223, 0.1639349, 0.1168466,
  0.2105114, 0.08210345, 0.1022912, 0.03018046, 0.1217543, 0.2123929, 
    0.04673881, 0.134833, 0.1524008, 0.1525073, 0.180029, 0.2138607, 
    0.0430823, 0.1285481, 0.4097655, 0.3382775, 0.3525541, 0.3929651, 
    0.1183251, 0.2384311, 0.2262792, 0.1917777, 0.2184732, 0.3288572, 
    0.1578879, 0.2448794, 0.3001541, 0.3202177, 0.176942,
  0.2780107, 0.08219033, 0.06856553, 0.0776766, 0.1339355, 0.1047515, 
    0.1615736, 0.08652887, 0.05903213, 0.07117444, 0.09932896, 0.08929724, 
    0.1801971, 0.1778359, 0.1120946, 0.1530924, 0.1863908, 0.1698816, 
    0.1592952, 0.1129596, 0.08184111, 0.08317842, 0.1040449, 0.08335883, 
    0.128989, 0.2787731, 0.2611275, 0.2044911, 0.2101735,
  0.1720848, 0.1209526, 0.1633253, 0.1552625, 0.1624105, 0.1769576, 0.21139, 
    0.07904048, 0.08505742, 0.0937202, 0.04289929, 0.05444399, 0.03079118, 
    0.04193898, 0.09949964, 0.09850167, 0.05493848, 0.05589949, 0.0761046, 
    0.07986479, 0.06052744, 0.08130622, 0.03002294, 0.2000063, 0.009111463, 
    0.02662962, 0.07447983, 0.1189219, 0.1727327,
  0.01739583, 0.006064945, 0.01316162, 0.006805213, 0.006320996, 0.007243844, 
    0.01934484, 0.03615226, 0.008021493, 0.001889075, 0.01109313, 
    0.009471578, 0.00107363, 0.006827906, 0.1746909, 0.01850788, 0.01748648, 
    0.01013426, 0.01243584, 0.02983385, 0.04048691, 0.02723519, 0.0119578, 
    0.4119794, 0.001559704, 0.007268441, 0.03120842, 0.04034632, 0.04560323,
  0.005358462, 0.002910158, 0.005329565, 0.0006320353, 0.002899133, 
    0.003728897, 0.003279007, 0.003591506, 0.0008326305, 0.0004740056, 
    -3.796231e-05, 0.01044983, 0.03718531, 0.0006923236, 0.001174707, 
    0.01190775, 0.003124538, 0.002041186, 0.002150243, 0.004102056, 
    0.004059636, 0.002068723, 0.003161375, 0.003536757, 0.02461465, 
    0.002886411, 0.002784511, 0.001479052, 0.001349184,
  0.01189777, 0.002026398, -2.302616e-05, 9.834718e-05, -0.001547236, 
    5.365663e-05, 0.0003212256, 0.001183815, 0.001343128, 0.000462138, 
    -5.214882e-05, 0.0001210183, 0.0003651496, 0.0004463732, 0.002490058, 
    0.001269707, 0.0008612502, 0.001082797, 0.0007133877, 0.0026797, 
    0.0003496267, 0.002403695, 0.004192945, 0.005463161, 0.07145347, 
    0.02365062, 4.536597e-05, 0.0006609621, 0.001603048,
  0.01338407, 3.409332e-07, 0.0002908311, 0.009485085, 0.0005179953, 
    8.425027e-05, 4.747111e-05, 0.0002069012, 0.0002858433, -0.000653933, 
    0.003408294, 0.0003357922, 0.004953244, 0.0002309504, 0.0001324171, 
    0.0002627888, 8.46381e-05, 3.470657e-05, 9.079199e-05, 2.846447e-05, 
    0.0005110705, 0.002558704, 0.02454978, 0.01414911, -6.260838e-06, 
    -7.622881e-06, -0.0001529001, 0.0004962078, 0.003908471,
  0.015151, 0.0135973, 0.005675669, 0.003871747, 0.0001063754, 0.0003768011, 
    0.0003369142, 0.0004022202, 0.03364874, 0.04927402, 0.0003067934, 
    0.00228554, 0.002670429, 0.0003848898, 0.0001607321, 0.0001600266, 
    0.0003559776, 0.0003890828, 0.0005923392, 0.0001637642, 0.0004839566, 
    0.003426217, 0.02829753, 0.0969943, 0.1005801, 0.0001941687, 0.001475604, 
    0.0002421936, 0.0008394108,
  0.01175622, 0.001582284, -8.06494e-05, 0.004536068, 8.635275e-08, 
    1.68346e-06, 0.02603684, 1.752369e-05, -0.001586214, 0.0006228725, 
    0.0001966714, 0.0007744735, 0.001284715, 0.0008554721, 0.0001105774, 
    9.206618e-05, 0.0002559205, 0.0006864893, 0.002739128, 0.002237041, 
    0.001448843, 0.0009903732, 0.227673, 0.06233914, 0.0001543132, 
    0.0001505748, 0.001234632, 0.007657882, 0.02938983,
  3.29857e-07, 4.439375e-08, 4.936505e-10, 3.488815e-09, 4.588509e-08, 
    0.003417752, -0.0002715809, 0.0003050136, 0.174172, -0.0003636408, 
    0.001028736, 4.640221e-05, 3.28671e-05, 2.123128e-05, 8.027681e-06, 
    5.749997e-05, 6.383276e-05, 0.001256484, 0.01539502, 0.03288063, 
    0.0226746, 0.0364816, 8.790193e-06, -0.001458592, 6.135619e-06, 
    1.858568e-05, 0.001455323, 0.003961991, 2.050063e-07,
  3.804147e-07, -5.433267e-06, -9.934975e-06, -1.281484e-06, 2.554281e-08, 
    1.843995e-08, -0.0007186038, 0.07363603, 0.2089571, 0.01315419, 
    0.06470475, 0.01636456, 0.005083236, 0.003377402, 0.003887071, 
    0.001334194, 0.0004422295, 0.004655226, 0.008069865, 0.02654804, 
    4.305579e-07, 0.08255287, 0.002592022, 0.002529408, 0.002552585, 
    0.001567638, 0.001327248, 0.004063907, 0.01105997,
  0.004996758, 0.0008470035, -0.0002039114, 0.1533888, -3.196661e-05, 
    1.292225e-07, 0.01106457, -3.123553e-05, -4.74005e-05, 0.00606428, 
    0.0961011, 0.1434065, 0.1928249, 0.2441832, 0.2337237, 0.16797, 
    0.1196013, 0.04977577, 0.0493473, 0.03665538, 0.002750679, 0.04774836, 
    0.02975618, 0.03901634, 0.01228936, 0.04384118, 0.02554011, 0.01968053, 
    0.06760237,
  0.06796473, 0.02477218, 0.02217057, 0.002018061, 0.0005140438, 
    1.041733e-06, 0.003322744, 0.07458403, 0.03710933, 0.06368054, 0.1016841, 
    0.1137028, 0.3683307, 0.3381568, 0.2729285, 0.2128663, 0.2443874, 
    0.1964915, 0.1174496, 0.05008734, 0.03072576, 0.002758193, 0.06476478, 
    0.08499544, 0.1328484, 0.1637985, 0.09140338, 0.05785311, 0.04686978,
  0.03923964, 0.01645529, 0.001831145, 0.04171127, 0.07393464, 0.03340146, 
    0.05640963, 0.04384588, 0.09877767, 0.07334047, 0.191863, 0.143915, 
    0.1299966, 0.1503162, 0.199438, 0.1933662, 0.1703782, 0.2553463, 
    0.08441395, 0.01587328, 0.006775334, -0.0007322153, 0.06500507, 
    0.03664976, 0.1015212, 0.06137997, 0.09942629, 0.09389903, 0.06530111,
  0.2270249, 0.08838384, 0.09534353, 0.2063411, 0.1631427, 0.2576028, 
    0.1416224, 0.05864801, 0.007887312, 0.01837253, 0.01927982, 0.03580821, 
    0.01143143, 0.1501885, 0.1906544, 0.2019027, 0.04809208, 0.1043288, 
    0.1807214, 0.2316919, 0.06328169, 0.1358707, 0.03365656, 0.2035079, 
    0.4049662, 0.0708416, 0.07053322, 0.214373, 0.3991133,
  0.3958412, 0.1728949, 0.3133538, 0.3650075, 0.3390494, 0.3563282, 
    0.3036958, 0.2889712, 0.2448274, 0.2093019, 0.2050455, 0.1991396, 
    0.2125453, 0.2275724, 0.2225054, 0.1567714, 0.1579712, 0.1499866, 
    0.1255176, 0.1170085, 0.07344926, 0.09363155, 0.08331665, 0.1880608, 
    0.166206, 0.07543266, 0.1271988, 0.3825663, 0.4928276,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -2.08573e-05, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.0004435529, 0, 0, 0, 6.121424e-05, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.912622e-05, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -0.0001238291, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0.0004643498, 0.000677878, 0, 0, 0, 0.001622323, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, -3.349386e-05, 0.001592889, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.0006604705, 0, 0, 0, 0, 0, -0.0001417488, 
    2.90029e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -5.131907e-05, 3.501876e-05, 0, 0, 
    0.00059015, 0, 0, -1.101328e-05, 0.002721648, 0.003048449, -6.649791e-06, 
    -6.603955e-06, -7.97432e-07, 0, 0, -3.136976e-06, 0,
  0, 0, 0, 0, 0, 0, 0.002915208, 0.0006142465, -1.022567e-06, 0, 0, 
    0.003425351, 0, -7.49586e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0006420799, 0, 
    -4.810146e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, -0.0001416677, 0.003541244, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.002428566, 0, 0, -4.725392e-06, 0, -5.40324e-05, 
    -0.0001701074, 1.610616e-05, -5.751279e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.682674e-06, -1.184458e-06, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.000215163, 0.0005011387, 
    -1.967132e-05, 8.329836e-05, 0.002240462, -3.377849e-05, 0.0003607585, 
    0.001941241, 0.004653485, 0.01130533, -2.754105e-05, -6.603955e-06, 
    -2.99638e-06, -4.005085e-05, 0, 0.0006234038, 0.001816469,
  0, 0, 0, 0, 0, 0, 0.007581248, 0.001566333, 4.309223e-05, 0, -5.0755e-05, 
    0.005199347, 0.0002060963, 0.0003089726, 0, 0, 0, 0, 0, 0, 1.788749e-05, 
    -3.571498e-05, 0, 0.002711772, -1.359397e-05, -0.0001726285, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, -0.0003016456, 0.005291833, 0.000877107, 
    -4.596034e-06, -1.975442e-07, -1.173943e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -8.630892e-09, 0, 0.0001286545, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -7.779681e-05, 0.003621532, 0, 0, -6.47877e-05, 0, 
    -0.0002431457, 0.0004441621, 0.002297871, 6.147196e-05, -3.303764e-07, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, -2.554857e-05, 0, 0, 0, 0.0003582514, 0, 0, 0, 4.964995e-06, 
    1.718611e-05, -5.086169e-06, 0, 0, 0, 0, 0, 0, 0, -3.121268e-05, 
    -8.72064e-06, 0, 0, 0, 0,
  7.605973e-08, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001593217, 0.0006844338, 
    0.0006735165, 0.0001675453, 0.004101374, 5.060917e-05, 0.00288607, 
    0.006844465, 0.01742383, 0.0185699, -0.0001939459, 2.55823e-05, 
    -1.850495e-05, -8.736997e-05, 5.854917e-05, 0.001386891, 0.004006988,
  0, 0, 0, 0, 0, 0.0009638776, 0.0198428, 0.00258436, 0.0001461742, 
    -7.56073e-06, 0.0006220129, 0.01477378, 0.001352288, 0.0004168396, 0, 0, 
    0, 0, 0, 0, -6.402816e-05, 0.0001831606, 0, 0.006829421, 0.0003709875, 
    0.0002857991, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, -0.0007060029, 0.00831639, 0.002748947, 0.0003194331, 
    -1.66872e-06, -6.701962e-05, 7.685828e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 1.523721e-05, -4.697094e-08, -2.886929e-06, 
    -3.022211e-05, 0.006237626, -4.904509e-05, 0, 0, 0, 0, 0, 0, 0, 
    -9.180073e-06, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -2.200271e-05, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.005636784, 0, -1.200552e-05, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -0.0003468261, 0.0067828, 0, 0, 0.0006831763, 0, 
    0.002419814, 0.01484131, 0.007563019, 0.0004928212, -3.730347e-05, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, -3.832286e-05, 2.141793e-05, 0, 2.121699e-06, 0.001741472, 
    1.419685e-05, 0.0008362332, 0.001378368, -0.0001139671, 6.824431e-05, 
    -1.693113e-05, 0, 0, 0, 0, 0, 0, 0, 0.0006180982, 0.002922812, 0, 0, 0, 0,
  5.324181e-07, 0, 0.0004587585, -2.782251e-05, 0, 0, 0, 0, 0, -1.387612e-05, 
    0, -4.848861e-07, 0.004201767, 0.0007584423, 0.001235979, 0.003777902, 
    0.00598207, 0.0007411257, 0.005944678, 0.01083896, 0.02884186, 
    0.03428793, -0.0004756982, 0.0001428415, -0.0001487916, -0.000113955, 
    0.0007266556, 0.00753145, 0.006754105,
  0, 0, 0, 0, 0, 0.00348895, 0.04679144, 0.007421579, 0.003596738, 
    -7.441319e-05, 0.001751236, 0.01813001, 0.004547527, 0.002429716, 0, 0, 
    0, 0, 0, 0, -0.0001064253, 9.180554e-05, 0, 0.01259935, 0.002375253, 
    0.0001986399, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0.0007438473, 0.0004863449, 0.01463552, 0.005997476, 
    0.004268813, -1.087418e-06, 0.005553497, 0.0008422485, 0, 0, 0, 0, 0, 0, 
    -1.454842e-05, 0, 0.0003934949, 0.0008354677, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, -9.90342e-06, 7.39149e-05, -3.342099e-05, 
    0.0009453935, 0.0007585337, 0.01668103, 0.0008373871, 0, 0, 0, 0, 0, 0, 
    0, -9.297172e-05, 0, -9.68017e-06, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -0.0001637418, -0.0001027821, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -4.226983e-06, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -1.608025e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.007854547, 0, 0.0002172451, 
    -5.433183e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, -1.434429e-05, 0, 0.0007335976, 0.016017, -1.639378e-05, 0, 
    0.002425072, 0, 0.01377828, 0.03226017, 0.01475029, 0.001838023, 
    -5.669313e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, -2.904764e-05, 0, 0, 0, -4.366711e-05, 0.0009931655, 0, -2.700737e-05, 
    0.004745517, 0.0003592172, 0.00257229, 0.003127361, -0.0003302463, 
    0.0001470424, -2.405021e-05, 0, 0, 0, 0, 0, 0, 0, 0.002829052, 
    0.006251966, 0, -1.56103e-06, 0, 0,
  0.0006048518, 0.001462602, 0.002060748, -3.773267e-05, 0, 0, 0, 
    -4.197095e-05, -1.69873e-06, 0.0001568547, 0, -3.974562e-05, 0.008922727, 
    0.005682665, 0.002519635, 0.01444062, 0.008871127, 0.001202696, 
    0.01331414, 0.019714, 0.04971024, 0.06461467, -0.0007244641, 
    0.0002463511, -0.0002445152, 0.003298548, 0.001126761, 0.01938085, 
    0.01015721,
  0, 0, 0, 0, 0, 0.008987835, 0.08022439, 0.01290472, 0.01312429, 
    -0.0002521987, 0.005388435, 0.0233742, 0.01084006, 0.003614706, 0, 0, 0, 
    0, 0, 0, -0.0001368582, 0.000295191, -1.890815e-05, 0.01502162, 
    0.01059646, 0.0008221456, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0.005511924, 0.005203702, 0.02327517, 0.01239684, 
    0.01057106, 2.235959e-05, 0.0165892, 0.008828486, -2.628498e-05, 0, 0, 0, 
    0, 0, -5.726315e-05, 0.0003647766, 0.0005997496, 0.00425744, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -7.57919e-08, 0, -4.19707e-05, 0.002698408, 0.001308594, 
    0.01260622, 0.004688414, 0.03111674, 0.009628069, -7.935451e-06, 0, 0, 0, 
    0, 0, 0, 0.001136727, 0.002600565, 5.972878e-05, -1.601668e-06, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -2.214232e-05, 0, -1.945215e-05, 0.0008337646, 
    0, 0, 2.255599e-05, 0, -1.955789e-05, 0, 0, 0, 0.003872095, 0.001384703, 
    0, -2.651458e-06, 0.000225636, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.396189e-06, 0, -9.957324e-06, 
    0.0007213526, 0, 0, 0, 0, 0, 0, -1.682709e-06, 0, 0, -5.952722e-06, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3.29308e-05, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.375929e-05, 0, 
    0, 0, 0, 0, 0, 0, 0.0003428445, 0.0002683227,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.526141e-05, 
    0.001363028, 0.001545964, 0, 0, 0, 0, 0.004313108, 0.005704949, 
    0.0003729496, -1.330131e-05, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.00618264, 0.0006532831, 
    0.003878991, 0.002384491, 0.002072323, 0, 0, 0, 0, 0, 0, -6.728457e-07, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.408813e-06, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, -1.058174e-05, 0, 0.006077385, 0.03854096, 0.0003017756, 
    -2.265625e-05, 0.0084068, 0, 0.02425112, 0.06870996, 0.03065561, 
    0.002610384, 0.0007827704, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0.002182414, -4.412774e-06, 0, 0, -5.976918e-05, 0.0009937368, 
    -4.431478e-06, 0.0004076021, 0.008299894, 0.004425444, 0.007446827, 
    0.003737112, -0.0004694949, 0.001375042, -0.0001137462, 0, 0, 0, 0, 0, 0, 
    0, 0.005750711, 0.009205342, 0, -2.645337e-05, 0, 0,
  0.002796699, 0.002876814, 0.003704374, 1.223352e-05, 0, 0, -2.978469e-06, 
    0.001647224, -4.80058e-05, 0.0007649277, 8.0408e-05, 0.001653829, 
    0.02562844, 0.01403505, 0.006510208, 0.0222488, 0.009914196, 0.004330523, 
    0.02517579, 0.03252378, 0.0947549, 0.09906323, 0.005102586, 0.001011282, 
    0.001717641, 0.01661612, 0.004084523, 0.03508941, 0.02015326,
  0, 0, 0, -1.760634e-06, -7.922865e-06, 0.01288488, 0.1151081, 0.02079787, 
    0.05104603, 0.002639827, 0.02392977, 0.03894066, 0.0252736, 0.009310601, 
    0, 0, 0, 0, 0, 0, 0.004840312, 0.002235497, -0.0002031774, 0.0269495, 
    0.01287473, 0.002270761, -2.723263e-05, 0, 0,
  0, 0, 0, 0, 0, 0, 0.01250999, 0.01078598, 0.03939299, 0.02627433, 
    0.01654383, 0.001432519, 0.02945731, 0.01993215, 8.111203e-05, 
    -5.415185e-06, 0, 0, 0, 0, 5.706489e-05, 0.001582337, 0.005344361, 
    0.00953502, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -7.525625e-06, 0, -0.000155359, 0.008681728, 0.01174374, 
    0.02628808, 0.01044793, 0.05161625, 0.04105971, -5.71038e-05, 
    0.001138464, 0, 0, 0, 0, 0, 0.0031048, 0.009961697, 0.001115552, 
    -1.513007e-05, 0, 0, 0,
  0, 2.442264e-05, 3.99778e-05, 0, 0, 0.0003094027, 0, 0, -4.980815e-06, 
    -8.485223e-06, 1.510731e-06, 0.001871783, 0.007545867, -1.212866e-05, 
    0.001980075, 0.001417587, -1.292069e-06, 0.00184513, 0, 0, -7.26208e-06, 
    0.006669871, 0.006752629, -4.744556e-05, 0.0005522565, 0.002149539, 0, 
    0.002026208, -5.028807e-06,
  0.0002684105, 2.685616e-06, -9.931145e-06, 0, 0, -5.868028e-07, 
    0.002346341, 0, 0, -0.0001642388, 0.0002009289, -5.861109e-05, 
    0.00154919, 0.001141418, 2.477901e-05, -4.603668e-05, 0, 0, 0, 0, 
    -0.0001579746, 0, -0.0001263506, 5.774403e-05, 0, 0, 0, -4.414583e-10, 0,
  0, 0, 0, -3.527447e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -1.599118e-10, -1.148276e-09, 5.151595e-09, -1.353742e-09, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.001492191, 0, 0, 0, 0, 0,
  0, -5.435111e-05, 0, -9.345007e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -1.186001e-05, 0, 0, 0.001710085, 0.0008546427, 0, 0, 0, 0, 0, 0, 
    0.003240663, 0.0004745509,
  0, 0, 0, 0, 6.091267e-05, -8.058401e-06, 0, 0, 0, 0, 0, 0, 0, 0.0003777973, 
    -1.764287e-05, 0, 3.07615e-05, 0.0001010711, 0.002920715, 0.01280782, 
    0.0008038798, 0, 0, 0, 0.006451823, 0.00903589, 0.006146447, 
    -0.0001946328, -7.111855e-06,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -4.221562e-06, 0.005520219, 
    0.01200182, 0.01123323, 0.00639553, 0.01243305, 0, 0, 0, 0, 0, 
    -1.275056e-05, -3.430522e-05, 0, 0, 0,
  0, 0, 0, -1.887237e-15, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.780519e-05, 
    0.0004367465, 0.002994751, 0.0005034914, -6.36391e-07, 0, 0, 0, 
    3.425011e-06, 0, 8.626762e-05, 0, 0, 0, -1.41214e-08, 0,
  0, 0, 0, 0, 1.472839e-06, 0, 0.02298186, 0.06382738, 0.0004429449, 
    -0.0005241127, 0.01345349, 0.0003263458, 0.03303751, 0.1087293, 
    0.05785885, 0.004976762, 0.003794695, 0, 0, 0, -5.740073e-09, 
    2.23647e-07, -3.918101e-08, -3.584595e-08, 0, 0, 0, 0, 0,
  0, 0.004511734, -3.384215e-05, 0, 0, 0.0001964995, 0.0007642015, 
    0.007443905, 0.005379611, 0.03474208, 0.01433496, 0.0206526, 0.01503971, 
    0.005391449, 0.0198905, 0.0007451492, 0, 0, -5.876091e-05, -1.634404e-05, 
    -1.148042e-07, 1.059025e-07, 1.597883e-05, 0.02348281, 0.01212192, 
    -5.897552e-05, -7.649438e-05, 7.195355e-10, -6.137828e-06,
  0.009751162, 0.005390513, 0.008292072, 0.001832071, 1.466971e-05, 
    7.818234e-05, 0.0006472624, 0.005359909, 0.001889989, 0.003259574, 
    0.0007376142, 0.01062556, 0.08483591, 0.05464529, 0.02360227, 0.03636405, 
    0.01142758, 0.01611877, 0.04068403, 0.04956703, 0.1734788, 0.1443557, 
    0.04052465, 0.003492648, 0.006867643, 0.02605223, 0.007239462, 
    0.07242996, 0.03593424,
  0, 0, -6.050281e-08, 0.001241921, 0.004042187, 0.04660746, 0.1704895, 
    0.1164332, 0.09562414, 0.01186357, 0.05756716, 0.06160316, 0.0626891, 
    0.02818833, 2.509412e-05, -1.051787e-05, -4.254801e-10, 0, 0, 
    -4.534696e-06, 0.01526559, 0.005648731, 0.0004681596, 0.04146853, 
    0.02243077, 0.004871143, -0.000113883, -1.427747e-06, 0,
  0, 0, 0, 0, 0, 1.154413e-08, 0.04802991, 0.01772884, 0.04824506, 0.1079939, 
    0.02759744, 0.01594291, 0.06925968, 0.03438391, 0.0001691211, 
    -1.704923e-05, 0, 0, 0, 0, -3.8708e-05, 0.01256098, 0.02296718, 
    0.03722911, -1.57571e-05, 0, 0, 0, 0,
  0.0002765236, 0, 0, 0, 5.71403e-08, 4.648894e-05, -2.558922e-05, 
    0.0002618879, 0.01083614, 0.03477227, 0.02767849, 0.04512867, 0.01385889, 
    0.08543812, 0.06788854, 0.0003676054, 0.001778516, 0, 0, 0, 0, 
    -1.048567e-05, 0.01429769, 0.01276829, 0.003726234, 0.001860879, 
    2.669742e-06, 0, 0,
  0, 0.005027556, 0.002419941, 0, 0, 0.0006963979, -2.63762e-05, 
    0.0002120322, 0.0007691957, 0.009114967, 0.002627439, 0.01293788, 
    0.03030017, 0.004491362, 0.009783087, 0.004637339, 0.004674583, 
    0.008303777, -2.622039e-05, 0, 0.003184245, 0.01740507, 0.01497764, 
    -0.0001405297, 0.01158713, 0.003389056, 0.0001066258, 0.007452771, 
    0.001460919,
  0.004545779, 0.005594894, -0.0002029182, 0, 0, -0.0001601491, 0.004732183, 
    0, 0.00341228, 0.003326361, 0.002163541, -3.8735e-05, 0.008295386, 
    0.009808261, 0.0006138359, 0.001436543, 0, 0, 0, -7.471001e-06, 
    0.001299881, -0.0001422686, 0.006308041, 0.007749846, 0.001277255, 
    8.613311e-05, 0.001839279, -0.000143446, 0.0005868882,
  0, -3.443101e-08, -4.283067e-07, -0.0001321082, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, -0.0001215254, 0, 0, -2.669935e-09, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5.150781e-10, 5.009015e-08, -7.146801e-09, 2.872472e-08, -4.083745e-11, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -1.430114e-05, 0.003662582, 0, 0, 0, 0, 0,
  0, 0.00419991, -2.059607e-06, 0.001323947, 0, 6.939741e-05, 0, 0, 
    -2.078261e-05, -1.017351e-05, 0, 0, 0, 0, 0, 0, 7.003628e-06, 0, 
    -0.00011497, 0.00258607, 0.003302654, -2.411262e-05, -1.219409e-05, 
    0.0008860102, 0, 0, 0, 0.004020773, 0.000607584,
  8.416443e-05, 0.0002342194, -1.03465e-05, -1.251614e-05, 0.005935765, 
    -0.0001041541, 0, 0, 0, 0, 0, -6.09721e-06, -4.838238e-07, 0.001812953, 
    0.00056509, -0.0001822903, 0.0007047099, 0.003541367, 0.01054604, 
    0.03754288, 0.006868365, -3.644933e-05, 0.0004194795, -7.469418e-06, 
    0.009316093, 0.01194391, 0.01062382, 0.0011042, 0.003066011,
  0, 0, 0, 0, 2.343695e-11, -4.484675e-07, 0, 0, 0, 0, 0, 2.443393e-09, 0, 
    -3.025096e-07, 0.02015465, 0.02743149, 0.0282771, 0.01730309, 0.03185924, 
    0.0001278604, -2.75892e-05, 0, 1.568907e-05, 0, -1.574995e-05, 
    0.00104513, 0, -3.165381e-05, 3.483297e-05,
  6.263612e-06, 3.067944e-08, 0, 8.764345e-07, 2.557093e-10, 0, -1.95812e-08, 
    8.559137e-05, 0, 0, 0, -1.048191e-10, -2.652808e-08, 0.001052993, 
    0.009824723, 0.01803716, 0.008225475, -2.331115e-05, 0.00102175, 0, 
    9.853743e-08, 0.0006829296, 1.321966e-05, 0.002912127, -4.766226e-08, 
    -2.810643e-08, 0, -4.93145e-10, 0,
  4.148047e-10, -7.281238e-08, -3.890783e-07, -2.864992e-10, 3.783957e-05, 
    4.019767e-06, 0.03796852, 0.109145, 0.006209565, 0.0002616828, 
    0.01400766, -0.0002284363, 0.07160328, 0.1977202, 0.1720355, 0.005765029, 
    0.009779488, 0, 0, -1.551956e-06, -4.768157e-05, 9.15788e-05, 
    -5.351156e-06, -4.671424e-06, -4.782836e-07, -4.895636e-12, 
    -4.351698e-11, -2.226608e-06, 0,
  9.286989e-06, 0.01649311, 0.007012088, 0, -5.291193e-09, 0.005694798, 
    0.002487782, 0.03651817, 0.04076369, 0.0678587, 0.1050018, 0.09895854, 
    0.07209305, 0.05966174, 0.08693268, 0.01624614, -1.932608e-06, 
    1.550249e-06, 0.001366592, 0.008967, 0.0009033549, 0.02053179, 
    0.005070772, 0.04789591, 0.01718169, -0.0001502217, 0.001385103, 
    6.467132e-05, 7.405829e-05,
  0.05553514, 0.02241351, 0.01787604, 0.00745387, -0.000589609, 0.007254991, 
    0.06919427, 0.4462243, 0.2126997, 0.2173202, 0.2306844, 0.1657173, 
    0.2307243, 0.1626211, 0.1972085, 0.0935538, 0.01117756, 0.03838786, 
    0.08539084, 0.1197234, 0.3163446, 0.280722, 0.1223041, 0.02460786, 
    0.01620933, 0.04135617, 0.01708629, 0.1295935, 0.06815537,
  1.558749e-07, 1.054543e-05, 0.001439662, 0.03150296, 0.1419351, 0.2463429, 
    0.3688657, 0.2578535, 0.4278274, 0.1491183, 0.2402719, 0.1641224, 
    0.272913, 0.05832208, 0.0001940141, 0.0007777802, 7.063107e-06, 
    -7.491436e-08, 1.250446e-07, 0.006617845, 0.1451482, 0.04185823, 
    0.02679699, 0.095443, 0.034619, 0.0163184, 1.496886e-05, -2.723303e-06, 
    -4.312985e-08,
  0, 0, -9.920775e-10, 1.3052e-05, 0.000449486, -2.002539e-06, 0.0438107, 
    0.04003511, 0.0649347, 0.1201849, 0.1199841, 0.1438043, 0.2282945, 
    0.09250618, 0.002097071, 0.006130859, 0.000460481, 1.087631e-06, 
    -2.010792e-07, 2.012867e-05, 0.001736879, 0.1128791, 0.2562814, 
    0.1403117, 0.0004217577, -2.557777e-09, 3.577124e-07, -1.38338e-11, 0,
  0.000214625, -2.731897e-06, 0, -1.55126e-11, 1.259926e-07, 0.001150908, 
    0.0006058729, 0.007752475, 0.09803123, 0.09377296, 0.1204278, 0.1198506, 
    0.1079415, 0.1393913, 0.1044723, 0.02473164, 0.009174019, 5.965298e-05, 
    1.211887e-05, 0, -2.331883e-05, 0.0002051657, 0.0278736, 0.08111083, 
    0.02388392, 0.005868416, 0.002115912, 0.0007533773, 0,
  0.001212697, 0.01197765, 0.004367162, 0, -6.716068e-05, 0.002679928, 
    0.000165828, 0.006870979, 0.005394918, 0.02406337, 0.02358331, 
    0.05521561, 0.07143739, 0.01441864, 0.02133395, 0.0120675, 0.01152587, 
    0.01909648, -0.0001965115, -8.41924e-06, 0.01328555, 0.03017772, 
    0.02263998, 0.00252294, 0.02384357, 0.009361706, 0.006470053, 0.02397877, 
    0.01215972,
  0.006310558, 0.008697505, 0.003810201, 0, 0.00111561, 0.0007338018, 
    0.004995447, 0.000454777, 0.006852536, 0.01059101, 0.0122245, 
    0.004963052, 0.01409633, 0.01417219, 0.002600793, 0.002883058, 0, 0, 
    -8.205838e-05, 0.0002088996, 0.002648745, -0.0002999836, 0.01248302, 
    0.01244457, 0.006786427, 0.005324722, 0.004135535, -0.0003350386, 
    0.01482208,
  0, -7.831605e-05, 0.0004304107, 0.0020997, -6.651097e-05, -1.126462e-05, 
    -1.98782e-05, 0, 0.0003381848, 0.002512157, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.007109818, 0, -1.899552e-05, -1.35405e-09, 0, 0, -3.166731e-06, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001448811, -2.08164e-06, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, -1.93582e-09, -1.017851e-07, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0001880128, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, -5.252089e-06, 0, 0, 0, 0, 0, 1.213791e-06, 0, -1.948738e-06, 0, 
    0.002039846, 0, 0.0006203714, -1.256145e-05, 0, 0, 0, 0, 0.0003925815, 
    0.0004504228, 0.00461737, 0, 0, 0, 0, 0,
  0.004579911, 0.008028606, -5.576441e-05, 0.004329955, -7.628751e-05, 
    0.004308409, -5.884845e-05, -7.33344e-05, 0.002214872, -0.0002387599, 
    -4.798358e-05, 0.003034576, 0.002725251, 0, 0, -1.98769e-06, 
    0.0004917877, 6.020509e-05, 5.626137e-06, 0.007729494, 0.01183355, 
    0.000426321, -1.472287e-05, 0.004024049, -4.018843e-05, 0.0002189911, 
    1.821904e-05, 0.005896931, 0.004933977,
  0.005887028, 0.005330077, -3.408947e-05, -9.425681e-05, 0.01076835, 
    0.00372261, 0.005816538, 0.001122263, -3.709973e-06, -2.888814e-08, 
    5.618644e-05, -4.304465e-05, -1.932632e-05, 0.005494828, 0.003918914, 
    0.003576689, 0.009125569, 0.01610098, 0.02778322, 0.06095067, 0.02533492, 
    -1.955149e-05, 0.00376226, 0.001704908, 0.01458176, 0.01285873, 
    0.02145997, 0.006993323, 0.009660401,
  8.365309e-06, 6.48843e-08, -1.94016e-07, -5.3337e-09, -4.266234e-07, 
    -0.0001219303, 0, -2.52766e-09, 3.417175e-07, 7.541838e-07, 3.153848e-06, 
    3.241606e-06, -5.634409e-09, 3.588256e-07, 0.05538518, 0.05812757, 
    0.05400438, 0.03430817, 0.06752162, 0.01052287, 3.852196e-05, 
    -5.827765e-07, 0.000203272, 0.005466194, 0.002530699, 0.007655304, 
    0.0008250413, 1.597099e-05, 0.005729448,
  1.536098e-05, 2.626755e-06, 1.204313e-06, -6.394445e-08, -1.255915e-09, 
    -9.861946e-09, 0.005339348, 0.001961869, 1.373105e-05, 2.64843e-06, 
    1.132127e-08, 1.020121e-06, 3.054231e-07, 0.02701653, 0.0784795, 
    0.06424128, 0.0343833, 0.0115566, 0.0008370269, -1.634653e-07, 
    8.072922e-06, 0.008015214, 0.0001294804, 0.01073824, 0.0001179942, 
    -3.203584e-06, 0.0008876117, 1.155374e-05, 1.316607e-05,
  2.832354e-06, 0.007583587, 8.546854e-06, 5.976039e-06, 0.01562002, 
    0.001705501, 0.09189446, 0.2017468, 0.01405474, 0.005196899, 0.02034594, 
    0.001452622, 0.129833, 0.2320645, 0.215516, 0.03771288, 0.01111366, 
    -5.718314e-07, 2.544724e-06, 0.0002805395, 1.031356e-05, 0.0188454, 
    0.004253461, 0.007365779, -3.990214e-05, 0.00203308, 3.606215e-05, 
    0.000324426, 3.758921e-06,
  0.03748845, 0.2671829, 0.170454, 0.0008388732, 4.462659e-05, 0.0849415, 
    0.1864319, 0.339883, 0.3245735, 0.2185961, 0.1216291, 0.1292086, 
    0.1519056, 0.07417732, 0.09251121, 0.01594501, 0.000445212, 
    -3.714105e-06, 0.001122808, 0.06245655, 0.06370303, 0.09572682, 
    0.1351821, 0.2011944, 0.07119793, 0.001900591, 0.01197011, 0.04101146, 
    0.007578847,
  0.3947739, 0.3590686, 0.2192216, 0.01750047, 0.0149795, 0.07787184, 
    0.1899941, 0.3988047, 0.1788905, 0.204088, 0.1573748, 0.1026792, 
    0.2097854, 0.1607302, 0.2320214, 0.1063489, 0.03061651, 0.06997296, 
    0.1055489, 0.1309204, 0.3682782, 0.3713637, 0.3759577, 0.1509304, 
    0.06249424, 0.1124849, 0.1004858, 0.3308101, 0.3544974,
  2.323702e-05, 0.007523951, 0.004101448, 0.02029651, 0.1017709, 0.2385262, 
    0.3373469, 0.2025088, 0.3776726, 0.1036434, 0.1760869, 0.1245893, 
    0.2482311, 0.1295734, 0.1551284, 0.1144699, 0.0004463344, 1.565904e-05, 
    4.747678e-05, 0.01105453, 0.08489695, 0.04588574, 0.05117101, 0.1289324, 
    0.2211833, 0.03726102, 0.001641502, 0.008726953, -0.0001008789,
  3.574678e-06, 0, -2.430139e-09, 4.852057e-06, 0.0001521215, -5.442061e-06, 
    0.04110208, 0.07758266, 0.1476264, 0.1037745, 0.08958955, 0.1110974, 
    0.2069321, 0.225637, 0.06160065, 0.003576702, 0.05553194, 0.004761329, 
    8.515596e-05, 0.002870244, 0.04355338, 0.1233028, 0.2548648, 0.2996334, 
    0.1033469, 0.03429925, 0.001277828, 0.002136994, 1.549354e-08,
  0.007629293, 0.006636272, -4.549075e-07, -1.636985e-10, -1.194211e-05, 
    0.003143256, 0.01147342, 0.06455718, 0.1576315, 0.1629832, 0.2471694, 
    0.2002355, 0.1957794, 0.2734084, 0.2741509, 0.1458597, 0.05485924, 
    0.0300768, 0.03007716, -2.49503e-05, 0.0005211203, 0.05273303, 
    0.08345903, 0.1654493, 0.1988572, 0.1103565, 0.03957454, 0.02094856, 
    0.006741796,
  0.005878384, 0.02235326, 0.006168073, -7.921415e-06, 0.01147882, 
    0.005976485, 0.001773123, 0.01072647, 0.01441556, 0.05927031, 0.1253577, 
    0.1726345, 0.1579501, 0.0710184, 0.1014001, 0.09346894, 0.04662934, 
    0.08043037, 0.05486077, 0.004248251, 0.01734812, 0.05302988, 0.04437499, 
    0.05090431, 0.05075309, 0.0637309, 0.0782534, 0.08371753, 0.03782991,
  0.009095863, 0.01372595, 0.01163165, -5.158912e-06, 0.0008590707, 
    0.000467239, 0.009868667, 0.002089693, 0.0118951, 0.02552047, 0.03871946, 
    0.04501943, 0.08443271, 0.05870217, 0.03258301, 0.00733517, 
    -0.0002312225, -5.19842e-05, 0.002663293, 0.002388245, 0.006593308, 
    -0.000347107, 0.02180792, 0.01795788, 0.06639627, 0.057463, 0.0231601, 
    0.00464123, 0.02706254,
  -1.796467e-05, 0.003306275, 0.006604193, 0.006887539, 0.001945873, 
    -0.0001319114, 0.0004344354, 0.003153173, 0.001267491, 0.007087413, 
    0.002441778, 0, 0, 0.0005408186, -2.796514e-05, 0, 0, 0, 0, 0, 
    0.01329942, -8.051841e-06, -0.0009651793, 0.002183543, -2.350791e-05, 0, 
    0.0005710895, -2.080657e-05, 0.001394189,
  0, -6.263701e-07, 3.378603e-09, -0.0003428017, -2.351282e-05, 0, 0, 0, 
    -0.0005659902, 0.004914476, -0.0001388956, 0, 0.001322473, -0.0001545098, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, -4.78032e-11, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.03174e-06, 0, 0, 
    0.002474098, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, -2.657928e-05, 0, 0, 0, -5.651579e-07, 0.0009974035, 
    -5.881589e-05, -1.194545e-05, -7.640051e-05, 0, 0.004219931, 
    2.891457e-05, 0.001677501, 6.975675e-05, -3.701003e-05, 0, -1.068729e-05, 
    0, 0.0007620797, 0.002704072, 0.009285058, 0, 0, 0, 0, 0,
  0.02745637, 0.01860982, 0.0001901525, 0.009395375, 0.002083459, 0.00703895, 
    0.0004501945, -0.0001502229, 0.003960542, 0.003954269, 0.005109174, 
    0.004258879, 0.007811178, -7.213283e-05, 0.003567488, -9.333817e-05, 
    0.005994217, 0.002828107, 0.006581161, 0.01299886, 0.02164825, 
    0.008176616, 0.00875861, 0.01097575, 0.0005135277, 0.0006859069, 
    0.001542515, 0.007090656, 0.0181288,
  0.01514581, 0.006187401, 0.0002809716, -2.35411e-05, 0.01354624, 
    0.01025967, 0.008331305, 0.003262563, 0.000163896, -1.120704e-05, 
    0.003089485, 0.0008675287, 4.283013e-06, 0.01364643, 0.01032564, 
    0.01356052, 0.03128001, 0.04969564, 0.06819261, 0.1113995, 0.05276987, 
    0.01626489, 0.02407364, 0.01623267, 0.03272049, 0.02247164, 0.03886504, 
    0.02755905, 0.02225642,
  0.001002838, 0.0002287387, -3.6451e-05, 3.187678e-06, 2.041245e-05, 
    1.801783e-05, 6.723629e-06, -4.283726e-06, 0.001322846, 0.0002566261, 
    7.490512e-06, 0.0001257843, -6.281299e-05, 0.0005301289, 0.08802254, 
    0.08139398, 0.09360155, 0.06980706, 0.1314572, 0.04450502, 0.04215836, 
    0.01575787, 6.579402e-05, 0.001403576, 0.01370427, 0.02356129, 
    0.01072318, 0.002274375, 0.01690974,
  3.808583e-06, 6.845538e-07, 1.952016e-06, 0.0002222974, -2.010981e-08, 
    1.257305e-09, 0.0006034364, 0.001012024, 1.275929e-06, 1.394244e-06, 
    1.406965e-08, 1.613521e-07, 2.226094e-07, 0.03380833, 0.05879025, 
    0.1060566, 0.04054293, 0.01589064, 0.00615924, 4.212272e-05, 
    7.104942e-06, 0.000239342, 2.769371e-05, 0.001691875, 4.279471e-05, 
    0.0001778818, 2.493581e-05, 4.02893e-06, 4.052217e-06,
  2.460908e-06, 0.0001532197, 6.86106e-06, 9.055872e-07, 0.006181324, 
    0.0002933087, 0.05396677, 0.1797334, 0.006393299, 0.006025302, 
    0.01685845, 0.0003211364, 0.09916634, 0.1901642, 0.1688246, 0.02406281, 
    0.00644541, 5.22687e-06, 3.856068e-07, 1.463116e-05, 5.030046e-06, 
    0.0006236069, 0.0008213413, 0.004495937, 3.180523e-06, 7.741112e-05, 
    1.771521e-06, 3.413636e-05, 7.603963e-07,
  0.007517306, 0.2036119, 0.07871979, 0.0001814531, 4.365026e-05, 0.03952978, 
    0.07056283, 0.2592414, 0.2803788, 0.1827422, 0.06928755, 0.09304417, 
    0.1104889, 0.05482878, 0.07102013, 0.009421199, 0.0002477676, 
    9.343347e-05, -0.0001361429, 0.004251075, 0.009286977, 0.06367639, 
    0.04679739, 0.1836074, 0.05743746, 0.0007356466, 0.0005517533, 
    0.01335863, 0.0001988768,
  0.3155177, 0.3191514, 0.1553192, 0.08851133, 0.01128154, 0.03570143, 
    0.09809894, 0.2537044, 0.1368263, 0.1074348, 0.06432286, 0.06094566, 
    0.160362, 0.137285, 0.1658548, 0.08698714, 0.01906954, 0.04425651, 
    0.07801235, 0.1029276, 0.3717965, 0.3086772, 0.3083025, 0.108042, 
    0.04656782, 0.0765653, 0.07744659, 0.2858696, 0.3167114,
  0.001782272, 0.007385977, 0.006492018, 0.01022633, 0.06531943, 0.185225, 
    0.3339942, 0.1661309, 0.3621107, 0.07299244, 0.1470831, 0.1077619, 
    0.2343942, 0.1142774, 0.1256256, 0.07846513, 9.974375e-05, 7.054752e-06, 
    1.25212e-05, 0.01427625, 0.04454412, 0.02836324, 0.02902224, 0.08639783, 
    0.171245, 0.02552198, 0.01057597, 0.007840762, -4.397329e-05,
  0.001993112, 0, -3.857946e-09, 0.001515736, 0.0001062166, -3.560174e-06, 
    0.06539638, 0.2038377, 0.1926186, 0.09361464, 0.07892032, 0.1090142, 
    0.1701833, 0.1797518, 0.04622228, 0.03384563, 0.03545287, 0.004325713, 
    0.0005390296, 0.000113616, 0.03939035, 0.07785494, 0.2037452, 0.2785721, 
    0.08834137, 0.04318007, 0.001523587, 0.001440757, -8.225875e-06,
  0.05725993, 0.02190083, 0.001433784, 8.441503e-10, -6.119108e-05, 
    0.006934084, 0.0238998, 0.1047221, 0.2078088, 0.1812549, 0.29484, 
    0.154252, 0.152964, 0.2607175, 0.2881523, 0.2001965, 0.1236938, 
    0.06594252, 0.01435747, 0.001558791, 0.008474397, 0.03731209, 0.07590098, 
    0.1317487, 0.1923191, 0.1965304, 0.06112758, 0.03113526, 0.01635652,
  0.1259205, 0.08094262, 0.05938564, 0.0257536, 0.08647574, 0.1055614, 
    0.06041428, 0.0177877, 0.02798039, 0.1805774, 0.2066633, 0.1758012, 
    0.174842, 0.1218707, 0.162177, 0.1463026, 0.1341652, 0.181877, 0.1267688, 
    0.04929297, 0.1274832, 0.1285741, 0.08498409, 0.0830358, 0.06793295, 
    0.08575097, 0.1240894, 0.1768472, 0.149232,
  0.08424623, 0.0433647, 0.1138222, 0.05606613, 0.1070521, 0.1268649, 
    0.06922437, 0.02937474, 0.03280764, 0.1032197, 0.2011487, 0.1551372, 
    0.1181944, 0.110642, 0.08665529, 0.03591001, -0.0003742666, 0.0002777281, 
    0.01314437, 0.005397231, 0.03173522, 0.05154603, 0.05170799, 0.0368165, 
    0.1089602, 0.07558336, 0.03938823, 0.03036305, 0.07703713,
  0.0003917409, 0.03154358, 0.06105084, 0.0844404, 0.02606751, 0.009669418, 
    -1.778885e-05, 0.005195853, 0.004955668, 0.02629294, 0.01646705, 
    0.01749541, 0.02063206, 0.02251335, -0.0008623828, -4.802977e-05, 0, 
    -6.564794e-05, -1.512224e-06, -2.879354e-05, 0.01862951, -2.026125e-05, 
    -0.001450517, 0.006963371, 0.008385429, 0, 0.002135236, 0.002484975, 
    0.006139377,
  0, 3.742496e-05, 0.001285809, 0.001282351, -7.342732e-05, 0, 0, 
    -7.428036e-06, -0.001086847, 0.006508603, 0.002652129, -6.354484e-05, 
    0.001952072, 0.006813371, 0.008284842, 0.001418774, 0, 0, 0, 0, 0, 
    2.760139e-08, 0, -1.756157e-07, 3.202536e-07, 0, 0, -1.844783e-07, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, -2.319662e-05, 0, 0, 0, 0, 0, 0, -3.298945e-05, 
    -5.737038e-05, -0.0001271502, -6.266681e-06, 0, 0.002899113, 0.004771505, 
    0, 0, 0, 0, 0, 0, 0,
  0, -8.195708e-06, 1.785078e-05, -9.016212e-05, 0.0001727665, 0, 0, 
    0.0006977103, 0.0009379614, -4.065885e-05, 0.001822162, -0.0001719961, 
    6.983255e-05, 0.006034998, 0.00344559, 0.005358589, 0.001420337, 
    -0.0001285771, 0, 0.0001070245, -7.362483e-05, 0.003096949, 0.01158918, 
    0.01554657, -2.687113e-05, 0, -1.270094e-05, 0.003274133, 0,
  0.04705479, 0.04018208, 0.007717132, 0.01922842, 0.009255496, 0.01107319, 
    0.001471321, 0.002999273, 0.007166768, 0.02057602, 0.02290251, 
    0.007777618, 0.00964307, 0.0005203864, 0.008339448, 0.006125345, 
    0.01290752, 0.01585643, 0.03287202, 0.03275568, 0.06086305, 0.04892958, 
    0.02980398, 0.03520028, 0.008650445, 0.002241183, 0.008157454, 
    0.01688289, 0.03934277,
  0.05392625, 0.02976936, 0.008043155, 0.03282603, 0.02957723, 0.02447281, 
    0.01725695, 0.009948558, 0.004501201, 0.001731621, 0.02347249, 
    0.00951566, 0.01193545, 0.01946693, 0.01690012, 0.03029498, 0.09409289, 
    0.102775, 0.09836922, 0.1818054, 0.1434813, 0.08460823, 0.08062733, 
    0.04836695, 0.08224358, 0.08919472, 0.09128976, 0.09561219, 0.1024653,
  0.01351238, 0.005140553, 0.001436653, 0.001524786, 0.0006374866, 
    0.002785749, 0.0006338324, -1.780444e-05, 3.575631e-05, 1.885428e-05, 
    4.713665e-05, 0.002060828, 0.004342628, 0.006859228, 0.1016112, 
    0.08944301, 0.0974305, 0.1080663, 0.1746608, 0.1003515, 0.04401618, 
    0.01779138, 0.01381997, 0.01176803, 0.007924771, 0.0284522, 0.02223857, 
    0.02795255, 0.0493781,
  8.542975e-07, 3.65047e-07, 7.788742e-07, 0.005499272, -8.159426e-06, 
    1.077995e-07, -0.0001407084, 0.0003873602, 1.026322e-06, 4.094689e-07, 
    3.153153e-08, 7.094168e-08, 9.090552e-08, 0.05512284, 0.0505528, 
    0.09311493, 0.05106111, 0.01271019, 0.006555687, -1.016145e-07, 
    1.906703e-06, 6.003631e-06, 5.678612e-06, 0.0006827486, 4.437446e-05, 
    0.0008365241, 1.236397e-06, -1.551617e-05, 1.392247e-06,
  6.445931e-07, 1.661294e-05, 1.613996e-06, 5.499704e-07, 0.003457102, 
    0.0004462426, 0.04773825, 0.1942762, 0.004375643, 0.006826229, 
    0.01675184, 0.0006217127, 0.07861855, 0.1696443, 0.1511076, 0.02485914, 
    0.005202022, 3.680069e-06, 1.494127e-08, 1.006006e-06, 2.305761e-06, 
    3.243984e-05, 0.006893686, 0.0005700495, 1.00179e-06, 2.418155e-05, 
    3.114749e-07, 3.041844e-06, 1.61913e-07,
  0.001311368, 0.1651032, 0.04162667, 0.0002217346, 0.0002535541, 0.028146, 
    0.03615895, 0.1709257, 0.2554125, 0.1798684, 0.05267099, 0.07680728, 
    0.093917, 0.05891871, 0.06223699, 0.01091617, 0.0005988384, 
    -6.267269e-05, -9.321543e-05, 5.998856e-06, 0.00617046, 0.02731491, 
    0.004767782, 0.165323, 0.04548896, 0.002016621, -4.920501e-05, 
    0.001265027, 1.085233e-05,
  0.269225, 0.3002715, 0.1379626, 0.06664744, 0.007588502, 0.0259766, 
    0.0606948, 0.1069791, 0.1124071, 0.05912533, 0.02108822, 0.05448167, 
    0.1271776, 0.1211912, 0.1208784, 0.0820494, 0.02337889, 0.0411041, 
    0.06596342, 0.1074631, 0.3806211, 0.2786266, 0.2671883, 0.08763378, 
    0.04760393, 0.06719066, 0.07267129, 0.264557, 0.3090827,
  9.053486e-05, 0.00146766, 0.005881486, 0.005210464, 0.05498218, 0.1491559, 
    0.3306468, 0.1261761, 0.3268594, 0.05835986, 0.1161343, 0.09392153, 
    0.1925364, 0.1113897, 0.08009644, 0.05901684, 0.0006026079, 1.601496e-05, 
    6.761842e-05, 0.01608814, 0.03386385, 0.02770467, 0.02403848, 0.07419422, 
    0.1103654, 0.02141042, 0.01277542, 0.007714315, 0.0001797518,
  0.01361179, 0, -3.773491e-09, 3.029784e-05, 1.654025e-05, -1.666248e-06, 
    0.06258995, 0.1725268, 0.1863522, 0.09188485, 0.07094637, 0.0945494, 
    0.1648988, 0.190105, 0.02709736, 0.02977569, 0.01987961, 0.004343816, 
    0.002064303, 0.0001131775, 0.04072903, 0.07587397, 0.1551026, 0.260681, 
    0.08305801, 0.02266855, 2.110048e-05, 8.330453e-05, 5.770225e-05,
  0.04183884, 0.01782026, 0.003284748, -4.009334e-08, 0.0008140823, 0.01049, 
    0.03640786, 0.1300269, 0.2167794, 0.1731259, 0.2634065, 0.1412203, 
    0.1388926, 0.2420932, 0.2855885, 0.1650696, 0.1054899, 0.07604742, 
    0.002099362, -1.72583e-05, 0.01355402, 0.01492399, 0.07121634, 0.1125415, 
    0.1561961, 0.1895176, 0.04714618, 0.02511068, 0.01663445,
  0.122198, 0.1417644, 0.1020946, 0.04610759, 0.06636819, 0.1182521, 
    0.09476316, 0.05484515, 0.1449083, 0.2377678, 0.1689689, 0.1580961, 
    0.164017, 0.07703799, 0.1556334, 0.139343, 0.1374017, 0.1952242, 
    0.1422232, 0.08586735, 0.1310563, 0.112715, 0.08990432, 0.1334102, 
    0.08539464, 0.09768722, 0.1065245, 0.1490684, 0.1262429,
  0.135538, 0.1261342, 0.1352975, 0.06958617, 0.1091716, 0.1017116, 
    0.1280879, 0.04920292, 0.1036718, 0.1596251, 0.2279661, 0.1837442, 
    0.1311636, 0.1690578, 0.10016, 0.1042281, 0.05896207, 0.05433414, 
    0.0549442, 0.07510538, 0.2057728, 0.164508, 0.1957394, 0.1116889, 
    0.1493619, 0.1037951, 0.06701297, 0.07220253, 0.1460941,
  0.052496, 0.1216572, 0.1535384, 0.198246, 0.1139937, 0.07973861, 
    0.05932871, 0.1232272, 0.05047567, 0.1841948, 0.07681325, 0.06587196, 
    0.1495544, 0.1103235, 0.0837532, 0.05381755, 0.04910396, 0.02279703, 
    0.02946487, 0.01814083, 0.0508802, 0.02682984, 0.01351401, 0.01906371, 
    0.06607809, -0.0001806316, 0.003218504, 0.1236527, 0.05806329,
  0.003202979, 0.004550732, 0.06347543, 0.03420147, 0.0170469, 0.01617826, 
    0.0166686, 0.02277423, 0.01241051, 0.05877667, 0.04536276, 0.0472257, 
    0.02645389, 0.02649988, 0.02993097, 0.03798303, 0.03737523, 0.021621, 
    0.0285719, 0.001594982, -0.0005908431, -0.0003488681, -1.729815e-07, 
    -0.0006381088, 7.570105e-06, -1.559616e-05, -0.0004116142, -0.001135558, 
    0.01685322,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -8.038148e-05, 
    0.000431561, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, -0.0001888294, 0, 0, 0, 0, 0, 0, 0.002648276, 
    0.001193938, 0.001189634, 1.591836e-05, 0, 0.01430177, 0.008690385, 
    -3.393114e-06, 0, 0, 0, 0, 0, 0,
  -0.0001578178, 0.009238054, 0.02308191, 0.009153379, 0.001923483, 
    0.0001921786, 0, 0.002692953, 0.002488704, 0.002848126, 0.01155722, 
    0.006338918, 0.0002391857, 0.006190367, 0.006587724, 0.013934, 
    0.004924493, 0.001554579, 0.0009342707, 0.003519784, 0.005429738, 
    0.02016444, 0.01807554, 0.02252709, 0.002625648, 0, 0.0001625835, 
    0.007963328, 2.667635e-06,
  0.1219015, 0.1575766, 0.1160399, 0.1462627, 0.0872601, 0.04114626, 
    0.01572651, 0.01180879, 0.01931916, 0.03589394, 0.03709284, 0.03067682, 
    0.02401714, 0.003722935, 0.0102267, 0.02969899, 0.05217901, 0.0664951, 
    0.07483272, 0.09688623, 0.1416837, 0.09205824, 0.08551899, 0.06701383, 
    0.04326467, 0.04423729, 0.05839035, 0.05843206, 0.1166417,
  0.1741042, 0.08162662, 0.07131872, 0.05058098, 0.05204464, 0.075525, 
    0.08582354, 0.05328937, 0.04064821, 0.05361448, 0.05650054, 0.03862015, 
    0.01718796, 0.02061773, 0.02107308, 0.04008611, 0.1097812, 0.1710609, 
    0.1634234, 0.2274583, 0.1726138, 0.1233004, 0.1242208, 0.07860934, 
    0.1388026, 0.1463448, 0.1747333, 0.1810144, 0.1976656,
  0.01750788, 0.008362403, 0.006676947, -9.638216e-05, 0.0102294, 
    0.009113099, 0.0005930389, 0.001306155, -5.35711e-05, 5.041092e-06, 
    0.002869906, 0.01033366, 0.01533954, 0.02807616, 0.11491, 0.09465554, 
    0.1078011, 0.1103493, 0.1757897, 0.0898439, 0.04287807, 0.01028304, 
    0.01034066, 0.007360069, 0.01069436, 0.0409168, 0.01063489, 0.03917184, 
    0.04860893,
  1.280261e-07, 1.079088e-07, 3.289709e-07, 0.00622153, 2.51997e-05, 
    -1.660025e-05, -4.706447e-05, 0.0002129931, 5.945672e-06, 3.686524e-08, 
    3.0582e-08, 2.728883e-07, 2.690107e-08, 0.07244475, 0.05681472, 
    0.07575966, 0.05371576, 0.01027958, 0.003637985, -5.82869e-08, 
    2.20012e-07, 3.765495e-07, 7.933708e-07, 3.55828e-06, 0.0001870805, 
    0.0007275819, 6.13389e-08, 0.0002926912, 4.600717e-07,
  2.074628e-07, 6.435705e-06, 3.227179e-07, -2.533521e-06, 0.003229038, 
    0.0002397956, 0.04985172, 0.1945857, 0.01270352, 0.008259087, 0.01775147, 
    0.001432695, 0.07157842, 0.1500452, 0.132513, 0.02235538, 0.004946269, 
    7.212344e-05, 5.207516e-08, 4.62452e-07, 2.636024e-06, 3.823102e-06, 
    0.00340387, 0.0004401966, 1.314768e-06, 7.858594e-06, 3.183417e-07, 
    2.359132e-06, 2.76281e-07,
  6.176768e-05, 0.1394894, 0.02433805, 0.0001039868, 0.0002954323, 
    0.01764587, 0.02125147, 0.0931382, 0.1984494, 0.1617279, 0.0380519, 
    0.05835586, 0.07899781, 0.05750535, 0.06188215, 0.02094645, 0.0006811846, 
    -4.809272e-06, -0.0001306715, -5.381456e-05, 0.002518009, 0.003859627, 
    0.005529063, 0.1445076, 0.03591121, 0.002483233, 0.0001150149, 
    0.0003310755, 3.307461e-06,
  0.2055299, 0.2432757, 0.1006723, 0.05484711, 0.01048498, 0.01386334, 
    0.05010783, 0.04062768, 0.1058047, 0.0426328, 0.01117495, 0.03879507, 
    0.09045924, 0.1034822, 0.08730678, 0.07037609, 0.02527093, 0.03539554, 
    0.0642932, 0.1124079, 0.379903, 0.2454778, 0.209133, 0.06199644, 
    0.04133962, 0.06043955, 0.06021002, 0.244265, 0.2744556,
  0.002111974, 4.942434e-05, 0.0009846499, 0.01478833, 0.05920804, 0.1123327, 
    0.3278881, 0.1076682, 0.2760901, 0.03783942, 0.09401616, 0.08318377, 
    0.1576739, 0.1145061, 0.05062278, 0.03757598, 5.067688e-05, 2.141496e-05, 
    6.443264e-05, 0.01660022, 0.03057902, 0.02640935, 0.01648351, 0.0715498, 
    0.05951956, 0.02177898, 0.002958922, 0.008604039, 0.0007813173,
  0.01631881, -7.449129e-08, 1.941128e-08, 5.066233e-06, 1.325629e-05, 
    -1.253964e-05, 0.06435328, 0.1501515, 0.1554973, 0.08963825, 0.06034916, 
    0.05796685, 0.1475865, 0.1794911, 0.03453149, 0.04107371, 0.008780429, 
    -4.815812e-06, 0.005232643, 5.283404e-05, 0.04822818, 0.05999671, 
    0.1140332, 0.2528623, 0.07485983, 0.01145515, 0.003752831, 3.695986e-05, 
    0.001912129,
  0.02454443, 0.01165838, 0.001369144, -1.556486e-06, 0.006079561, 
    0.01329186, 0.1073554, 0.1402229, 0.2066148, 0.141359, 0.2471662, 
    0.148175, 0.1457542, 0.2402745, 0.2907848, 0.1293786, 0.09387036, 
    0.07772914, 0.001342867, 0.0007619458, 0.0118508, 0.01522989, 0.06974401, 
    0.1022776, 0.1444189, 0.1554061, 0.04520865, 0.02067139, 0.01517816,
  0.1055439, 0.1354026, 0.06143657, 0.02961363, 0.04724026, 0.09432957, 
    0.08638364, 0.1069188, 0.183951, 0.1991559, 0.137925, 0.1482685, 
    0.1616181, 0.04456879, 0.1404159, 0.1259272, 0.1308349, 0.18588, 
    0.1370748, 0.08450893, 0.1006253, 0.0859502, 0.07877076, 0.1294465, 
    0.09360054, 0.1049547, 0.1019825, 0.1241599, 0.1161695,
  0.1748487, 0.178956, 0.1238224, 0.064527, 0.07612132, 0.08704954, 
    0.1599299, 0.1320384, 0.1291686, 0.1293448, 0.2314174, 0.1824571, 
    0.1710676, 0.1679022, 0.1003669, 0.1837478, 0.1435366, 0.1713998, 
    0.1576143, 0.1267206, 0.2376349, 0.1985987, 0.2239734, 0.1614331, 
    0.2254995, 0.1654996, 0.07624351, 0.1320876, 0.2057652,
  0.1437299, 0.1939118, 0.2600379, 0.2483473, 0.1665842, 0.1330135, 
    0.1347055, 0.1801305, 0.1862776, 0.2209587, 0.1425271, 0.1350455, 
    0.160182, 0.1471951, 0.1522082, 0.1791167, 0.1721254, 0.0960355, 
    0.122674, 0.09929895, 0.1562288, 0.06857374, 0.1242709, 0.05454769, 
    0.1285905, 0.001674097, 0.007128729, 0.2444813, 0.2072401,
  0.04576436, 0.08622721, 0.1405658, 0.09238292, 0.09139968, 0.09269958, 
    0.08536825, 0.08303849, 0.1132216, 0.1515377, 0.1364488, 0.1154808, 
    0.09798866, 0.08175193, 0.088871, 0.1274917, 0.1435151, 0.1147899, 
    0.1267092, 0.1167934, 0.05723505, 0.06189633, 0.00798047, 0.003218748, 
    0.003580964, 0.003225896, 0.001401164, 0.03444913, 0.07005591,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0002022144, 
    0.001085671, 0, 0, 0, 8.537545e-05, 0.0008900997, 0, 0, 0, 0, 0,
  0, 0.01193046, 0.02733343, 0.005602823, 0, 0, -6.10181e-08, -7.340041e-06, 
    -0.0004104085, 0, 0, -5.58411e-05, 4.034637e-05, -0.000390553, 
    0.0002024044, 0.005368578, 0.003179541, 0.007676322, 0.002059249, 
    -0.0005125684, 0.0188188, 0.02003611, 0.001084544, -9.222822e-06, 
    -4.384285e-06, 0, 0, 0, 0,
  -0.0001192807, 0.02251511, 0.07997135, 0.08355573, 0.06322459, 0.01314312, 
    0.0001173845, 0.003512274, 0.007942745, 0.01034614, 0.03879265, 
    0.03506137, 0.0589755, 0.03736556, 0.02630818, 0.03833663, 0.0386953, 
    0.04280279, 0.0123163, 0.01031469, 0.02830101, 0.04238012, 0.0413962, 
    0.06286543, 0.0285978, 0.0003275146, 0.01006297, 0.01525224, 0.005952614,
  0.1645053, 0.2264886, 0.205774, 0.2273051, 0.2182131, 0.1762931, 0.122844, 
    0.09669157, 0.07236572, 0.1186037, 0.152321, 0.15085, 0.1365617, 
    0.06112146, 0.06215897, 0.05641491, 0.08018178, 0.1188397, 0.1200853, 
    0.1540072, 0.1926749, 0.1190742, 0.1217361, 0.1059624, 0.1119532, 
    0.1714111, 0.1814353, 0.1348572, 0.1652354,
  0.1817043, 0.09179375, 0.06621864, 0.03653422, 0.03448311, 0.07114288, 
    0.0969202, 0.09673513, 0.1074552, 0.07808783, 0.0551259, 0.1034096, 
    0.04756135, 0.03263771, 0.02223683, 0.0621249, 0.139354, 0.1851934, 
    0.1681536, 0.2295282, 0.1805842, 0.1396522, 0.1476314, 0.1498301, 
    0.1568686, 0.129747, 0.167779, 0.1693172, 0.1651662,
  0.02275581, 0.005234607, 0.008616564, 0.0005688484, 0.01703613, 0.01402766, 
    5.446098e-05, 0.01139001, 0.0009215096, 0.0005957035, 0.02373274, 
    0.02750027, 0.0292972, 0.03173129, 0.1119532, 0.1202981, 0.1078217, 
    0.09265553, 0.149123, 0.0761488, 0.02772825, 0.007714777, 0.000989655, 
    0.005900359, 0.009275176, 0.03584344, 0.01002714, 0.04093973, 0.04565163,
  7.02321e-08, 2.300979e-08, 1.653245e-07, 0.01039181, 0.004376924, 
    -1.325045e-06, -8.631629e-06, 5.069107e-05, 4.77287e-06, 9.180119e-08, 
    7.183976e-09, 5.402052e-07, -8.135806e-07, 0.06845023, 0.05072253, 
    0.06087233, 0.03300926, 0.005318903, 0.001497198, 3.022975e-07, 
    -1.436005e-06, -4.713316e-09, 1.080421e-07, -2.74225e-06, 0.0002616316, 
    0.003650066, -5.41993e-06, 0.007083053, 5.505794e-07,
  -1.246098e-10, 3.833204e-06, 6.473137e-08, 0.0001410963, 0.002511085, 
    9.367199e-05, 0.05978252, 0.1852058, 0.01181731, 0.01282153, 0.0174589, 
    0.00353734, 0.058606, 0.1311584, 0.09573098, 0.0168493, 0.005066699, 
    1.944528e-05, 1.941669e-08, 3.030788e-07, 9.94726e-07, 3.391803e-07, 
    5.609724e-05, 0.0003117356, 2.379941e-07, 1.441455e-06, 6.180982e-07, 
    3.328e-07, 1.697256e-07,
  5.226139e-05, 0.1100189, 0.01654817, 5.399109e-05, 0.0004813017, 
    0.01291548, 0.01320614, 0.04272357, 0.1196296, 0.1682559, 0.03103727, 
    0.05454475, 0.05701808, 0.03948083, 0.05600176, 0.01720335, 0.0006327037, 
    3.330538e-05, -1.374029e-05, -1.307898e-05, -6.052176e-05, 0.0006798565, 
    0.01121181, 0.1155656, 0.04246761, 0.002287267, 0.002687539, 
    6.820676e-05, 1.132007e-06,
  0.1555193, 0.1823302, 0.07835669, 0.0722388, 0.007157112, 0.007963893, 
    0.04162534, 0.02369282, 0.07200629, 0.02172973, 0.007257737, 0.01707738, 
    0.06033165, 0.07470313, 0.05910714, 0.06191133, 0.02701267, 0.02853248, 
    0.07243815, 0.1217852, 0.376232, 0.2164788, 0.1651044, 0.04377132, 
    0.03492672, 0.06194463, 0.04862571, 0.2036047, 0.2627298,
  0.0007850883, 0.0002511156, 1.762918e-05, 0.01286082, 0.07998501, 
    0.08912935, 0.3310261, 0.09723846, 0.2338022, 0.01725561, 0.0876599, 
    0.07521617, 0.1012336, 0.09962668, 0.03643612, 0.02161727, 5.452192e-05, 
    2.148685e-05, 0.0003811784, 0.01296556, 0.03173834, 0.02404815, 
    0.0109355, 0.06584791, 0.03500398, 0.01599638, 0.001015953, 0.005007714, 
    0.0007171555,
  0.01578054, -1.239477e-05, -5.69157e-11, 4.962601e-07, 8.723947e-06, 
    -4.744645e-05, 0.05544255, 0.1401772, 0.1555108, 0.08919173, 0.06380375, 
    0.04070808, 0.1336581, 0.1591082, 0.03418789, 0.03786909, 0.003368657, 
    9.692819e-07, 0.01412017, 0.001476738, 0.03820832, 0.04152222, 
    0.07599527, 0.2449964, 0.05918955, 0.007106977, 2.218211e-06, 
    1.275878e-05, 0.002615014,
  0.01571626, 0.01015131, 0.001400978, 8.828699e-07, 0.02120818, 0.01560839, 
    0.1591747, 0.1402637, 0.1690502, 0.1185672, 0.2293268, 0.1627014, 
    0.1144735, 0.2248027, 0.2803172, 0.09986267, 0.07788914, 0.07005636, 
    0.0008572131, 0.000736838, 0.007962817, 0.01104957, 0.06024212, 
    0.0868325, 0.1345713, 0.127426, 0.04025348, 0.0159677, 0.01187554,
  0.1073393, 0.1262279, 0.03989468, 0.02796738, 0.04423309, 0.07912668, 
    0.07651765, 0.1005042, 0.1773944, 0.1904283, 0.1165621, 0.1409436, 
    0.140019, 0.03829246, 0.1315604, 0.1107275, 0.1172989, 0.1774834, 
    0.1338895, 0.07879727, 0.07848182, 0.06983528, 0.06860229, 0.1229636, 
    0.0915656, 0.09615048, 0.1086355, 0.1123387, 0.1176973,
  0.1739199, 0.1801758, 0.1096727, 0.05631904, 0.05280775, 0.06548497, 
    0.168581, 0.1325617, 0.1083173, 0.1163352, 0.2019072, 0.1661707, 
    0.1607711, 0.1553245, 0.09242773, 0.1834419, 0.1584803, 0.2178634, 
    0.2407258, 0.1555771, 0.2164939, 0.1788233, 0.1972586, 0.1553824, 
    0.2010034, 0.1512942, 0.07683966, 0.1525913, 0.198981,
  0.1595342, 0.1933075, 0.22514, 0.2175105, 0.1425915, 0.1400622, 0.1463612, 
    0.1817585, 0.1681875, 0.1820488, 0.1347992, 0.1243834, 0.1457981, 
    0.1128119, 0.1392784, 0.1893723, 0.1987545, 0.08907556, 0.1085221, 
    0.09072342, 0.1408096, 0.08402957, 0.1494073, 0.08032171, 0.1307053, 
    0.03734579, 0.0234737, 0.2388917, 0.2218011,
  0.08511925, 0.1396899, 0.1721932, 0.08164697, 0.08472835, 0.07882389, 
    0.1010331, 0.07335034, 0.1092125, 0.1283411, 0.1449439, 0.1313686, 
    0.1478763, 0.1554497, 0.1313755, 0.1429433, 0.1828458, 0.142915, 
    0.1476081, 0.1593494, 0.1586694, 0.158153, 0.08690117, 0.02827271, 
    0.05491906, 0.02916178, 0.05477811, 0.07806721, 0.08971449,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002669572, 0.001735117, 
    0.00767244, -5.696932e-05, 0, 0, 0.0001343824, 0.001594943, 
    -3.286719e-05, 0, 0, 0, 0,
  -0.0001179288, 0.02173078, 0.04634716, 0.04099308, -0.0007323122, 0, 
    0.0004013109, -4.767109e-05, -0.0006409824, -1.201691e-05, -5.590743e-06, 
    -6.46129e-05, 0.002795294, 0.02118024, 0.02649422, 0.01645788, 
    0.02764775, 0.05710061, 0.04556831, 0.03645648, 0.04524583, 0.03819874, 
    0.02374204, 0.002273263, 0.00056524, -2.956214e-07, -3.142202e-07, 
    -5.411417e-07, 0,
  0.03338126, 0.05566866, 0.1209566, 0.1727074, 0.144794, 0.07752271, 
    0.04397546, 0.05543052, 0.08507935, 0.07523137, 0.1761057, 0.1584976, 
    0.2001205, 0.1629352, 0.1282521, 0.1062832, 0.1134841, 0.1048522, 
    0.04140685, 0.08994116, 0.09650443, 0.07048228, 0.07688301, 0.1289372, 
    0.04831054, 0.05090216, 0.06794348, 0.03927256, 0.02597376,
  0.2346252, 0.2921457, 0.2263944, 0.2131284, 0.2157232, 0.2104379, 
    0.1488655, 0.1482308, 0.1922961, 0.222912, 0.2142202, 0.2052604, 
    0.2166479, 0.1452479, 0.1050297, 0.1048642, 0.1495114, 0.167273, 
    0.1619125, 0.1826124, 0.2451061, 0.185707, 0.1587611, 0.1340645, 
    0.1575027, 0.2357035, 0.2404679, 0.1725609, 0.2191972,
  0.1740382, 0.093173, 0.05509282, 0.03252842, 0.0279694, 0.08018596, 
    0.08905797, 0.1068638, 0.1050224, 0.08100728, 0.05053127, 0.09858663, 
    0.04620104, 0.04802914, 0.03031441, 0.07147181, 0.1363589, 0.1989849, 
    0.1858184, 0.2470371, 0.2137403, 0.1419504, 0.1551828, 0.2142229, 
    0.1394988, 0.1263884, 0.1641713, 0.1489934, 0.1509932,
  0.01910403, 0.01719989, 0.008697226, 0.005071485, 0.02860775, 0.02146441, 
    -0.0005347731, 0.007013911, 0.0003057194, 0.005374641, 0.03228286, 
    0.02702563, 0.03232365, 0.03140988, 0.1065854, 0.114808, 0.1042754, 
    0.08801154, 0.1264791, 0.06347395, 0.01703912, 0.005345069, 0.005860434, 
    0.005988254, 0.008646987, 0.0353117, 0.01109618, 0.04453664, 0.0400589,
  9.662423e-08, 3.305372e-10, 7.753076e-08, 0.01183782, 0.01169094, 
    -1.733045e-06, -8.49128e-05, -5.923198e-06, 6.549212e-06, 7.478529e-08, 
    1.123213e-09, 5.57445e-07, 0.002352448, 0.07361214, 0.04029969, 
    0.05472244, 0.01895184, 0.003586045, 0.000649206, -3.101102e-07, 
    -6.244471e-07, -1.042026e-10, 1.115365e-07, 6.668485e-06, 0.0001154629, 
    0.01205279, -2.336567e-06, 0.02333776, -1.829819e-06,
  4.235464e-09, 4.527546e-06, 1.80313e-08, 0.0001970784, 0.003173345, 
    0.000298811, 0.04750696, 0.1738976, 0.01320111, 0.0108817, 0.01791548, 
    0.02304715, 0.0500436, 0.1374998, 0.08447148, 0.01772844, 0.01210631, 
    3.480431e-06, 2.409678e-09, 6.950774e-08, 1.756846e-07, 3.790981e-07, 
    3.10505e-06, 0.0003377766, 8.020319e-07, 3.006694e-07, 8.996793e-06, 
    2.272744e-07, 3.234728e-08,
  2.96096e-05, 0.07731348, 0.01971786, 0.0009193891, 0.000619075, 0.01030685, 
    0.00974493, 0.02269846, 0.0806852, 0.1935713, 0.02991256, 0.04020471, 
    0.05472568, 0.03506087, 0.05224095, 0.0242374, 0.0009545371, 
    -4.304325e-05, 0.003975634, -1.925678e-06, -1.431227e-05, 0.0001546232, 
    0.01344244, 0.09954689, 0.05470967, 0.007312807, 0.00502927, 
    0.0002573498, 1.066569e-06,
  0.1162232, 0.1324656, 0.07679851, 0.0715036, 0.005180985, 0.005812009, 
    0.02838656, 0.01581476, 0.05664001, 0.01279815, 0.00495559, 0.009045701, 
    0.04535056, 0.07008892, 0.05038324, 0.05411275, 0.03221337, 0.04269277, 
    0.07690565, 0.1278822, 0.3633084, 0.209548, 0.1359814, 0.03614575, 
    0.03418312, 0.05650552, 0.03597518, 0.1826712, 0.2302484,
  0.006792814, 0.000271172, 1.139736e-05, 0.01456815, 0.07294799, 0.1122943, 
    0.2884001, 0.09457685, 0.2068172, 0.01094566, 0.09137746, 0.07109977, 
    0.07031718, 0.09094956, 0.02046583, 0.01286112, 5.422761e-05, 
    2.476264e-05, 5.918021e-05, 0.005296231, 0.03996802, 0.02529394, 
    0.00817547, 0.06561642, 0.02650842, 0.008037435, 0.01109719, 0.00162836, 
    0.004870983,
  0.02540069, -0.0001363322, -1.670344e-11, 4.503859e-08, 5.171216e-06, 
    -1.84133e-05, 0.04677039, 0.1437161, 0.1455373, 0.08146939, 0.06708555, 
    0.02740412, 0.1291228, 0.1567721, 0.01941643, 0.03221475, 0.0003521466, 
    4.365376e-08, 0.01913865, -2.945392e-06, 0.03318939, 0.03255824, 
    0.05064049, 0.2193355, 0.04145642, 0.005642243, 0.0004629182, 
    2.172391e-06, 0.02270796,
  0.01127467, 0.01109308, 0.00095683, 9.161288e-05, 0.03079413, 0.01869337, 
    0.1629572, 0.1296612, 0.1302525, 0.09407911, 0.1831195, 0.14681, 
    0.1184327, 0.2231193, 0.2700108, 0.07198237, 0.077434, 0.05395275, 
    0.0009802785, 0.0001387858, 0.01409384, 0.008591649, 0.05302362, 
    0.07488114, 0.1399936, 0.09591055, 0.03132792, 0.01305542, 0.01137441,
  0.09849297, 0.1201399, 0.0271133, 0.01902264, 0.0357177, 0.06568088, 
    0.06785567, 0.1053305, 0.1658581, 0.1850722, 0.1012282, 0.1320418, 
    0.1341694, 0.04112742, 0.1271079, 0.1035623, 0.1195156, 0.1626659, 
    0.1263912, 0.07259247, 0.05967524, 0.05961261, 0.05870201, 0.1221832, 
    0.08360342, 0.08936672, 0.09055742, 0.1127096, 0.1024565,
  0.1709738, 0.1838013, 0.1042168, 0.0568248, 0.03768675, 0.05601166, 
    0.1555513, 0.1268467, 0.09210697, 0.1065355, 0.175162, 0.1290283, 
    0.1588791, 0.1432667, 0.09638701, 0.187325, 0.147388, 0.2161224, 
    0.2403758, 0.1334838, 0.1730152, 0.1385104, 0.1622953, 0.1522637, 
    0.172431, 0.1371484, 0.06733333, 0.1500283, 0.191188,
  0.1530513, 0.1863547, 0.1989657, 0.1948533, 0.128117, 0.1318358, 0.148564, 
    0.1605373, 0.1272492, 0.1449673, 0.09837126, 0.119561, 0.1305481, 
    0.08349258, 0.1307642, 0.1810427, 0.1730722, 0.07413122, 0.0940029, 
    0.07488004, 0.1296564, 0.0835383, 0.1748084, 0.1112714, 0.1301923, 
    0.1810866, 0.1481244, 0.2275107, 0.201002,
  0.08949561, 0.152605, 0.1795678, 0.09380413, 0.08880523, 0.07828373, 
    0.1036757, 0.08623505, 0.1072463, 0.1068811, 0.1283849, 0.1684995, 
    0.175735, 0.1816669, 0.1515777, 0.156615, 0.1978838, 0.1326146, 
    0.1301407, 0.1496489, 0.166584, 0.1702285, 0.1590949, 0.0743205, 
    0.1391332, 0.06604078, 0.150175, 0.08514989, 0.08330145,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3.941166e-07, -0.0003712115, 
    0.01418658, 0.02544557, 0.02035151, 0.01726837, -0.0001420609, 0, 0, 
    0.001390764, 0.04647757, 0.03596747, 0.009844851, 0.01494798, 
    -2.050387e-05, 0,
  0.0156611, 0.02337574, 0.07340544, 0.09052461, -0.00324379, -0.0002343478, 
    0.02219593, -0.0001592686, -0.0005892768, -0.0009947657, 8.314777e-06, 
    0.0004306753, 0.01217733, 0.1502758, 0.1343995, 0.09489078, 0.104385, 
    0.141877, 0.123898, 0.1122058, 0.1480298, 0.1349147, 0.1241612, 
    0.04954048, 0.02816823, 0.01059037, 0.01140163, 0.00231311, 0.008611642,
  0.09539422, 0.1051007, 0.1763983, 0.2006592, 0.1880285, 0.129537, 
    0.06662578, 0.1068151, 0.1047037, 0.1287712, 0.2517045, 0.2024336, 
    0.22941, 0.2072223, 0.1579213, 0.151044, 0.2249725, 0.2248606, 0.1658789, 
    0.1883319, 0.2114842, 0.2247863, 0.1630944, 0.248529, 0.161454, 
    0.1362341, 0.1309132, 0.09960474, 0.1088522,
  0.2831137, 0.3135616, 0.2158856, 0.2057482, 0.2193276, 0.2207969, 
    0.1810859, 0.1555229, 0.2245135, 0.2422031, 0.2302528, 0.203234, 
    0.1976707, 0.1275977, 0.1286888, 0.1772314, 0.1677527, 0.2397989, 
    0.1977318, 0.2103699, 0.2507735, 0.1750229, 0.1989475, 0.1608209, 
    0.1773982, 0.248013, 0.2657574, 0.1909108, 0.2469558,
  0.1464279, 0.09110085, 0.04025664, 0.02754215, 0.03131691, 0.07363974, 
    0.08590476, 0.1074397, 0.09427737, 0.08769657, 0.05664564, 0.08586655, 
    0.03201624, 0.03555711, 0.02855297, 0.07677154, 0.1298693, 0.2009429, 
    0.198632, 0.2408953, 0.2142124, 0.1493025, 0.1691535, 0.2444673, 
    0.1112275, 0.1158779, 0.1424385, 0.1359613, 0.1322048,
  0.01779165, 0.03457698, 0.008546527, 0.01353902, 0.04313606, 0.0338207, 
    0.0001328465, -0.0001603671, -4.779366e-06, 0.002104803, 0.02619182, 
    0.01223103, 0.03083133, 0.02612673, 0.08387007, 0.1207667, 0.09936982, 
    0.075106, 0.1217276, 0.04867483, 0.01739394, 0.003712794, 0.0020375, 
    0.0002830336, 0.009145525, 0.04126222, 0.01133222, 0.0434459, 0.03384416,
  1.134966e-08, -2.323593e-10, -3.588451e-08, 0.01550057, 0.01432872, 
    -3.807473e-07, 0.0004470855, 6.715578e-07, 2.698039e-06, 5.361228e-08, 
    3.329858e-10, 3.318603e-07, 0.001017625, 0.07545281, 0.04376503, 
    0.05180946, 0.01049658, 0.0009878079, 0.0001407489, 6.125089e-07, 
    -1.572322e-07, 2.055221e-08, 9.616499e-08, 2.855907e-05, 0.0004790107, 
    0.005795069, -1.491823e-05, 0.0265884, -6.444746e-05,
  -3.099482e-09, 6.93444e-06, 7.881939e-08, 0.0001319907, 0.004198902, 
    0.0007110276, 0.03126099, 0.1681529, 0.01047318, 0.009057157, 0.0119938, 
    0.03077757, 0.05190327, 0.1412627, 0.08981093, 0.02205181, 0.01788092, 
    8.133653e-06, 8.241869e-07, 5.162634e-09, 1.080057e-07, 2.807219e-07, 
    1.472737e-06, 0.0003902144, 2.674016e-07, 2.292427e-07, 0.0001023493, 
    1.265591e-07, 6.463038e-08,
  4.994956e-05, 0.06308462, 0.03443096, 0.003759445, 0.0008939803, 
    0.009389744, 0.009391858, 0.01749966, 0.0642432, 0.2234046, 0.03009348, 
    0.03186534, 0.04446507, 0.03713478, 0.06154164, 0.02238816, 0.001958866, 
    -7.807293e-05, 0.005913169, 3.385043e-06, -0.0001305537, -6.358699e-06, 
    0.02476616, 0.08708637, 0.07200562, 0.01297149, 0.01569854, 0.001130588, 
    2.63609e-06,
  0.1021985, 0.11297, 0.09244104, 0.08670873, 0.01831258, 0.01617013, 
    0.0208295, 0.01205743, 0.05781157, 0.009270853, 0.004491354, 0.008517154, 
    0.0406174, 0.06182607, 0.04524425, 0.05744708, 0.04293369, 0.05482927, 
    0.07662163, 0.1491183, 0.3505038, 0.1986136, 0.1082589, 0.03150157, 
    0.03890739, 0.0583196, 0.03365088, 0.1807833, 0.2152915,
  0.04155526, 0.0005196459, 5.236891e-05, 0.03343761, 0.08863684, 0.1094257, 
    0.2195934, 0.1110593, 0.1917726, 0.008150959, 0.1040647, 0.07593278, 
    0.06370752, 0.08292162, 0.01153257, 0.00994257, 5.381876e-05, 
    1.740579e-05, 0.0001237881, 0.01297965, 0.03014441, 0.02646284, 
    0.006808661, 0.0623408, 0.01831731, 0.006125494, 0.0133504, 0.001615996, 
    0.02934809,
  0.04944043, -8.732302e-05, 0, 2.247121e-08, -1.780679e-05, -1.075677e-05, 
    0.02979377, 0.1587985, 0.1487894, 0.08209901, 0.06273688, 0.0190121, 
    0.1227016, 0.1335928, 0.01517939, 0.02425946, 3.350906e-05, 
    -2.497238e-07, 0.03329553, 1.314391e-05, 0.03619289, 0.02708407, 
    0.03751464, 0.1730387, 0.03156087, 0.004242368, 1.989018e-06, 
    6.957508e-07, 0.04620667,
  0.01328625, 0.01150344, 0.001036761, 0.000199352, 0.04185954, 0.01401305, 
    0.1495656, 0.1205432, 0.1083018, 0.08002761, 0.1441325, 0.1373135, 
    0.1022082, 0.2449357, 0.2463956, 0.05504481, 0.05874785, 0.05084689, 
    0.001604883, 0.0001391413, 0.0388503, 0.006868945, 0.0522282, 0.07990444, 
    0.118488, 0.06514147, 0.01944173, 0.00926451, 0.007352524,
  0.07372318, 0.1196185, 0.02606841, 0.01668677, 0.03440401, 0.06217898, 
    0.05666326, 0.0974813, 0.1557911, 0.1794048, 0.09079005, 0.1238562, 
    0.1259396, 0.03281388, 0.1236233, 0.1032974, 0.09935542, 0.1640705, 
    0.1353206, 0.07198527, 0.05443426, 0.05580403, 0.05151883, 0.1251716, 
    0.0753848, 0.08445567, 0.0931818, 0.116113, 0.1073109,
  0.1501484, 0.1691441, 0.09992975, 0.04718517, 0.02229555, 0.06195078, 
    0.1374175, 0.1363268, 0.08131596, 0.09960042, 0.1456239, 0.1181621, 
    0.1433485, 0.1305645, 0.1042022, 0.2045205, 0.1456622, 0.2099264, 
    0.235941, 0.1263435, 0.1313189, 0.1141837, 0.156641, 0.153176, 0.1498571, 
    0.1260229, 0.07091677, 0.1366854, 0.1743272,
  0.1507425, 0.1891059, 0.1874952, 0.1830042, 0.1265785, 0.1153948, 
    0.1463736, 0.1448595, 0.1187504, 0.1337119, 0.07096037, 0.1196163, 
    0.115843, 0.06142604, 0.1484675, 0.170394, 0.1410307, 0.06519519, 
    0.08280353, 0.06871968, 0.1364055, 0.09443724, 0.1860216, 0.1230445, 
    0.1233192, 0.2049086, 0.2294786, 0.2100421, 0.186088,
  0.09806636, 0.1701443, 0.1927306, 0.1066729, 0.08253603, 0.06050159, 
    0.09594318, 0.08300759, 0.07626852, 0.09874493, 0.1248776, 0.1827474, 
    0.1955952, 0.2081534, 0.1826069, 0.1665685, 0.2114207, 0.1370541, 
    0.1196857, 0.1478021, 0.1730428, 0.1680503, 0.1595604, 0.08046885, 
    0.2105339, 0.1807156, 0.2194206, 0.07803807, 0.08205395,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.009520083, 0.08706271, 0.1285906, 
    0.1518776, 0.08180089, 0.03587512, 0.0009179618, -0.0004178851, 
    1.146585e-05, 0.009165776, 0.07767239, 0.07668839, 0.05206295, 
    0.06609548, 0.0006789163, 0,
  0.05798323, 0.05288481, 0.1858795, 0.1994144, 0.01537472, -0.001079193, 
    0.03475579, 0.0002165323, 0.0007984407, 0.004169872, -7.600054e-05, 
    0.0009799692, 0.07283808, 0.1741707, 0.2250435, 0.1784264, 0.1798474, 
    0.2450132, 0.2323058, 0.2400717, 0.2829297, 0.2683742, 0.2596768, 
    0.1735136, 0.1172889, 0.05371371, 0.06751142, 0.06217546, 0.06189189,
  0.1187538, 0.1900075, 0.2309496, 0.2524472, 0.2067486, 0.158164, 
    0.08682402, 0.1391542, 0.1583926, 0.1651058, 0.2929681, 0.2539898, 
    0.2591507, 0.2302748, 0.1910803, 0.179416, 0.2593294, 0.2425464, 
    0.1948674, 0.1824982, 0.2166839, 0.2632354, 0.197087, 0.2784242, 
    0.2268998, 0.1947626, 0.181509, 0.167365, 0.1439331,
  0.3220257, 0.3198377, 0.2328993, 0.2104136, 0.2108083, 0.2218063, 
    0.1869559, 0.1611107, 0.2817318, 0.2619618, 0.228882, 0.200226, 
    0.1798741, 0.120513, 0.1220155, 0.1842466, 0.17389, 0.2320132, 0.1897704, 
    0.2174061, 0.2623689, 0.2100808, 0.187389, 0.1981349, 0.1652659, 
    0.2525517, 0.2573284, 0.1918657, 0.2481279,
  0.1535928, 0.08529269, 0.04248044, 0.0220214, 0.03456591, 0.06484491, 
    0.08687458, 0.1102433, 0.09928075, 0.07660796, 0.06292773, 0.08830144, 
    0.02517111, 0.02688951, 0.02374325, 0.06239506, 0.1256163, 0.1992567, 
    0.2161587, 0.226142, 0.2194062, 0.1456559, 0.1534175, 0.2529172, 
    0.08176111, 0.1123423, 0.1247943, 0.1501941, 0.1227347,
  0.01479371, 0.04623178, 0.01814783, 0.02169604, 0.04110053, 0.03819378, 
    0.005308679, 0.0005026353, -3.603651e-06, 0.0004521891, 0.0209089, 
    0.009295165, 0.03689493, 0.01718904, 0.07288744, 0.1158573, 0.09021469, 
    0.05777419, 0.1148759, 0.04241504, 0.01408615, 0.006980597, 0.003027046, 
    0.0004090369, 0.008047614, 0.0564857, 0.0155014, 0.04270118, 0.03085971,
  -7.767682e-08, 0, -1.434496e-07, 0.02085876, 0.03072993, 2.595426e-05, 
    0.005078903, 2.906357e-06, 1.548733e-06, 2.328524e-08, 2.827668e-12, 
    2.98187e-07, 0.0009294037, 0.07770787, 0.04289243, 0.04066723, 
    0.01130925, 0.0004653028, 0.001685314, -3.106139e-07, -9.215744e-07, 
    2.704881e-08, 8.425188e-08, 4.25076e-07, 0.0002724527, 7.653268e-05, 
    -0.0001505331, 0.02751954, 0.003395675,
  4.431492e-08, 3.066201e-06, 3.089167e-08, 9.572936e-05, 0.008203337, 
    0.001509243, 0.01989772, 0.1395555, 0.01023378, 0.01124768, 0.004735229, 
    0.02856479, 0.06083817, 0.1356027, 0.07879185, 0.02710305, 0.01409405, 
    2.258412e-05, 9.948356e-06, 5.514922e-09, -2.444682e-11, 4.891424e-08, 
    7.155654e-07, 0.0006064428, -0.0001260972, 1.377643e-07, 0.000219491, 
    8.586958e-05, 3.331329e-08,
  0.0008094869, 0.05572743, 0.03324717, 0.002406781, 0.001583518, 
    0.009031262, 0.008300311, 0.01238883, 0.07584622, 0.2459858, 0.02748344, 
    0.03255556, 0.0375827, 0.03186635, 0.06191542, 0.02134234, 0.005101097, 
    -7.413424e-05, 0.001619062, 0.0002657678, -0.0001698557, 3.407662e-05, 
    0.02035749, 0.08856207, 0.08748503, 0.02830292, 0.02387739, 0.001763715, 
    3.361144e-06,
  0.09585937, 0.115607, 0.0960166, 0.1165777, 0.01651002, 0.01375109, 
    0.01698863, 0.009371373, 0.03893064, 0.008225181, 0.003573277, 
    0.006292832, 0.04212381, 0.04695204, 0.0423332, 0.06761631, 0.05334155, 
    0.07132103, 0.07759474, 0.190811, 0.3416647, 0.1621696, 0.0814352, 
    0.03389588, 0.04241681, 0.05495256, 0.05509365, 0.2070647, 0.2181385,
  0.02400291, 0.00270002, 1.082878e-05, 0.01645449, 0.07963821, 0.07819258, 
    0.2126702, 0.127557, 0.2095363, 0.006206739, 0.109524, 0.07807101, 
    0.06884397, 0.07429802, 0.009877597, 0.007040187, 4.615041e-05, 
    1.022492e-05, 0.0001629244, 0.01206244, 0.02881377, 0.02539539, 
    0.005336607, 0.07559239, 0.01593995, 0.008953372, 0.01679998, 
    0.001274102, 0.02354595,
  0.03731185, -3.738122e-05, 8.717324e-11, 1.687816e-08, -1.356298e-05, 
    -6.696035e-05, 0.03215201, 0.1664621, 0.1537071, 0.09090045, 0.0621702, 
    0.01833209, 0.1192936, 0.1138704, 0.004830107, 0.02554688, 8.624726e-06, 
    -2.308926e-07, 0.02095703, 0.0001943638, 0.04175515, 0.02192105, 
    0.03284721, 0.1452948, 0.02120166, 0.00264887, 5.911544e-07, 
    4.105501e-07, 0.03623243,
  0.01731839, 0.005466778, 0.0007394753, 0.0001141749, 0.05633467, 
    0.01531223, 0.1557083, 0.09975114, 0.09798387, 0.07537831, 0.1166369, 
    0.1151647, 0.0971009, 0.239498, 0.219294, 0.05736227, 0.04886999, 
    0.04755687, 0.001144926, 0.0001615521, 0.09930295, 0.006743762, 
    0.0700999, 0.08936085, 0.1166086, 0.0592044, 0.01493912, 0.008255473, 
    0.004223301,
  0.05451003, 0.113989, 0.03100467, 0.01889274, 0.03085096, 0.07235222, 
    0.06175167, 0.08678041, 0.1460587, 0.1841272, 0.091287, 0.09730693, 
    0.1228716, 0.03451955, 0.1032385, 0.1075609, 0.105716, 0.1755262, 
    0.1122636, 0.0798449, 0.05297449, 0.05389771, 0.05279854, 0.1110781, 
    0.07503273, 0.07614198, 0.0895238, 0.1266935, 0.1422945,
  0.1660514, 0.1634348, 0.1049319, 0.04629345, 0.01445839, 0.06516763, 
    0.1320421, 0.1495422, 0.0799144, 0.09422275, 0.1110665, 0.1067513, 
    0.1473121, 0.1319139, 0.1039375, 0.1942685, 0.1501621, 0.2262648, 
    0.2416269, 0.1166961, 0.1100116, 0.1059669, 0.1358235, 0.1486675, 
    0.1553315, 0.1233494, 0.06140836, 0.157455, 0.1608086,
  0.1863108, 0.2429154, 0.1876083, 0.1660712, 0.1269835, 0.1056195, 0.133244, 
    0.1240959, 0.1196172, 0.1192399, 0.0678812, 0.1386436, 0.09574739, 
    0.0510725, 0.1304845, 0.1646962, 0.1124628, 0.06344749, 0.06166777, 
    0.06662694, 0.1388616, 0.1086459, 0.1906105, 0.1469244, 0.1353017, 
    0.2089496, 0.2366276, 0.2030035, 0.212554,
  0.1123776, 0.1827, 0.2008881, 0.1229787, 0.07433837, 0.05571627, 0.0895023, 
    0.06802315, 0.08449347, 0.1091334, 0.1523352, 0.1908906, 0.2173769, 
    0.2554275, 0.1930127, 0.1764034, 0.2341121, 0.146821, 0.1264497, 
    0.1591543, 0.1883392, 0.1546484, 0.1649805, 0.09182408, 0.2108996, 
    0.2071948, 0.2203448, 0.06959799, 0.08862444,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.013948e-06, 0.1068444, 0.1629395, 
    0.166644, 0.1861793, 0.1271242, 0.1166222, 0.01999651, 0.01088428, 
    -0.001337272, 0.03907703, 0.1232335, 0.1558121, 0.1397012, 0.1469933, 
    0.04063392, 0.0001391863,
  0.1528188, 0.1681877, 0.2628091, 0.2501452, 0.07262664, 0.0006699112, 
    0.09170003, 0.01467463, 0.01565121, 0.02444059, 0.002336408, 0.006909316, 
    0.1414771, 0.2464444, 0.3128556, 0.2346406, 0.2053375, 0.3027171, 
    0.2662164, 0.2627576, 0.2784426, 0.2588796, 0.2463272, 0.2033518, 
    0.1382275, 0.153741, 0.1557851, 0.1389049, 0.1558713,
  0.1395257, 0.2208214, 0.2597421, 0.2792874, 0.2364795, 0.1844848, 
    0.0866365, 0.1714182, 0.1748263, 0.1590636, 0.3261386, 0.2611206, 
    0.2495642, 0.2644551, 0.1967687, 0.1832749, 0.2595993, 0.2376374, 
    0.1977563, 0.1786175, 0.2218773, 0.2668611, 0.2135412, 0.2919389, 
    0.2156923, 0.22455, 0.2016625, 0.1660945, 0.1313449,
  0.3161179, 0.2998019, 0.2190959, 0.2042107, 0.1999887, 0.2155478, 
    0.1884756, 0.1707858, 0.2795225, 0.2759219, 0.2248722, 0.162638, 
    0.1680878, 0.1127965, 0.1329341, 0.159372, 0.148299, 0.2201856, 
    0.2099798, 0.2095518, 0.2457086, 0.1900512, 0.1884177, 0.1891705, 
    0.156351, 0.2492606, 0.2648751, 0.1965094, 0.236939,
  0.1445691, 0.08036044, 0.04670871, 0.02083924, 0.03992865, 0.06210734, 
    0.09101445, 0.1205214, 0.09508526, 0.0668318, 0.06383561, 0.08670619, 
    0.03104971, 0.02695347, 0.02371768, 0.06487962, 0.1210664, 0.1794406, 
    0.2043119, 0.2124737, 0.2020587, 0.138168, 0.1562747, 0.2773773, 
    0.06358722, 0.1011912, 0.1305782, 0.1428704, 0.115521,
  0.014976, 0.04352319, 0.02964386, 0.01245551, 0.04679161, 0.02859021, 
    0.01188437, 0.002016725, 4.705242e-05, 0.001912191, 0.00821584, 
    0.009090846, 0.03812206, 0.01355778, 0.06839734, 0.0801678, 0.1090981, 
    0.04796908, 0.1254788, 0.04229897, 0.01455205, 0.008646863, 0.00556477, 
    0.0005251181, 0.006451999, 0.06890513, 0.01882691, 0.04387214, 0.03342221,
  -1.060456e-05, -3.548031e-11, -1.054264e-07, 0.03025568, 0.03667803, 
    0.0004275264, 0.009123707, 0.0001875583, 9.832816e-07, 1.33721e-09, 
    7.523815e-11, 4.4419e-07, 0.002897965, 0.07503477, 0.05199941, 
    0.02971916, 0.01236952, 0.002949869, 0.0001630496, -3.078012e-06, 
    -5.144393e-06, 3.263696e-08, 7.263736e-08, 1.367117e-07, 0.0002604966, 
    5.987128e-05, 0.0002542741, 0.02737561, 0.007335752,
  4.980427e-08, 2.012755e-06, 2.506554e-06, 0.0001144621, 0.0119248, 
    0.00639388, 0.02533528, 0.1416713, 0.009437571, 0.01477543, 0.003109998, 
    0.01473904, 0.07162587, 0.1374834, 0.08873361, 0.03855376, 0.0212811, 
    0.0007726342, 6.448358e-05, 5.043648e-08, 2.039075e-08, 1.569277e-07, 
    8.328381e-06, 0.001024492, -9.37502e-06, 6.212789e-09, 6.04825e-06, 
    3.609993e-05, 6.504977e-08,
  0.002467229, 0.063736, 0.04093474, 0.01100805, 0.001412438, 0.008699858, 
    0.009187643, 0.01299782, 0.09725949, 0.258823, 0.02824119, 0.03925904, 
    0.04227958, 0.03640994, 0.06175733, 0.01388687, 0.01577562, 0.0002374068, 
    -9.85276e-05, 0.006389168, 0.001884364, 0.0006809126, 0.01957816, 
    0.06844825, 0.09363358, 0.05630206, 0.03302136, 0.02239279, 0.007470751,
  0.08936877, 0.1194403, 0.0937999, 0.1847885, 0.01669819, 0.02748491, 
    0.02159726, 0.009200823, 0.03723316, 0.007235488, 0.00381839, 
    0.006315432, 0.04230694, 0.05308032, 0.04649194, 0.07837054, 0.05476785, 
    0.08315724, 0.07904425, 0.2112674, 0.3416339, 0.1408001, 0.08896906, 
    0.04236971, 0.04665134, 0.05138551, 0.07750464, 0.2026826, 0.2184302,
  0.003769117, 0.0007492015, 1.642172e-05, 0.0008395029, 0.05456841, 
    0.07942858, 0.2452807, 0.1505471, 0.2705268, 0.01351169, 0.1463336, 
    0.08336806, 0.07830256, 0.07416549, 0.009090014, 0.003258898, 
    8.196803e-05, 6.800239e-05, 0.006191563, 0.021227, 0.04591284, 
    0.02665705, 0.004746667, 0.08000071, 0.01118109, 0.0116759, 0.0114492, 
    0.0004308755, 0.00350492,
  0.007098417, -5.446044e-06, -1.235664e-10, 2.164348e-08, 0.0006263481, 
    -2.476014e-05, 0.05068787, 0.1719602, 0.16955, 0.1008622, 0.06579043, 
    0.02585823, 0.1253293, 0.1100437, 0.001298093, 0.02457581, 7.770914e-06, 
    3.154922e-06, 0.01526032, 6.125339e-05, 0.0491244, 0.02430024, 
    0.04079234, 0.1340895, 0.01620782, 0.002421197, 1.202447e-05, 
    2.046416e-07, 0.01146556,
  0.01545726, 0.0004959857, 0.001057272, 0.0004922378, 0.05091158, 0.0124108, 
    0.1665623, 0.06044277, 0.0786115, 0.08732642, 0.107665, 0.1072484, 
    0.1000423, 0.2299334, 0.1918026, 0.05916933, 0.02404815, 0.03374572, 
    0.001738359, 0.0002520633, 0.1263911, 0.01676591, 0.07578176, 0.1047623, 
    0.117791, 0.05226018, 0.0179378, 0.007285682, 0.003549634,
  0.06690719, 0.09812964, 0.03152123, 0.02011637, 0.02905467, 0.07244266, 
    0.07632619, 0.09435848, 0.1389789, 0.1968494, 0.08601964, 0.07603276, 
    0.12228, 0.03182013, 0.1123998, 0.1177112, 0.1164528, 0.173734, 
    0.1256612, 0.07681644, 0.05167233, 0.04810509, 0.04470148, 0.1111232, 
    0.09643088, 0.06573278, 0.0968568, 0.1038096, 0.1234273,
  0.1468371, 0.157672, 0.1012395, 0.06219723, 0.01412172, 0.06117957, 
    0.1048395, 0.1467996, 0.07665853, 0.1046663, 0.09849457, 0.1105454, 
    0.1531042, 0.1171014, 0.1065497, 0.2237408, 0.2154669, 0.2356362, 
    0.2884741, 0.1262434, 0.08199882, 0.1215159, 0.1493483, 0.1596413, 
    0.1797443, 0.1299198, 0.07591964, 0.1652995, 0.1740957,
  0.1966522, 0.2455572, 0.1984539, 0.1617409, 0.1256931, 0.09677042, 
    0.1251909, 0.1687953, 0.1051816, 0.1125773, 0.08497041, 0.1294612, 
    0.0889075, 0.04499911, 0.1028884, 0.1308071, 0.07897975, 0.06073765, 
    0.04610156, 0.0620732, 0.1477792, 0.1065049, 0.1877968, 0.1635385, 
    0.1423163, 0.2119516, 0.2301002, 0.1936977, 0.2044392,
  0.1037742, 0.1913503, 0.2268111, 0.1388223, 0.08556052, 0.06072962, 
    0.09947414, 0.05714322, 0.1217627, 0.1390888, 0.1821253, 0.2243327, 
    0.2736718, 0.3226141, 0.249598, 0.2300909, 0.269553, 0.2165766, 
    0.1417697, 0.1646869, 0.252881, 0.1998618, 0.19225, 0.1208914, 0.2280344, 
    0.2127062, 0.2084283, 0.06965523, 0.07388927,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  -9.909024e-05, -4.007819e-06, 0, 0, 0, 0, 0, 0, -2.705829e-08, 0, 
    -1.386252e-06, 8.666985e-05, 0.0007098507, 0.1686279, 0.1593839, 
    0.1704404, 0.1990605, 0.2059925, 0.152998, 0.0383988, 0.02520563, 
    0.006869948, 0.08071948, 0.1801987, 0.1843408, 0.1803378, 0.207394, 
    0.1147712, 0.004155538,
  0.2537373, 0.2300283, 0.2905399, 0.3014347, 0.1157634, 0.01474127, 
    0.1189619, 0.04347223, 0.05227064, 0.05972124, 0.03741278, 0.04046839, 
    0.2368463, 0.2769854, 0.3282404, 0.2768796, 0.1984186, 0.3152755, 
    0.2609846, 0.2798899, 0.296847, 0.249614, 0.2167746, 0.1988209, 
    0.1640422, 0.1587048, 0.1725209, 0.1724094, 0.2405556,
  0.1446626, 0.2280777, 0.2587916, 0.2798682, 0.2343237, 0.2116055, 0.104983, 
    0.2033919, 0.2266887, 0.2015898, 0.3041355, 0.2674176, 0.2445783, 
    0.2544623, 0.1813517, 0.1845116, 0.2380995, 0.2129932, 0.188346, 
    0.1710109, 0.2106693, 0.2548459, 0.2030472, 0.2669756, 0.1837966, 
    0.2177877, 0.1956244, 0.1662369, 0.131467,
  0.3028455, 0.287237, 0.2184381, 0.2113396, 0.1978574, 0.2088405, 0.2027304, 
    0.1844512, 0.2675533, 0.2445175, 0.2034417, 0.1463736, 0.1556832, 
    0.124366, 0.1357197, 0.1678154, 0.1495564, 0.2068592, 0.2031434, 
    0.2037938, 0.2348421, 0.1752405, 0.1738005, 0.1702948, 0.156094, 
    0.2264541, 0.2691522, 0.2104186, 0.2341984,
  0.1511814, 0.08200896, 0.04384218, 0.03255622, 0.04808161, 0.06033437, 
    0.08433305, 0.1168713, 0.09593049, 0.0777539, 0.07117074, 0.08055351, 
    0.04077894, 0.03008064, 0.02041766, 0.06120038, 0.114146, 0.165308, 
    0.1903534, 0.1951382, 0.1855095, 0.1359872, 0.161925, 0.2904194, 
    0.05131629, 0.08630589, 0.1293427, 0.1425311, 0.1146636,
  0.01691214, 0.02807944, 0.04357348, 0.009158303, 0.06284458, 0.02510474, 
    0.009387344, 0.004069963, 0.0005176132, 0.004095911, 0.0005133469, 
    0.02106556, 0.05347671, 0.02178452, 0.06220568, 0.05824275, 0.1151489, 
    0.0373575, 0.1224266, 0.04246034, 0.01621493, 0.01262915, 0.007246604, 
    0.003499792, 0.007039316, 0.08299684, 0.02091439, 0.03983277, 0.03142314,
  -8.845265e-07, -1.850667e-09, -1.959602e-07, 0.04207591, 0.04239972, 
    0.0006036765, 0.0186947, -8.253327e-06, 2.386557e-06, 1.310067e-07, 
    1.396961e-08, 3.95104e-05, 0.01366943, 0.07382502, 0.05547763, 
    0.02061459, 0.008302665, 0.005630273, -1.546232e-05, 3.786664e-05, 
    -2.825988e-05, 4.239236e-08, 1.189404e-07, 2.752799e-06, 0.0002735642, 
    2.563297e-05, 0.001967506, 0.02600423, 0.002025604,
  1.102024e-07, 8.320704e-06, 3.669932e-05, 0.001051475, 0.02450482, 
    0.00159638, 0.0380843, 0.1497412, 0.01908015, 0.01216564, 0.00557228, 
    0.005216119, 0.08087704, 0.1418335, 0.1130489, 0.04925305, 0.03436216, 
    0.001069852, 0.0001073313, 1.386418e-07, 1.143072e-07, 5.579197e-07, 
    1.354237e-05, 0.0007996936, -1.046175e-06, 6.504594e-08, -7.966889e-06, 
    0.000104945, 2.231938e-07,
  0.004121163, 0.07857019, 0.05981909, 0.01443295, 0.001063261, 0.01030112, 
    0.0207161, 0.02065718, 0.1395548, 0.300394, 0.04357944, 0.06147032, 
    0.05512115, 0.04951937, 0.06691657, 0.01451676, 0.02402303, 0.0002997668, 
    0.001608598, 0.003832927, 0.009771682, 0.001383316, 0.02320135, 
    0.06046242, 0.1070119, 0.06781942, 0.03919129, 0.002653909, 0.01546235,
  0.1094376, 0.1399216, 0.1008008, 0.2405948, 0.01506144, 0.02562218, 
    0.03946196, 0.01964446, 0.05059529, 0.0107174, 0.006836038, 0.01445773, 
    0.05594269, 0.06650022, 0.06538764, 0.0891123, 0.05662528, 0.1047086, 
    0.102989, 0.2400496, 0.3830135, 0.1430773, 0.1072032, 0.05895781, 
    0.05853036, 0.06711145, 0.09390426, 0.2329896, 0.251497,
  0.007196733, 0.002968982, 0.0001281301, 4.828003e-05, 0.03666236, 
    0.08954108, 0.29967, 0.20739, 0.342098, 0.03872387, 0.1733337, 0.1071156, 
    0.113991, 0.07875921, 0.008915653, 0.00283492, 9.359091e-05, 
    9.409993e-05, 0.005611307, 0.03553917, 0.07440808, 0.03126026, 
    0.006172813, 0.08095044, 0.01705118, 0.01659158, 0.004557594, 
    0.0002654458, 0.003664799,
  0.0002545509, 2.722188e-06, -1.1409e-10, 5.5703e-08, 0.0007060869, 
    0.00081178, 0.06904373, 0.1966839, 0.2065276, 0.1139326, 0.07537364, 
    0.04457065, 0.154673, 0.1054377, 0.002178957, 0.02817533, 1.003646e-05, 
    1.574755e-05, 0.008159442, 0.00125265, 0.06192458, 0.03595445, 
    0.06706705, 0.1458095, 0.01653069, 0.002448127, 4.189201e-05, 
    1.222934e-06, 0.001180082,
  0.01806085, 1.93351e-05, 0.00861381, 0.002177649, 0.02180539, 0.01221736, 
    0.1637304, 0.03100587, 0.06353753, 0.08784902, 0.111877, 0.1148673, 
    0.1144131, 0.2445416, 0.1991721, 0.06129239, 0.01860499, 0.02986916, 
    0.001590704, 0.0003305625, 0.06610179, 0.02220721, 0.08413802, 0.1393433, 
    0.1347347, 0.07017342, 0.02403335, 0.007863327, 0.002879217,
  0.05269414, 0.09241609, 0.03711206, 0.0243915, 0.03237848, 0.07822868, 
    0.09660758, 0.1059244, 0.1290255, 0.1918779, 0.07703273, 0.07599442, 
    0.1196897, 0.03954263, 0.1084465, 0.122226, 0.1077683, 0.2046863, 
    0.1228403, 0.07908133, 0.05267014, 0.05513455, 0.05544959, 0.1330373, 
    0.09483684, 0.06296784, 0.08673699, 0.09765054, 0.1145281,
  0.1427852, 0.1770824, 0.1106266, 0.05461767, 0.01243079, 0.05796542, 
    0.1177026, 0.156936, 0.07452089, 0.1044039, 0.08740771, 0.1160275, 
    0.1753378, 0.125065, 0.125226, 0.1988801, 0.1967895, 0.2391185, 
    0.3616118, 0.1430224, 0.06414207, 0.1072737, 0.1768497, 0.1975249, 
    0.1590132, 0.1635474, 0.06020244, 0.2171066, 0.1832819,
  0.2107765, 0.2305439, 0.1721306, 0.1459348, 0.1234488, 0.09644222, 
    0.1144057, 0.1640679, 0.1122904, 0.1252523, 0.1089463, 0.1400905, 
    0.09068397, 0.03240498, 0.08359411, 0.1302776, 0.10068, 0.06263592, 
    0.04781878, 0.06651425, 0.1464759, 0.1010061, 0.2063171, 0.1890978, 
    0.1966012, 0.2226998, 0.2202815, 0.1666978, 0.1987458,
  0.09884105, 0.1624019, 0.2085267, 0.1467086, 0.1227376, 0.08510598, 
    0.104506, 0.075966, 0.08512098, 0.1270983, 0.1658654, 0.2129314, 
    0.2457515, 0.2916521, 0.2405135, 0.2240002, 0.2587991, 0.1969058, 
    0.17018, 0.174437, 0.2150849, 0.1870762, 0.2359076, 0.136433, 0.2308304, 
    0.2059351, 0.1773351, 0.07188955, 0.06347828,
  1.341797e-05, 3.779102e-06, -5.859766e-06, -1.549863e-05, -2.51375e-05, 
    -3.477637e-05, -4.441524e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -4.156769e-05, -3.192882e-05, -2.228995e-05, -1.265108e-05, 
    -3.012216e-06, 6.626652e-06, 1.626552e-05, 2.112906e-05,
  -0.002178703, -0.0002003084, 0.002371695, -5.783856e-05, 0, -4.223028e-05, 
    0.0001901192, -3.346406e-05, 1.919127e-05, 0.0003336427, 0.001293382, 
    0.001539013, 0.001804817, 0.1781393, 0.1770859, 0.1856423, 0.1839998, 
    0.2211672, 0.1999802, 0.06899141, 0.05035758, 0.02858903, 0.1300953, 
    0.1778684, 0.184363, 0.1963458, 0.2567317, 0.1751521, 0.02702342,
  0.2560489, 0.2476744, 0.3422548, 0.3569559, 0.1441335, 0.02513448, 
    0.1420196, 0.0537164, 0.1059398, 0.0893407, 0.06892809, 0.1222156, 
    0.3121661, 0.3014504, 0.3246397, 0.2847937, 0.2209506, 0.3055481, 
    0.2842721, 0.2876883, 0.3017313, 0.2451469, 0.2171015, 0.2021103, 
    0.1617696, 0.1525149, 0.1572896, 0.1656265, 0.2569574,
  0.1561754, 0.2354507, 0.2703831, 0.2877244, 0.2359327, 0.2203632, 
    0.1111652, 0.2260866, 0.2225129, 0.2034291, 0.2889862, 0.257536, 
    0.2489838, 0.2528824, 0.1634411, 0.1758461, 0.2357766, 0.2272695, 
    0.2062484, 0.2011534, 0.2447502, 0.2534424, 0.189663, 0.2686704, 
    0.1864466, 0.2176612, 0.1787227, 0.147316, 0.1417426,
  0.3141247, 0.2888469, 0.2111561, 0.2187869, 0.2033105, 0.2035022, 
    0.1913235, 0.2017928, 0.2528261, 0.2267886, 0.2027471, 0.149653, 
    0.1454412, 0.1547365, 0.1360668, 0.158836, 0.1583218, 0.1910231, 
    0.2059765, 0.1844899, 0.2060348, 0.1860697, 0.1804099, 0.1669192, 
    0.1467459, 0.2211404, 0.2701785, 0.2337707, 0.2516311,
  0.1311, 0.0844023, 0.04980304, 0.04359828, 0.05255952, 0.06575774, 
    0.08990961, 0.1200198, 0.09994908, 0.09373317, 0.07830071, 0.07299475, 
    0.04480751, 0.04340148, 0.02455117, 0.05399021, 0.1118157, 0.1504785, 
    0.1671005, 0.174749, 0.169113, 0.1353368, 0.1633558, 0.2939309, 
    0.04524007, 0.08674243, 0.1150478, 0.1574585, 0.1021952,
  0.01660032, 0.02883067, 0.05904864, 0.009266804, 0.06018434, 0.02732045, 
    0.0148407, 0.006679924, 0.003570422, 0.009430801, 0.00957855, 0.03396716, 
    0.07721656, 0.02720523, 0.07166688, 0.04750338, 0.1076836, 0.03707593, 
    0.1219845, 0.05259397, 0.01693314, 0.017317, 0.02434646, 0.007894686, 
    0.01123908, 0.102635, 0.02051035, 0.04056405, 0.03427345,
  9.411254e-05, -1.226878e-05, -1.390405e-09, 0.02863441, 0.04524016, 
    0.0007688461, 0.03316464, 0.0003359709, 2.761768e-06, 1.199431e-07, 
    5.898443e-08, 0.0007747949, 0.02153264, 0.07213951, 0.06256646, 
    0.01049182, 0.009555065, 0.008869105, 0.009295317, 0.001703684, 
    -3.614232e-05, 2.007977e-07, 2.092533e-07, 1.423223e-06, 0.0003526953, 
    5.453537e-05, 0.005564678, 0.02168243, 3.497913e-05,
  2.868713e-07, 1.347726e-05, 0.0004382392, 0.001197331, 0.01773623, 
    0.005346301, 0.04664655, 0.1410235, 0.02607444, 0.002234258, 0.009291438, 
    0.01339887, 0.09471424, 0.1641378, 0.1109493, 0.05080486, 0.04035664, 
    0.00272169, 0.0001927844, 1.37592e-07, 1.047893e-07, 1.276183e-06, 
    1.530296e-05, 0.001285968, -1.459141e-07, 7.446284e-07, 1.034959e-05, 
    0.0001513983, 2.464412e-07,
  0.02404265, 0.07531714, 0.0903655, 0.01158966, 0.001358294, 0.01029606, 
    0.03550877, 0.02577739, 0.1929297, 0.3271542, 0.05027501, 0.07394999, 
    0.06365144, 0.06011007, 0.06533984, 0.01279628, 0.01871915, 0.00249649, 
    0.01243327, 0.0002154209, 0.004644957, 0.0007781869, 0.02398743, 
    0.08222754, 0.1179044, 0.0574465, 0.03626201, 0.003296156, 0.0145153,
  0.1344925, 0.1819861, 0.1032224, 0.3023463, 0.006479893, 0.01934285, 
    0.05463676, 0.02938877, 0.06664902, 0.01414949, 0.009292117, 0.01843939, 
    0.0789597, 0.08143631, 0.07988983, 0.09912372, 0.06347841, 0.1125472, 
    0.1284843, 0.2790966, 0.4245274, 0.156141, 0.14728, 0.07807622, 
    0.06257866, 0.09449321, 0.115434, 0.2742575, 0.2874906,
  0.005556184, 0.005233871, 0.004144053, 1.372705e-05, 0.02023499, 
    0.07894266, 0.3537491, 0.2450832, 0.4067039, 0.04846621, 0.160787, 
    0.1158607, 0.1322217, 0.09550004, 0.009875672, 0.004249936, 8.363641e-05, 
    1.116195e-05, 0.004089525, 0.01390858, 0.0909209, 0.03265501, 
    0.006277608, 0.08748432, 0.01806386, 0.007860822, 0.00286004, 
    0.0002021393, 0.0006999666,
  7.140567e-05, 1.03098e-07, 3.903879e-10, 6.697066e-08, 6.768516e-05, 
    -0.0001531171, 0.05969002, 0.2518936, 0.2350975, 0.102915, 0.07457167, 
    0.04736397, 0.1752339, 0.1180892, 0.005901837, 0.03248294, 4.492849e-05, 
    2.321657e-05, 0.002229285, 0.001004593, 0.09662738, 0.04062183, 
    0.07814509, 0.1681332, 0.01939475, 0.002709952, 8.98771e-05, 
    7.980963e-07, 0.0001060674,
  0.01816689, 0.0003551972, 0.007019557, 0.003661208, 0.01013697, 
    0.006292236, 0.1636739, 0.01302685, 0.04760521, 0.08683397, 0.1313205, 
    0.1128568, 0.1357144, 0.2582327, 0.2140615, 0.05796207, 0.01963153, 
    0.03195649, 0.001637593, 0.0005838671, 0.01893559, 0.02760374, 
    0.09223662, 0.1744976, 0.1576614, 0.09906991, 0.0341469, 0.008692427, 
    0.002645853,
  0.05314085, 0.09112085, 0.03578827, 0.04644621, 0.02831908, 0.0884399, 
    0.09399106, 0.1045963, 0.1099656, 0.1758218, 0.08402917, 0.08316264, 
    0.133757, 0.04035996, 0.1131049, 0.1381582, 0.1315818, 0.1806716, 
    0.1175502, 0.07961787, 0.05811526, 0.06659224, 0.07774857, 0.1393855, 
    0.0977433, 0.07542832, 0.08729943, 0.1066606, 0.121111,
  0.2049336, 0.1722878, 0.1240169, 0.0607521, 0.01913857, 0.07578815, 
    0.1291027, 0.1566152, 0.07890051, 0.1057145, 0.09951381, 0.1304452, 
    0.1939064, 0.1340477, 0.1445295, 0.2286216, 0.2568335, 0.2435889, 
    0.3877924, 0.1872188, 0.06521714, 0.1145885, 0.146717, 0.137943, 
    0.1427896, 0.1541141, 0.08274138, 0.248465, 0.1580331,
  0.2362945, 0.2444815, 0.1725003, 0.1390241, 0.1087568, 0.08514935, 
    0.1053277, 0.165914, 0.08597123, 0.131601, 0.1155517, 0.1389903, 
    0.1141136, 0.0408311, 0.1191646, 0.09690624, 0.06521418, 0.05441142, 
    0.07775996, 0.06699381, 0.1542143, 0.1267718, 0.1874652, 0.1859804, 
    0.1538548, 0.2185275, 0.2085036, 0.2125928, 0.2316506,
  0.1123226, 0.1682227, 0.2384641, 0.1726177, 0.1381583, 0.1031066, 
    0.1182762, 0.07208581, 0.0550262, 0.1305293, 0.2216646, 0.2324044, 
    0.2743571, 0.3032396, 0.266511, 0.2717307, 0.3311886, 0.2396264, 
    0.1668777, 0.1565108, 0.1961799, 0.1931243, 0.2417262, 0.1355582, 
    0.2258713, 0.1777207, 0.1554924, 0.07085509, 0.08911664,
  6.10212e-05, 5.603315e-05, 5.10451e-05, 4.605704e-05, 4.106899e-05, 
    3.608093e-05, 3.109288e-05, 4.394443e-05, 3.547128e-05, 2.699814e-05, 
    1.852499e-05, 1.005184e-05, 1.578692e-06, -6.894455e-06, 2.094211e-05, 
    2.648026e-05, 3.201841e-05, 3.755657e-05, 4.309472e-05, 4.863288e-05, 
    5.417103e-05, 4.954218e-05, 5.746523e-05, 6.538828e-05, 7.331133e-05, 
    8.123438e-05, 8.915742e-05, 9.708047e-05, 6.501165e-05,
  -0.005564602, -0.0008649079, 0.004945267, 0.007221162, 0.001168615, 
    -0.0001366702, -0.0007175027, -0.001150642, 0.001674848, 0.006992616, 
    0.00220224, 0.00147763, 0.01540927, 0.1779604, 0.2305244, 0.2458083, 
    0.1849339, 0.2275886, 0.2024371, 0.1087025, 0.1374664, 0.06998155, 
    0.1625777, 0.1744549, 0.1803492, 0.1982604, 0.2597877, 0.2019849, 
    0.07661287,
  0.2542518, 0.2563049, 0.3679003, 0.3848339, 0.1686116, 0.05196764, 
    0.1420936, 0.05065398, 0.1323779, 0.1346375, 0.1252277, 0.1852319, 
    0.3232186, 0.345093, 0.3581384, 0.3029645, 0.2193518, 0.3397663, 
    0.3077143, 0.3311989, 0.3249866, 0.2483227, 0.2442478, 0.2251077, 
    0.1741155, 0.1382313, 0.1488173, 0.1537257, 0.2554685,
  0.1689648, 0.2260018, 0.2843355, 0.3019235, 0.2253972, 0.2071991, 
    0.1459582, 0.2272528, 0.2230627, 0.1885596, 0.288803, 0.2948971, 
    0.244209, 0.2619055, 0.1762947, 0.1815116, 0.2365675, 0.2337238, 
    0.1938097, 0.2076584, 0.2410209, 0.3286905, 0.2060238, 0.2697446, 
    0.1907844, 0.2276241, 0.2016859, 0.1559665, 0.1659622,
  0.3074983, 0.2914494, 0.2052042, 0.1974442, 0.2069099, 0.2009672, 
    0.2117245, 0.2371002, 0.2738319, 0.2261768, 0.2305461, 0.15084, 
    0.1456925, 0.1354239, 0.1553435, 0.1668218, 0.1572845, 0.195442, 
    0.1950294, 0.1783223, 0.2049377, 0.1994126, 0.1518774, 0.1651427, 
    0.1515651, 0.2218998, 0.2665946, 0.2072067, 0.2537259,
  0.1390741, 0.0852294, 0.05417729, 0.03781653, 0.05800898, 0.07455565, 
    0.09985734, 0.1421634, 0.1235307, 0.1078522, 0.09002895, 0.08178167, 
    0.04846266, 0.05412566, 0.02747509, 0.05360844, 0.1119807, 0.1515882, 
    0.1441218, 0.173841, 0.1545016, 0.1402907, 0.1799266, 0.2947718, 
    0.03634681, 0.09054435, 0.1086073, 0.152273, 0.1048677,
  0.01748932, 0.03230738, 0.06714876, 0.01120442, 0.0682262, 0.02635003, 
    0.02522684, 0.01034928, 0.005681707, 0.01323024, 0.03090546, 0.03457177, 
    0.1003282, 0.04098974, 0.07347098, 0.04315493, 0.1076576, 0.04105945, 
    0.129896, 0.06881975, 0.03247166, 0.03408407, 0.03647319, 0.00939865, 
    0.01687807, 0.1249554, 0.02255725, 0.04716226, 0.03289591,
  9.281914e-08, -8.095278e-05, 9.335652e-05, 0.03699205, 0.06509717, 
    0.01347358, 0.0503102, 0.0006133317, 6.350123e-07, 1.349725e-07, 
    2.928966e-07, 0.0002857194, 0.05291191, 0.06820339, 0.05326736, 
    0.005584977, 0.03576534, 0.01689736, 0.02365293, 0.001909877, 
    -1.634903e-05, 3.400315e-08, 1.433027e-07, 7.137092e-07, 0.003894442, 
    0.0003684965, 0.007283207, 0.01358224, -0.0002905588,
  3.549554e-07, 4.268551e-05, 0.0003840631, 0.001169874, 0.02803729, 
    0.005588823, 0.05014585, 0.1365902, 0.02861261, 3.677466e-05, 0.01825996, 
    0.04244435, 0.0984161, 0.1494089, 0.110866, 0.05624267, 0.055002, 
    0.00686861, 0.0002095865, 1.385208e-07, 2.059209e-07, 1.575469e-06, 
    1.842403e-05, 0.003437358, 1.765434e-05, 3.737813e-06, 0.002194066, 
    3.138102e-05, 2.173562e-07,
  0.01979688, 0.0872811, 0.1178102, 0.005355192, 0.000419506, 0.01092114, 
    0.03690201, 0.01940275, 0.1770243, 0.3462563, 0.04652901, 0.06328684, 
    0.05369797, 0.05261964, 0.04767304, 0.01286673, 0.006849804, 0.008164207, 
    0.006130821, 0.0001501196, 0.0008719699, 0.0002720203, 0.02506948, 
    0.1073924, 0.130315, 0.03936891, 0.03256562, 0.01154209, 0.02341009,
  0.1121538, 0.2002978, 0.08465032, 0.3869671, 0.002769745, 0.006610938, 
    0.03968035, 0.02576463, 0.04467707, 0.01111543, 0.007678389, 0.01459718, 
    0.06057673, 0.05976431, 0.06340799, 0.0866713, 0.07248516, 0.09408721, 
    0.1264328, 0.2637182, 0.3806334, 0.1308754, 0.1444976, 0.08347096, 
    0.05020476, 0.08985484, 0.08799195, 0.2488905, 0.298276,
  0.001694909, 0.001409886, 0.006168058, 5.983439e-06, 0.001261907, 
    0.05101377, 0.2660509, 0.2052059, 0.4308771, 0.04692092, 0.1351052, 
    0.103091, 0.08673515, 0.08128487, 0.01575295, 0.005683755, 0.0001285849, 
    6.165101e-06, 0.005061235, 0.002434913, 0.0560158, 0.03541117, 
    0.006016145, 0.08044504, 0.01429485, 0.00579378, 0.002712803, 
    7.081938e-05, 0.0005130056,
  1.996503e-05, 4.288845e-07, 6.158637e-09, 7.009896e-08, 2.633763e-05, 
    -5.050897e-05, 0.06893376, 0.3197962, 0.2733377, 0.09497022, 0.07460158, 
    0.04360461, 0.163734, 0.09921296, 0.005868562, 0.02998655, 3.682581e-05, 
    1.222317e-05, 0.0002380152, 0.0002492979, 0.09018495, 0.03001238, 
    0.05677337, 0.1506211, 0.01551615, 0.002647562, 0.0003864526, 
    5.296914e-07, 2.780432e-05,
  0.01609552, 0.001784377, 0.01982601, 0.007609759, 0.01348452, 0.001938552, 
    0.1593815, 0.003623365, 0.04253361, 0.08519035, 0.1361995, 0.09477902, 
    0.1432056, 0.2666099, 0.2481075, 0.07129143, 0.05241213, 0.02685019, 
    0.004955159, 0.0007984964, 0.003955392, 0.0456102, 0.1072057, 0.1855402, 
    0.1610398, 0.08029034, 0.07352633, 0.01232801, 0.001044052,
  0.06766441, 0.09221556, 0.03863577, 0.03916259, 0.0427973, 0.1040113, 
    0.09298683, 0.1012085, 0.09402251, 0.1651597, 0.0946961, 0.1197374, 
    0.1410725, 0.05058605, 0.1201278, 0.1702394, 0.1335823, 0.1970086, 
    0.1388623, 0.08095983, 0.06161872, 0.106621, 0.1069733, 0.1540779, 
    0.09507514, 0.08067767, 0.09078134, 0.1215665, 0.124128,
  0.1886291, 0.178012, 0.1510919, 0.08578125, 0.04035469, 0.07877707, 
    0.1340136, 0.1597995, 0.0806527, 0.115146, 0.119564, 0.1416413, 
    0.2267335, 0.1566227, 0.1478529, 0.2479916, 0.2319881, 0.3097502, 
    0.3445186, 0.1825541, 0.06577696, 0.1440698, 0.151577, 0.1798201, 
    0.1668967, 0.1432497, 0.06345002, 0.2028498, 0.1600532,
  0.2485748, 0.2329658, 0.1640965, 0.1490465, 0.1235316, 0.07183001, 
    0.1530821, 0.2185514, 0.08071874, 0.1280956, 0.1334113, 0.1351992, 
    0.08572756, 0.03280243, 0.08692253, 0.1092316, 0.07360844, 0.06875379, 
    0.06590761, 0.06904496, 0.1422694, 0.1403013, 0.2254018, 0.1524034, 
    0.2118438, 0.2298339, 0.1894223, 0.1951405, 0.1957813,
  0.08653636, 0.1714373, 0.2110778, 0.1764208, 0.1594073, 0.09739044, 
    0.134945, 0.08953972, 0.08120008, 0.1168354, 0.1893367, 0.2023716, 
    0.2368869, 0.2504158, 0.2479052, 0.2561157, 0.2396368, 0.1798672, 
    0.1434446, 0.1221951, 0.1876589, 0.1882293, 0.2544441, 0.1373503, 
    0.1839037, 0.1700745, 0.1418828, 0.07624424, 0.06018406,
  0.0004863774, 0.0004109764, 0.0003355754, 0.0002601744, 0.0001847735, 
    0.0001093725, 3.397148e-05, 0.000849969, 0.0006852715, 0.0005205739, 
    0.0003558764, 0.0001911788, 2.648126e-05, -0.0001382163, -0.001172759, 
    -0.001165145, -0.001157532, -0.001149918, -0.001142304, -0.001134691, 
    -0.001127077, -0.0006034635, -0.0003709786, -0.0001384937, 9.399122e-05, 
    0.0003264761, 0.0005589611, 0.000791446, 0.0005466982,
  0.03698276, 0.007683921, 0.02335577, 0.02845118, 0.01523767, 0.000616072, 
    -0.002094799, 0.004353263, 0.002495029, 0.007356497, 0.003472709, 
    0.01229887, 0.05168857, 0.1699825, 0.2275115, 0.2110008, 0.225478, 
    0.26105, 0.2146115, 0.1736351, 0.1983851, 0.1336632, 0.1832789, 
    0.1808785, 0.1803349, 0.2048319, 0.2597885, 0.1975124, 0.1071834,
  0.2614871, 0.2908301, 0.3892937, 0.4025167, 0.2216763, 0.08495287, 
    0.1421288, 0.1005758, 0.1565746, 0.1729846, 0.2348276, 0.2693487, 
    0.3017497, 0.381955, 0.3372428, 0.3366822, 0.27261, 0.3693376, 0.3612013, 
    0.3813394, 0.3660977, 0.3016147, 0.2363204, 0.3045279, 0.1743397, 
    0.134148, 0.1608039, 0.1433897, 0.2484934,
  0.1785344, 0.2477561, 0.2914795, 0.27872, 0.2151842, 0.2172389, 0.1519906, 
    0.2856499, 0.2956972, 0.1892038, 0.26662, 0.2788425, 0.2416506, 
    0.2606478, 0.1970176, 0.1939402, 0.2304955, 0.2687089, 0.2246847, 
    0.2290014, 0.2558917, 0.295235, 0.2384468, 0.3187476, 0.1985261, 
    0.2480432, 0.2049908, 0.1526868, 0.1892527,
  0.2953658, 0.2826312, 0.2127191, 0.2123468, 0.2130311, 0.2214312, 
    0.2530976, 0.2554799, 0.2690036, 0.2310913, 0.2489847, 0.164055, 
    0.1809987, 0.1596087, 0.179531, 0.1924365, 0.1544742, 0.1909171, 
    0.2070423, 0.1729687, 0.2038455, 0.2074042, 0.1573674, 0.1562598, 
    0.1450883, 0.2165241, 0.2784391, 0.1988384, 0.2372811,
  0.1435604, 0.08299501, 0.04937937, 0.04721094, 0.06526029, 0.08965333, 
    0.1070463, 0.1383539, 0.1358973, 0.1225296, 0.09727021, 0.1098921, 
    0.0660458, 0.05948947, 0.03128735, 0.06112703, 0.1091862, 0.1519821, 
    0.1331396, 0.1643889, 0.159546, 0.1373853, 0.1826154, 0.2893835, 
    0.02941741, 0.1003411, 0.1101002, 0.1625922, 0.1164983,
  0.02298374, 0.04039175, 0.07850467, 0.01587607, 0.07161576, 0.02964934, 
    0.02856366, 0.01634081, 0.008952927, 0.0149532, 0.03085868, 0.01876143, 
    0.1337156, 0.05417132, 0.0798213, 0.0480314, 0.1084796, 0.05795834, 
    0.1438758, 0.09561351, 0.04510847, 0.04766378, 0.03933263, 0.009642175, 
    0.03833642, 0.1433489, 0.03434559, 0.06768989, 0.04327864,
  9.503465e-08, 0.001518007, 0.003042984, 0.04288333, 0.07901049, 0.01386309, 
    0.06762951, 0.0003163479, -1.807182e-05, -3.055144e-07, -2.218015e-06, 
    2.92895e-05, 0.0530546, 0.07650515, 0.06413992, 0.005106387, 0.04173733, 
    0.01277428, 0.04619248, 0.006904599, 0.001306492, 7.893041e-08, 
    3.561274e-07, 8.43765e-07, 0.01040428, 0.004529273, 0.01609642, 
    0.01744502, 0.001468951,
  3.483088e-07, -0.0002214327, 0.0007971005, 0.004370248, 0.03055545, 
    0.01088411, 0.04255379, 0.1165509, 0.03186222, 0.001023889, 0.02213286, 
    0.04965357, 0.1052519, 0.1297919, 0.1017635, 0.06379973, 0.06136969, 
    0.01130814, 0.0003175336, 2.109228e-06, 3.278145e-07, 4.488191e-06, 
    4.925559e-05, 0.004015261, 0.001067301, 0.0004746208, 0.01070517, 
    4.311705e-05, 1.634146e-07,
  0.009273724, 0.08245603, 0.09638245, 0.003467964, 0.0003311202, 0.012052, 
    0.03480688, 0.01726547, 0.1345329, 0.2877602, 0.05342426, 0.05619683, 
    0.0458122, 0.04565385, 0.03853627, 0.01706462, 0.003417795, 0.0183467, 
    0.007959535, 0.000596726, 9.909978e-05, 0.0004385554, 0.02603091, 
    0.0983972, 0.1466028, 0.03338016, 0.01822556, 0.0176844, 0.0129413,
  0.06484806, 0.1316166, 0.0345091, 0.4487755, 0.001617068, 0.002831701, 
    0.03149458, 0.02431844, 0.0262388, 0.007805294, 0.007744259, 0.01293432, 
    0.04907269, 0.04702483, 0.05329804, 0.07833213, 0.06768963, 0.08257909, 
    0.12598, 0.2532775, 0.3224051, 0.1058297, 0.1161349, 0.07400112, 
    0.03167573, 0.07383983, 0.07431542, 0.2155288, 0.2393107,
  0.0002921502, 0.0002224141, 0.001255784, 1.75085e-06, 4.506136e-05, 
    0.02229687, 0.2086354, 0.195851, 0.3612755, 0.05008707, 0.121614, 
    0.1042631, 0.06639971, 0.0512358, 0.02467147, 0.01504217, 0.000188433, 
    0.0004071979, 0.007188231, 0.000215734, 0.04667814, 0.03681723, 
    0.006245327, 0.05473422, 0.01366881, 0.004154537, 0.001892397, 
    3.270258e-06, 0.0003202309,
  9.367195e-06, 1.593225e-07, -2.191759e-08, 5.558323e-08, 7.540038e-06, 
    -5.815195e-06, 0.06164301, 0.3536149, 0.3161135, 0.08595973, 0.07309115, 
    0.03822428, 0.1301039, 0.05120003, 0.007539166, 0.02067538, 0.0001285263, 
    -7.198054e-06, 1.64553e-05, 1.82795e-05, 0.03832794, 0.02341538, 
    0.04716175, 0.07235797, 0.01095828, 0.002880425, 0.0002681388, 
    1.994078e-07, 1.518714e-05,
  0.005679168, 0.002919833, 0.02125639, 0.008837771, 0.008959789, 
    0.005624408, 0.1188912, 0.0003033336, 0.03395101, 0.063868, 0.1211176, 
    0.08329264, 0.1390515, 0.2541493, 0.2005927, 0.06764852, 0.04725707, 
    0.05164439, 0.002336958, 0.0003364619, 4.765514e-05, 0.04572757, 
    0.1038827, 0.165527, 0.1497009, 0.09055159, 0.04311416, 0.01451967, 
    0.001288178,
  0.08571792, 0.1131132, 0.04198505, 0.04489064, 0.04485666, 0.09250963, 
    0.1013107, 0.1207231, 0.08988042, 0.1651052, 0.1042087, 0.1025635, 
    0.1356263, 0.08094084, 0.1175327, 0.1698456, 0.1721763, 0.21945, 
    0.1536284, 0.08894537, 0.07150888, 0.09959441, 0.1093014, 0.1761214, 
    0.09090878, 0.08791871, 0.09628152, 0.1370977, 0.1443264,
  0.2603121, 0.2211617, 0.1615885, 0.08749892, 0.05432168, 0.07837912, 
    0.1490598, 0.1845405, 0.095514, 0.1291907, 0.1614012, 0.1726009, 
    0.2653531, 0.1480339, 0.1625657, 0.2590201, 0.2188926, 0.3305614, 
    0.3623002, 0.1629488, 0.07984601, 0.1671478, 0.1747387, 0.1917184, 
    0.1633146, 0.1576783, 0.1079528, 0.2080957, 0.2121506,
  0.2202513, 0.2185651, 0.1877628, 0.1883355, 0.1408099, 0.08474327, 
    0.1328521, 0.1998589, 0.08295067, 0.1227994, 0.1340306, 0.1591169, 
    0.106268, 0.03991956, 0.07535286, 0.09817901, 0.07320983, 0.07102406, 
    0.06904497, 0.08763582, 0.1650942, 0.1217349, 0.2287558, 0.1674685, 
    0.1616582, 0.2756143, 0.1983728, 0.2082645, 0.2445542,
  0.1049576, 0.1759123, 0.2216516, 0.1801848, 0.1400556, 0.1158532, 
    0.1499874, 0.1053754, 0.1174668, 0.128612, 0.188674, 0.2282748, 
    0.2244668, 0.198134, 0.189091, 0.1608955, 0.23628, 0.1474912, 0.1672436, 
    0.1415216, 0.1809643, 0.1750533, 0.2400665, 0.1774521, 0.1877447, 
    0.14976, 0.1470054, 0.08588186, 0.1304193,
  0.009834158, 0.009580641, 0.009327124, 0.009073606, 0.008820089, 
    0.008566571, 0.008313053, 0.007977426, 0.007934829, 0.007892232, 
    0.007849636, 0.007807039, 0.007764442, 0.007721845, 0.003371346, 
    0.003489596, 0.003607846, 0.003726096, 0.003844346, 0.003962596, 
    0.004080846, 0.006370399, 0.006548263, 0.006726128, 0.006903992, 
    0.007081856, 0.00725972, 0.007437585, 0.01003697,
  0.08800703, 0.01513108, 0.02883951, 0.04521716, 0.02135108, 0.003475538, 
    0.002361006, 0.01175713, 0.01287631, 0.01101473, 0.005396258, 0.02534872, 
    0.07560405, 0.1661916, 0.2034707, 0.253172, 0.2732559, 0.2883182, 
    0.2111234, 0.2198755, 0.2470986, 0.1895353, 0.1856601, 0.1785712, 
    0.1887909, 0.199654, 0.2577813, 0.1861058, 0.1094543,
  0.28595, 0.3258466, 0.388105, 0.4397395, 0.2805269, 0.08239809, 0.1498482, 
    0.1266238, 0.2068719, 0.1904152, 0.2468518, 0.3179388, 0.2933137, 
    0.4103207, 0.3160565, 0.3084409, 0.2455788, 0.3548166, 0.372515, 
    0.3280368, 0.3539095, 0.297161, 0.2785314, 0.3132572, 0.1584633, 
    0.1316737, 0.1755278, 0.1519876, 0.2548006,
  0.1709017, 0.2424213, 0.2687089, 0.3197, 0.2796147, 0.2300929, 0.192516, 
    0.2986119, 0.2996382, 0.2081427, 0.2741029, 0.3234179, 0.2683048, 
    0.2960979, 0.2524752, 0.2442267, 0.2671298, 0.3006217, 0.2494344, 
    0.2889847, 0.3009522, 0.3210379, 0.2194814, 0.4219725, 0.193398, 
    0.266051, 0.235335, 0.1712585, 0.164685,
  0.3235727, 0.3200749, 0.2500322, 0.2234306, 0.2235077, 0.2415998, 
    0.2478574, 0.2777746, 0.2808716, 0.2427927, 0.2479301, 0.1805955, 
    0.2133797, 0.1813696, 0.1701612, 0.1961534, 0.164336, 0.2289637, 
    0.2103954, 0.1719059, 0.2281561, 0.1949238, 0.1683644, 0.1603519, 
    0.1783427, 0.2433527, 0.2827519, 0.2162009, 0.3185369,
  0.1488341, 0.09895765, 0.06443676, 0.05334888, 0.07149929, 0.1117654, 
    0.1329984, 0.1531041, 0.1434951, 0.1349876, 0.1217361, 0.1217287, 
    0.09441169, 0.07088733, 0.04275661, 0.08073647, 0.11649, 0.154283, 
    0.148267, 0.1673979, 0.1593593, 0.1567746, 0.1823904, 0.293529, 
    0.02807273, 0.1003501, 0.1310806, 0.1799384, 0.1336437,
  0.04033072, 0.03825384, 0.09894795, 0.02213612, 0.06285576, 0.02611442, 
    0.03714174, 0.02857602, 0.02126807, 0.0195843, 0.03337603, 0.007647347, 
    0.1684752, 0.06675899, 0.09399558, 0.05381148, 0.1138761, 0.07172196, 
    0.1512252, 0.1036589, 0.05732056, 0.07459891, 0.04209403, 0.01031995, 
    0.05647158, 0.176527, 0.04822085, 0.07124716, 0.05613513,
  -5.081444e-06, -3.073452e-05, 0.03670774, 0.05996899, 0.09217654, 
    0.04341106, 0.06863029, 0.007413235, 4.483981e-06, 1.542685e-05, 
    -0.0003060177, 0.009034782, 0.04588461, 0.1076071, 0.05915367, 
    0.003742369, 0.05566175, 0.007683326, 0.05924379, 0.02886258, 
    0.003618035, 3.531664e-05, 2.805697e-06, 8.182597e-07, 0.01758531, 
    0.02699488, 0.01886791, 0.0416675, 0.01119438,
  2.078003e-07, -7.478308e-05, 0.001369103, 0.01802435, 0.03611121, 
    0.01837421, 0.04315802, 0.1113707, 0.03275463, 0.002428126, 0.02926765, 
    0.04928836, 0.1259242, 0.1297307, 0.1014242, 0.070377, 0.07742494, 
    0.02692389, 0.002101482, 0.0001369486, 7.582075e-07, 2.450651e-06, 
    9.066401e-06, 0.009047788, 0.03791194, 0.02831936, 0.03904794, 
    9.675607e-05, 6.920901e-07,
  0.0007275696, 0.07432095, 0.09129095, 0.004622354, 0.0006908089, 
    0.01162559, 0.03103214, 0.01625804, 0.1136256, 0.2575042, 0.06138163, 
    0.04729483, 0.04205539, 0.04006108, 0.03256007, 0.02479453, 0.006807141, 
    0.00646131, 0.007832407, 0.0001337803, 9.682679e-05, 0.001521339, 
    0.03153948, 0.1236789, 0.158777, 0.04367742, 0.01588133, 0.007927725, 
    0.005969478,
  0.06038157, 0.09322841, 0.02035453, 0.4540641, 0.001776564, 0.003297548, 
    0.02990965, 0.02800931, 0.02100852, 0.006761719, 0.0119803, 0.01379947, 
    0.0437365, 0.03996575, 0.04933964, 0.0767324, 0.06089026, 0.07905347, 
    0.114708, 0.2450867, 0.2875464, 0.08999796, 0.1098595, 0.06748086, 
    0.02023943, 0.06958793, 0.0684449, 0.1978038, 0.2085616,
  6.690196e-05, 3.777665e-05, 1.277516e-05, 4.676313e-07, -8.219453e-07, 
    0.003803526, 0.1662093, 0.1939887, 0.363028, 0.05406557, 0.1121944, 
    0.1002284, 0.05236361, 0.0386825, 0.02783883, 0.03210843, 0.001412976, 
    0.003382464, 0.00986852, 4.225834e-05, 0.04203047, 0.04226065, 
    0.007207461, 0.0417005, 0.01454572, 0.003911771, 0.001068678, 
    2.589684e-07, 0.000169013,
  3.885525e-06, 6.59778e-08, 2.596539e-06, 2.507885e-08, 1.536797e-06, 
    -3.852992e-07, 0.05087523, 0.3728298, 0.3446206, 0.08235058, 0.08385432, 
    0.0314495, 0.109407, 0.0368978, 0.0125224, 0.01005966, -6.415635e-05, 
    -6.303014e-05, 3.67043e-06, 1.875064e-06, 0.01068763, 0.02501223, 
    0.04077126, 0.03842803, 0.01056367, 0.003879566, 0.001505135, 
    5.598787e-08, 1.049639e-05,
  0.0007376924, 0.007191128, 0.02458563, 0.02145897, 0.003211284, 
    0.003324839, 0.06962012, 6.645396e-05, 0.0212828, 0.05533055, 0.1166087, 
    0.07686377, 0.1334666, 0.2492121, 0.1764031, 0.07991722, 0.03302503, 
    0.03850698, 0.002655643, 4.307986e-05, 1.112852e-05, 0.03237909, 
    0.1084438, 0.1720434, 0.1388287, 0.05474851, 0.02449917, 0.0196388, 
    7.719122e-05,
  0.0811362, 0.1361981, 0.04636865, 0.04543107, 0.05161551, 0.08687826, 
    0.07995923, 0.1224383, 0.08937684, 0.1552556, 0.07480428, 0.09780771, 
    0.1015762, 0.06202921, 0.1271382, 0.16969, 0.1719529, 0.2627852, 0.16576, 
    0.1055222, 0.09436896, 0.08668379, 0.1068553, 0.2020191, 0.1095611, 
    0.1002771, 0.07791685, 0.1237702, 0.1335728,
  0.2921838, 0.2744916, 0.1712059, 0.08495747, 0.05013752, 0.06358708, 
    0.1470783, 0.201488, 0.1135591, 0.1459464, 0.1737044, 0.1976617, 
    0.289748, 0.144307, 0.1511026, 0.3057308, 0.2343587, 0.3804872, 
    0.4012727, 0.1746173, 0.1105314, 0.1897067, 0.1782798, 0.2104119, 
    0.1695766, 0.1704989, 0.1101227, 0.212637, 0.243765,
  0.2395497, 0.2514101, 0.2207682, 0.2054385, 0.1740086, 0.09616609, 
    0.2297909, 0.2134338, 0.09764275, 0.1506385, 0.1718151, 0.218684, 
    0.1139649, 0.04457895, 0.08969264, 0.09304778, 0.09419426, 0.07952099, 
    0.09183969, 0.1127504, 0.159315, 0.1265597, 0.2065172, 0.1357878, 
    0.1499743, 0.2307187, 0.2043507, 0.2148378, 0.2771946,
  0.09475278, 0.1685324, 0.2416072, 0.1700472, 0.1639248, 0.1185454, 
    0.1506965, 0.1509424, 0.09873345, 0.1218645, 0.1681347, 0.2190777, 
    0.265808, 0.2328942, 0.2031413, 0.2345607, 0.2326059, 0.1539318, 
    0.1556714, 0.1068423, 0.1780736, 0.1863522, 0.25904, 0.1362434, 
    0.1495233, 0.1427192, 0.1234624, 0.08227175, 0.07679629,
  0.02420903, 0.02415885, 0.02410866, 0.02405848, 0.02400829, 0.02395811, 
    0.02390793, 0.02178311, 0.02377613, 0.02576915, 0.02776217, 0.02975519, 
    0.03174821, 0.03374123, 0.02243379, 0.02012534, 0.0178169, 0.01550845, 
    0.0132, 0.01089156, 0.008583114, 0.01889409, 0.01925969, 0.0196253, 
    0.01999091, 0.02035652, 0.02072213, 0.02108774, 0.02424918,
  0.1042449, 0.04537813, 0.03109444, 0.03934005, 0.01736549, 0.002337854, 
    0.01467301, 0.01589445, 0.01739833, 0.01357926, 0.01804261, 0.02979654, 
    0.08120722, 0.1508806, 0.1698476, 0.2342084, 0.2773029, 0.293872, 
    0.1962076, 0.2222729, 0.2653565, 0.2095311, 0.1960797, 0.1850716, 
    0.1956569, 0.1920932, 0.2351216, 0.1796361, 0.1155571,
  0.3089519, 0.3719426, 0.3870873, 0.4381445, 0.3026825, 0.06815181, 
    0.1480909, 0.1710712, 0.2354678, 0.1957049, 0.2365073, 0.346156, 
    0.2964928, 0.378373, 0.2653602, 0.2378758, 0.2035067, 0.3861535, 
    0.2964977, 0.2744611, 0.2954105, 0.2514473, 0.2327148, 0.2496625, 
    0.1425987, 0.137531, 0.1611374, 0.1921431, 0.2499521,
  0.1626877, 0.2238621, 0.2996222, 0.342919, 0.2970634, 0.2669065, 0.1611032, 
    0.23804, 0.3095466, 0.2332249, 0.2712167, 0.3435539, 0.2537582, 
    0.2928213, 0.2694769, 0.250724, 0.2592168, 0.2713712, 0.2535493, 
    0.3079493, 0.3040603, 0.329784, 0.2340942, 0.402173, 0.2391156, 
    0.2518181, 0.2035527, 0.1642411, 0.1675376,
  0.3253003, 0.3484392, 0.2707959, 0.2485388, 0.2503115, 0.2783985, 
    0.2818663, 0.319688, 0.2939061, 0.2674906, 0.2696227, 0.211741, 
    0.2096555, 0.2009929, 0.214539, 0.2131155, 0.187748, 0.2432581, 
    0.2645081, 0.1730001, 0.219174, 0.2406008, 0.1780418, 0.1553511, 
    0.168158, 0.2441484, 0.3170947, 0.2267141, 0.3118314,
  0.1640305, 0.1112197, 0.0872499, 0.08699987, 0.09739672, 0.1444115, 
    0.1649518, 0.1761327, 0.1785835, 0.153598, 0.1506914, 0.1340373, 
    0.09287068, 0.09571219, 0.04940278, 0.1268576, 0.1317215, 0.1602987, 
    0.1669632, 0.1826237, 0.1774229, 0.1923309, 0.2003603, 0.3177326, 
    0.03146326, 0.10954, 0.1470541, 0.2098539, 0.1509524,
  0.06456529, 0.04777983, 0.1221538, 0.03127856, 0.06805677, 0.03616713, 
    0.04212279, 0.03397285, 0.03384773, 0.03141855, 0.03608886, 0.006576842, 
    0.1681546, 0.07026849, 0.108198, 0.07221089, 0.1222789, 0.07887252, 
    0.1655848, 0.1106641, 0.06058437, 0.08439758, 0.04801616, 0.0106271, 
    0.05122009, 0.1524286, 0.08816747, 0.07617936, 0.07325999,
  0.0001830478, -7.582688e-06, 0.1311731, 0.06187945, 0.08832645, 0.06158466, 
    0.07786919, 0.03005813, 0.0001550881, 0.0003226513, -0.0001236146, 
    0.01249545, 0.03410843, 0.1292921, 0.06637542, 0.00812145, 0.04636005, 
    0.009255108, 0.0635398, 0.09037223, 0.01216479, 0.005029297, 
    -3.655137e-05, 7.487211e-06, 0.01481456, 0.04615553, 0.04669938, 
    0.06398121, 0.01284398,
  1.418568e-07, -7.049938e-05, 0.008858553, 0.06390793, 0.04427182, 
    0.02442487, 0.0501846, 0.1085142, 0.03566374, 0.00618251, 0.04326054, 
    0.05514577, 0.1509698, 0.1407414, 0.09805162, 0.06566074, 0.07951943, 
    0.03424986, 0.01066429, 0.002070395, 5.556274e-05, 3.543981e-07, 
    1.307528e-06, 0.01046089, 0.03135809, 0.01625457, 0.1018964, 
    0.0009863471, 0.000217572,
  0.0001230786, 0.07305183, 0.08883251, 0.01627636, 0.00531624, 0.01699096, 
    0.02369588, 0.0168966, 0.08370265, 0.2504176, 0.06381024, 0.04509754, 
    0.03391308, 0.03640736, 0.02913282, 0.03276254, 0.0107459, 0.003530266, 
    0.00231143, 6.056169e-06, 6.909198e-05, 0.002501573, 0.02743752, 
    0.1532865, 0.1640681, 0.03155237, 0.01868205, 0.001444738, 0.002934042,
  0.05829674, 0.06692281, 0.01521696, 0.3696921, 0.0007864217, 0.004098078, 
    0.03071255, 0.03294111, 0.01915154, 0.007728058, 0.01598594, 0.0163045, 
    0.04140362, 0.03695738, 0.04661113, 0.07509778, 0.05793501, 0.08742343, 
    0.1228603, 0.2371505, 0.2633094, 0.09378738, 0.111535, 0.07368446, 
    0.01941415, 0.0706526, 0.07890195, 0.1995527, 0.184844,
  1.505991e-05, 6.593006e-07, 9.13103e-07, 1.282543e-07, -1.86278e-07, 
    -5.963895e-05, 0.1525042, 0.1794646, 0.3294579, 0.05489257, 0.09756494, 
    0.1002141, 0.044957, 0.03104721, 0.02533861, 0.03728535, 0.01162258, 
    0.008686012, 0.01159698, 7.293479e-05, 0.04455891, 0.04914015, 
    0.01035719, 0.02967812, 0.01875729, 0.006517634, 0.00105892, 
    -5.826026e-08, 9.128714e-05,
  1.983279e-06, 1.633284e-08, 2.928473e-08, 7.853433e-09, 5.439771e-07, 
    -4.635432e-08, 0.04230147, 0.3961515, 0.3325114, 0.08754871, 0.08618486, 
    0.02914201, 0.09893331, 0.03247873, 0.01636506, 0.01441069, 5.271968e-06, 
    -1.610036e-05, 5.259295e-07, 7.665226e-07, 0.002224738, 0.01988076, 
    0.03938849, 0.02329395, 0.01241738, 0.00872461, 0.003030116, 
    2.561529e-08, 7.328919e-06,
  0.0001434617, 0.006795278, 0.02527509, 0.02824285, -0.0002195836, 
    0.0001691057, 0.03897158, 2.214489e-05, 0.01177381, 0.0451502, 0.1185499, 
    0.07442547, 0.1357704, 0.2545028, 0.1639447, 0.07456188, 0.03127986, 
    0.03236245, 0.006644895, 4.825733e-05, -2.006958e-06, 0.01976716, 
    0.1131255, 0.1688897, 0.1327056, 0.04185268, 0.0248555, 0.02216992, 
    0.0001278058,
  0.07116724, 0.1337497, 0.04838366, 0.04392648, 0.02688533, 0.08848361, 
    0.07820745, 0.1394631, 0.1112321, 0.1272507, 0.06556001, 0.09414463, 
    0.1068314, 0.06763507, 0.1304087, 0.1818072, 0.2277365, 0.257978, 
    0.2031634, 0.1358082, 0.09623304, 0.08017783, 0.1135037, 0.2053385, 
    0.1452643, 0.115929, 0.09175125, 0.150248, 0.1406583,
  0.3185976, 0.3116463, 0.1667297, 0.09501541, 0.06099462, 0.1034902, 
    0.1672829, 0.2457862, 0.1028083, 0.1564314, 0.157019, 0.2398173, 
    0.2788859, 0.1353873, 0.1371177, 0.3756805, 0.3005206, 0.4183265, 
    0.4148272, 0.195061, 0.1337435, 0.2076014, 0.1938114, 0.2624035, 
    0.192424, 0.1941767, 0.1199705, 0.2353254, 0.3152981,
  0.263474, 0.2923789, 0.2327256, 0.1833718, 0.148579, 0.1095904, 0.2269396, 
    0.2425163, 0.1040537, 0.2108968, 0.193571, 0.2175772, 0.1163799, 
    0.05127943, 0.09522557, 0.1163148, 0.1517008, 0.08634269, 0.1199854, 
    0.1270029, 0.1533902, 0.1337089, 0.211522, 0.1201191, 0.1517395, 
    0.2181275, 0.1698272, 0.207219, 0.2989099,
  0.1097092, 0.1710905, 0.2274043, 0.2019676, 0.1843135, 0.1362004, 
    0.1394159, 0.1240542, 0.135711, 0.1748877, 0.1807051, 0.2410256, 
    0.3158686, 0.3222309, 0.2818795, 0.2936078, 0.2408062, 0.170949, 
    0.1648565, 0.1258354, 0.1903597, 0.2322512, 0.2652539, 0.1194612, 
    0.1310634, 0.1578656, 0.1312152, 0.07727046, 0.099273,
  0.04153079, 0.04124913, 0.04096748, 0.04068583, 0.04040417, 0.04012252, 
    0.03984086, 0.04257756, 0.04418289, 0.04578821, 0.04739354, 0.04899887, 
    0.0506042, 0.05220953, 0.03139702, 0.03022882, 0.02906062, 0.02789242, 
    0.02672422, 0.02555602, 0.02438782, 0.03902553, 0.03887006, 0.03871459, 
    0.03855911, 0.03840364, 0.03824817, 0.03809269, 0.04175611,
  0.1175527, 0.09448731, 0.03239055, 0.03508713, 0.015873, 0.002696326, 
    0.01861874, 0.01825076, 0.02493015, 0.02614595, 0.0389639, 0.03419447, 
    0.08316603, 0.140626, 0.1812806, 0.2060407, 0.208594, 0.2420582, 
    0.1807601, 0.2522069, 0.2739355, 0.2156336, 0.208192, 0.1924384, 
    0.198636, 0.1788869, 0.2323897, 0.1608024, 0.1124325,
  0.3133943, 0.3732938, 0.4134801, 0.4525236, 0.2870806, 0.0705682, 
    0.1490256, 0.2125452, 0.2535274, 0.1879566, 0.2491411, 0.3615896, 
    0.2955253, 0.3827877, 0.2981903, 0.2224704, 0.208504, 0.3545669, 
    0.2679451, 0.2923172, 0.26715, 0.2369742, 0.2064698, 0.2433943, 
    0.1227221, 0.104652, 0.1483719, 0.2125784, 0.2667073,
  0.1726362, 0.2513077, 0.3196073, 0.3620929, 0.2778939, 0.2630822, 
    0.1370094, 0.264544, 0.2714293, 0.2626845, 0.2720866, 0.3011823, 
    0.2582891, 0.2831005, 0.2880495, 0.2444269, 0.2354255, 0.2531116, 
    0.2586084, 0.2528463, 0.3065914, 0.2787042, 0.2272546, 0.3387079, 
    0.2410329, 0.2793268, 0.1690248, 0.161489, 0.186172,
  0.3105845, 0.3427542, 0.2798607, 0.308878, 0.2621099, 0.2765624, 0.3106926, 
    0.344539, 0.3085509, 0.2842429, 0.3601534, 0.1994938, 0.2605207, 
    0.2267459, 0.2382512, 0.2256955, 0.1872352, 0.2209735, 0.2488851, 
    0.2027878, 0.2264034, 0.2652384, 0.2192374, 0.1695461, 0.1387706, 
    0.2535815, 0.3181409, 0.2462296, 0.3016192,
  0.2047523, 0.1385408, 0.09381352, 0.1074694, 0.1277071, 0.1811973, 
    0.1866224, 0.2133567, 0.213602, 0.1716919, 0.1265491, 0.1186494, 
    0.08619605, 0.1118412, 0.0582516, 0.1535095, 0.1392058, 0.1750796, 
    0.1811896, 0.2113489, 0.1975, 0.2220771, 0.2198749, 0.3339892, 
    0.04436455, 0.1251252, 0.1763839, 0.2392451, 0.1806966,
  0.09819111, 0.06597614, 0.094232, 0.05535749, 0.05396168, 0.04955272, 
    0.04000823, 0.05577726, 0.04112349, 0.05953448, 0.04503024, 0.01465565, 
    0.1333971, 0.07449185, 0.09836094, 0.1061546, 0.1275544, 0.07676731, 
    0.1868561, 0.1255765, 0.0652476, 0.1059489, 0.05493397, 0.01281576, 
    0.05892926, 0.1085901, 0.08791748, 0.08491069, 0.08197021,
  0.002746131, 1.041259e-06, 0.04555992, 0.05838397, 0.07493526, 0.07028233, 
    0.06533838, 0.02585228, 0.005580198, 0.001280887, -6.920515e-06, 
    0.02328779, 0.02827144, 0.1717419, 0.1136184, 0.0169639, 0.03182294, 
    0.02469712, 0.06581105, 0.0895519, 0.09490421, 0.04649067, 0.005043412, 
    5.582537e-05, 0.01044074, 0.08837298, 0.07188798, 0.08500077, 0.03135016,
  1.090841e-07, -1.830973e-06, 0.02122852, 0.1307398, 0.03926616, 0.03074444, 
    0.06195433, 0.1163371, 0.03912461, 0.01342712, 0.07653077, 0.07551862, 
    0.155725, 0.1268666, 0.08494286, 0.05592812, 0.06922674, 0.02748052, 
    0.01853377, 0.009539546, 0.00287465, 2.092597e-06, 3.844574e-07, 
    0.01370843, 0.01833702, 0.001615321, 0.08122874, 0.009925109, 0.003233177,
  0.0002526789, 0.07228185, 0.05943276, 0.01571721, 0.01932478, 0.02411557, 
    0.017033, 0.016754, 0.07737262, 0.2436791, 0.06397036, 0.03872161, 
    0.02826042, 0.03210273, 0.02437872, 0.02896175, 0.01659289, 0.007675075, 
    0.00319089, 0.0004439472, 5.91742e-05, 0.001304671, 0.01139097, 
    0.1697635, 0.1575526, 0.02049313, 0.0189341, 0.003242953, 0.001576062,
  0.064132, 0.05954917, 0.01558276, 0.2928195, 0.000142048, 0.006279026, 
    0.03163688, 0.03216867, 0.01711775, 0.008237708, 0.0158733, 0.0196554, 
    0.03443157, 0.03242907, 0.04190401, 0.06642946, 0.05723887, 0.09296168, 
    0.120797, 0.2276451, 0.23271, 0.08521826, 0.1086882, 0.07538271, 
    0.01941375, 0.07502728, 0.09161635, 0.1919564, 0.1784597,
  5.284504e-07, 1.550276e-06, 3.312822e-07, 4.212777e-08, 1.243254e-07, 
    -0.0003478579, 0.156933, 0.1586915, 0.2916444, 0.04818649, 0.07290424, 
    0.09438122, 0.03903031, 0.02666921, 0.0215029, 0.04217032, 0.03747502, 
    0.009148891, 0.02038904, 0.001888136, 0.03599173, 0.05518845, 0.01213412, 
    0.02627865, 0.02860143, 0.01908517, 0.001127155, -1.129905e-06, 
    6.050349e-05,
  1.270799e-06, 1.82321e-09, 6.82138e-10, 1.748939e-09, 2.707118e-07, 
    -1.055845e-08, 0.03336025, 0.3843893, 0.3136548, 0.09489536, 0.08450131, 
    0.0308782, 0.09197284, 0.03037072, 0.02353913, 0.04887588, 0.00133635, 
    5.017378e-05, 1.343767e-07, 3.499961e-07, 0.0006039827, 0.01988654, 
    0.03918243, 0.01458523, 0.017494, 0.02727801, 0.008626094, 7.296362e-09, 
    5.646129e-06,
  1.141774e-05, 0.00678897, 0.02178438, 0.03918685, -0.0002383938, 
    -4.808995e-05, 0.02000777, 1.309516e-05, 0.003007655, 0.03658025, 
    0.1274602, 0.07331773, 0.1273754, 0.2612416, 0.1744285, 0.08248319, 
    0.05156034, 0.04601835, 0.008503235, 4.200372e-05, -7.197881e-08, 
    0.01408832, 0.1270133, 0.159527, 0.1253843, 0.03849282, 0.02864913, 
    0.04032417, 0.0001255009,
  0.08021943, 0.1389972, 0.05525259, 0.03843448, 0.02894687, 0.07494985, 
    0.07607696, 0.1483942, 0.1424308, 0.08990197, 0.06900144, 0.1019157, 
    0.1223174, 0.08688699, 0.1505423, 0.1639324, 0.2379827, 0.245664, 
    0.2032852, 0.1150848, 0.08669589, 0.08697343, 0.1199332, 0.2138086, 
    0.1962958, 0.1182946, 0.102255, 0.1555633, 0.1571041,
  0.291308, 0.309123, 0.1701196, 0.08910396, 0.06190821, 0.1229796, 
    0.1832018, 0.2414513, 0.09444366, 0.1504664, 0.1593094, 0.2395649, 
    0.2941088, 0.1606705, 0.1114677, 0.3895432, 0.3041286, 0.4365725, 
    0.4457498, 0.1927823, 0.1495247, 0.1998895, 0.1535584, 0.2724647, 
    0.2039302, 0.190418, 0.1519781, 0.2646391, 0.3257861,
  0.3057737, 0.3042549, 0.2572758, 0.1474385, 0.1153368, 0.09226201, 
    0.1831353, 0.2508015, 0.1223078, 0.2602477, 0.1810157, 0.2267711, 
    0.1056868, 0.06003891, 0.1022904, 0.1572971, 0.1556606, 0.07410739, 
    0.1592486, 0.1399509, 0.1586853, 0.1764595, 0.213149, 0.14649, 0.1236634, 
    0.2682529, 0.1695475, 0.194731, 0.3304425,
  0.1207877, 0.1827343, 0.2266618, 0.2284626, 0.2223434, 0.1322694, 
    0.1782461, 0.199218, 0.121549, 0.2130811, 0.2068989, 0.2655713, 
    0.3230916, 0.301685, 0.2669017, 0.2690756, 0.2391912, 0.1703275, 
    0.1861589, 0.1473579, 0.1779193, 0.2627572, 0.2329532, 0.1449747, 
    0.1342759, 0.1012328, 0.1378683, 0.0927113, 0.1015366,
  0.0599519, 0.0574755, 0.05499911, 0.05252271, 0.05004632, 0.04756992, 
    0.04509353, 0.05114345, 0.05258153, 0.05401961, 0.0554577, 0.05689578, 
    0.05833386, 0.05977194, 0.03680607, 0.0387275, 0.04064893, 0.04257037, 
    0.0444918, 0.04641324, 0.04833467, 0.06778579, 0.06690267, 0.06601956, 
    0.06513643, 0.06425332, 0.06337019, 0.06248707, 0.06193301,
  0.1174143, 0.1103957, 0.0487295, 0.03778814, 0.0161537, 0.003216708, 
    0.02585245, 0.02326344, 0.02469393, 0.04077611, 0.04177823, 0.03792898, 
    0.08829208, 0.1343202, 0.1897429, 0.2096207, 0.181144, 0.2011988, 
    0.1610461, 0.2530087, 0.2700796, 0.2312053, 0.2107918, 0.1902335, 
    0.1867083, 0.1757564, 0.2127497, 0.1548661, 0.1136274,
  0.3239068, 0.4062438, 0.4579467, 0.4378919, 0.2653407, 0.0693551, 
    0.1534395, 0.2432985, 0.2638682, 0.189111, 0.2595868, 0.3585841, 
    0.2934532, 0.3553317, 0.3011252, 0.2778558, 0.2072681, 0.3113575, 
    0.2797996, 0.2839604, 0.3252817, 0.2357183, 0.236245, 0.260568, 
    0.1091442, 0.1023006, 0.1432388, 0.2264588, 0.2439413,
  0.165379, 0.2350982, 0.4053652, 0.3869736, 0.2663128, 0.2378308, 0.1404404, 
    0.3176862, 0.2704773, 0.266143, 0.3204962, 0.3482256, 0.2816005, 
    0.3630576, 0.3411348, 0.2980366, 0.3305353, 0.286194, 0.3190327, 
    0.2474906, 0.3272606, 0.3057329, 0.2844765, 0.3568444, 0.2288646, 
    0.2977197, 0.1778718, 0.1963729, 0.1933036,
  0.3769823, 0.3574181, 0.3235915, 0.3119084, 0.2962312, 0.3329668, 
    0.3253905, 0.3817734, 0.3010985, 0.2865311, 0.3321761, 0.2121461, 
    0.2794837, 0.2471038, 0.2298893, 0.2485411, 0.2002872, 0.2276729, 
    0.2787956, 0.2547033, 0.2566252, 0.2495161, 0.2610138, 0.1831733, 
    0.1623346, 0.3002768, 0.3598292, 0.3588141, 0.3581886,
  0.2234235, 0.1796177, 0.1192935, 0.1424117, 0.1670213, 0.2192647, 
    0.2017187, 0.2495891, 0.219706, 0.1628508, 0.1400666, 0.132501, 
    0.09495911, 0.1231558, 0.06933331, 0.1563348, 0.1548093, 0.1890868, 
    0.1840302, 0.2392859, 0.2323784, 0.2271827, 0.2647683, 0.3520153, 
    0.06302852, 0.1725114, 0.2131265, 0.2423395, 0.1993455,
  0.1399437, 0.09043271, 0.06124198, 0.07846075, 0.06808724, 0.09155924, 
    0.0646079, 0.1091171, 0.0890393, 0.09366004, 0.03146793, 0.003717912, 
    0.1271001, 0.09285611, 0.09470058, 0.1198853, 0.147566, 0.1056852, 
    0.2718132, 0.1180391, 0.07142895, 0.1287023, 0.1187613, 0.01722682, 
    0.05685737, 0.1025421, 0.1551671, 0.115189, 0.1285386,
  0.06103488, -5.684281e-05, 0.01823025, 0.05747844, 0.0685095, 0.09388065, 
    0.08737095, 0.0500052, 0.02634846, 0.04622407, -1.126414e-07, 0.01473751, 
    0.05687881, 0.1729403, 0.1688192, 0.03121826, 0.07438961, 0.03791251, 
    0.07114585, 0.08340769, 0.1582908, 0.1224969, 0.06917335, 1.709001e-05, 
    0.00842564, 0.06845137, 0.06480176, 0.1631559, 0.111964,
  5.85465e-07, 1.654827e-07, 0.006733897, 0.1864751, 0.03957796, 0.04352364, 
    0.08603054, 0.1241007, 0.04317467, 0.0323306, 0.1047803, 0.08160125, 
    0.171052, 0.108527, 0.07980087, 0.04825477, 0.05956322, 0.02240926, 
    0.01768977, 0.01651417, 0.01022206, 0.000326559, 2.944005e-07, 
    0.02411866, 0.0009346543, -1.333348e-05, 0.06821835, 0.01857246, 
    0.009445826,
  0.001248498, 0.07961474, 0.04344067, 0.02524329, 0.02923985, 0.03119426, 
    0.01688517, 0.01637128, 0.06806241, 0.2196942, 0.06485083, 0.03438811, 
    0.0247906, 0.02922044, 0.02323682, 0.0273531, 0.02319616, 0.01056825, 
    0.009473994, 0.01035315, 0.0001541351, 0.006305535, 0.00534305, 
    0.1573125, 0.1534446, 0.01694163, 0.02067549, 0.01713199, 0.0001556096,
  0.06863698, 0.05780989, 0.01772691, 0.2425343, -8.595333e-05, 0.01221568, 
    0.03126558, 0.02896896, 0.01497517, 0.01009395, 0.0199405, 0.02524826, 
    0.02881275, 0.02988001, 0.03487124, 0.06238629, 0.06475259, 0.09747009, 
    0.1130051, 0.2012042, 0.1896992, 0.07609629, 0.106112, 0.07507995, 
    0.01992291, 0.06943428, 0.1020223, 0.176474, 0.1648028,
  -4.135556e-07, 6.510263e-07, 1.453709e-07, 1.574439e-08, 7.054425e-08, 
    0.0001921636, 0.1636253, 0.131033, 0.2567223, 0.04206142, 0.05027249, 
    0.08778045, 0.03480317, 0.02471023, 0.02007338, 0.05566309, 0.04052095, 
    0.04703996, 0.03050931, 0.00730391, 0.02769063, 0.05676787, 0.01234732, 
    0.02505506, 0.04752956, 0.04305165, 0.009871079, -2.035656e-06, 
    3.152156e-05,
  8.552262e-07, 1.467887e-09, 1.519081e-10, 5.210194e-10, 1.4101e-07, 
    -4.61184e-09, 0.02453114, 0.3634233, 0.3127403, 0.1033454, 0.07572381, 
    0.03748485, 0.08587222, 0.02652573, 0.02840263, 0.0791795, 0.02566292, 
    0.0005822345, 1.780165e-07, 1.729047e-07, 0.0002179156, 0.02063727, 
    0.04127416, 0.01230091, 0.01540813, 0.03968352, 0.04672586, 0.0001191792, 
    5.221843e-06,
  1.404411e-05, 0.00445404, 0.0205654, 0.06383795, -0.0001721484, 
    -6.243244e-06, 0.01320401, 8.196326e-06, -3.69277e-06, 0.03357911, 
    0.1445614, 0.07018617, 0.1356281, 0.2760902, 0.1879445, 0.08624342, 
    0.09164985, 0.09697821, 0.01739296, 2.396757e-05, 9.548188e-07, 
    0.01107016, 0.1414547, 0.1468957, 0.1185552, 0.0375873, 0.04973193, 
    0.06118519, 0.0005055424,
  0.1132726, 0.1435545, 0.1116928, 0.0290366, 0.01156814, 0.07958219, 
    0.0549435, 0.1373516, 0.1138283, 0.06536281, 0.07374967, 0.1332405, 
    0.1451866, 0.12272, 0.2141101, 0.1780191, 0.2702575, 0.3301311, 
    0.2561687, 0.1172108, 0.08783462, 0.124319, 0.1332869, 0.2189333, 
    0.1965956, 0.0978154, 0.1325718, 0.1787626, 0.2028609,
  0.3065972, 0.3095114, 0.170186, 0.07539239, 0.05755922, 0.09659051, 
    0.2082273, 0.231114, 0.1178438, 0.1621357, 0.1944555, 0.2397437, 
    0.3188943, 0.1974942, 0.129392, 0.3250569, 0.3037918, 0.4560021, 
    0.4439538, 0.1738313, 0.1425757, 0.2064856, 0.1709546, 0.2786216, 
    0.178385, 0.1978194, 0.214166, 0.3202942, 0.3587161,
  0.3529503, 0.3046509, 0.235248, 0.1463821, 0.1413095, 0.06951062, 
    0.1849132, 0.2778357, 0.1734216, 0.2910986, 0.1647542, 0.2772682, 
    0.1449385, 0.1275208, 0.1266782, 0.1353577, 0.159836, 0.07938658, 
    0.1678774, 0.1268478, 0.1997062, 0.158807, 0.2478486, 0.1742389, 
    0.1196813, 0.26548, 0.1925155, 0.2021146, 0.3238631,
  0.1500393, 0.2142359, 0.2434314, 0.2350481, 0.2228676, 0.2020058, 0.205897, 
    0.235214, 0.2451161, 0.3148325, 0.3068252, 0.3116042, 0.3134604, 
    0.2420195, 0.2684374, 0.2744828, 0.2647546, 0.178273, 0.1527111, 
    0.1939065, 0.1854034, 0.2597631, 0.2421097, 0.1573045, 0.1043144, 
    0.1283266, 0.1673378, 0.09193449, 0.1026794,
  0.08444641, 0.07964391, 0.07484141, 0.07003891, 0.06523641, 0.06043392, 
    0.05563142, 0.06204276, 0.06378279, 0.06552282, 0.06726284, 0.06900287, 
    0.0707429, 0.07248292, 0.06574182, 0.06860583, 0.07146984, 0.07433384, 
    0.07719785, 0.08006185, 0.08292586, 0.09477105, 0.09496951, 0.09516798, 
    0.09536644, 0.09556491, 0.09576337, 0.09596184, 0.0882884,
  0.09850796, 0.1200001, 0.0886455, 0.03846443, 0.01629112, 0.007063019, 
    0.03102008, 0.02815791, 0.03491709, 0.05982731, 0.04429134, 0.03996474, 
    0.1094581, 0.1351057, 0.2056293, 0.1984514, 0.1726324, 0.1724547, 
    0.1409387, 0.2225378, 0.2956904, 0.2574105, 0.2253045, 0.1700276, 
    0.1911714, 0.1599537, 0.1983762, 0.1380576, 0.1067242,
  0.3199783, 0.3878901, 0.4685925, 0.4122874, 0.2269058, 0.07560549, 
    0.1419359, 0.2629752, 0.2766571, 0.1824909, 0.2798927, 0.3477505, 
    0.2939612, 0.3111488, 0.3656216, 0.3134924, 0.2541043, 0.3411827, 
    0.3138069, 0.3226397, 0.3465465, 0.2986853, 0.2510172, 0.3003161, 
    0.0970918, 0.1057978, 0.1482401, 0.2606009, 0.2602901,
  0.1609178, 0.2674011, 0.5020806, 0.3839251, 0.3084693, 0.2935486, 
    0.1448932, 0.3667771, 0.3285321, 0.2878013, 0.362057, 0.3435564, 
    0.3533702, 0.4277431, 0.3677512, 0.3857247, 0.3822791, 0.3640762, 
    0.3705669, 0.3456773, 0.3914524, 0.3682684, 0.387091, 0.4233028, 
    0.3137926, 0.3193855, 0.2317917, 0.213316, 0.1859659,
  0.3982051, 0.3786434, 0.3370185, 0.366149, 0.3647557, 0.3220316, 0.3118268, 
    0.3640412, 0.2761344, 0.2868648, 0.2887603, 0.2615377, 0.2765525, 
    0.2581057, 0.2487523, 0.2337392, 0.2281914, 0.2557469, 0.3302714, 
    0.2877375, 0.3008795, 0.2715182, 0.2586104, 0.2111958, 0.2052995, 
    0.2908182, 0.4085958, 0.4027631, 0.414262,
  0.2427033, 0.2397004, 0.1255093, 0.2693053, 0.234267, 0.2784822, 0.236438, 
    0.248829, 0.2062422, 0.1401874, 0.160555, 0.1404893, 0.1106409, 
    0.1121798, 0.09720878, 0.142969, 0.1659447, 0.1902271, 0.1946802, 
    0.2159958, 0.2662509, 0.2339326, 0.3118542, 0.3966454, 0.1191592, 
    0.1779118, 0.1974003, 0.2089905, 0.1559013,
  0.1596695, 0.08350424, 0.0402008, 0.106587, 0.1791792, 0.1381618, 
    0.2054261, 0.2322352, 0.2242209, 0.1528692, 0.00369639, 0.001518349, 
    0.112896, 0.09637852, 0.1405058, 0.1447637, 0.1532722, 0.1506695, 
    0.2211283, 0.1065207, 0.1188696, 0.1163708, 0.2436923, 0.02501348, 
    0.06324864, 0.1026468, 0.1202024, 0.1668039, 0.1661571,
  0.2013285, -0.0002396994, 0.01236361, 0.07673471, 0.06838872, 0.1308646, 
    0.1316328, 0.1758032, 0.2840723, 0.07368901, -6.666033e-09, 0.001583681, 
    0.1404799, 0.1958259, 0.1327264, 0.0424656, 0.1120351, 0.04117883, 
    0.06920417, 0.1184315, 0.2499326, 0.3146389, 0.1396732, 1.139662e-05, 
    0.01784305, 0.03394982, 0.06377658, 0.2796758, 0.2843381,
  0.003346998, 1.768569e-06, 0.0005180232, 0.1448053, 0.04037832, 0.05031057, 
    0.1045004, 0.1187656, 0.04962408, 0.06186021, 0.1071895, 0.09833416, 
    0.1747472, 0.0818083, 0.0712058, 0.04327463, 0.05462604, 0.02797827, 
    0.02320523, 0.02592592, 0.0452771, 0.03052603, 1.868596e-06, 0.02075669, 
    0.00017059, -2.430315e-06, 0.07284308, 0.02784483, 0.03939357,
  0.0149116, 0.1406584, 0.03626895, 0.02256127, 0.03469145, 0.04202156, 
    0.01964672, 0.02104897, 0.05867608, 0.2086339, 0.06186474, 0.03093836, 
    0.02487963, 0.0262894, 0.02464538, 0.02901537, 0.01895732, 0.01140547, 
    0.01705217, 0.02883773, 0.004845226, 0.001280346, 0.003340413, 0.1596635, 
    0.1378452, 0.01793441, 0.02646766, 0.02933761, 0.005404915,
  0.08182753, 0.05475615, 0.01783961, 0.2184462, -0.0001651426, 0.02074165, 
    0.03095781, 0.02745713, 0.01400349, 0.01425184, 0.03465658, 0.03076537, 
    0.02608877, 0.02763037, 0.03641006, 0.05843265, 0.06099225, 0.0850177, 
    0.09948341, 0.1502142, 0.154708, 0.0644725, 0.1205417, 0.07334223, 
    0.02289017, 0.06018216, 0.1108237, 0.153524, 0.1519359,
  1.769672e-08, 3.785611e-07, 8.632754e-08, 9.874343e-09, 5.069325e-08, 
    0.003292219, 0.1477274, 0.1105599, 0.229884, 0.02980391, 0.03596738, 
    0.07635064, 0.03132876, 0.02674435, 0.02257366, 0.05195707, 0.1004166, 
    0.09709004, 0.05035239, 0.0098112, 0.02379607, 0.06264962, 0.01352885, 
    0.02412985, 0.05429965, 0.05406312, 0.034846, 1.091257e-05, 1.027473e-05,
  6.852812e-07, -2.163832e-10, 4.734276e-07, 2.984394e-10, 8.602989e-08, 
    -2.393994e-09, 0.01162071, 0.3406975, 0.3043703, 0.08652758, 0.06403486, 
    0.03934592, 0.07099991, 0.02492143, 0.03442675, 0.08168776, 0.09316055, 
    0.03814061, 1.320363e-06, 4.435053e-08, 0.0001157236, 0.02367721, 
    0.04306792, 0.01575516, 0.02159189, 0.03945569, 0.1108716, 0.01067111, 
    7.176471e-06,
  3.111112e-06, 0.002236175, 0.01771249, 0.08522506, -0.0001540431, 
    -2.515635e-06, 0.01189665, 9.515027e-07, -0.0001544498, 0.03270641, 
    0.1636695, 0.06943654, 0.1579859, 0.2873079, 0.2022397, 0.1326234, 
    0.1371803, 0.1325846, 0.03198652, 1.824014e-05, 1.703374e-06, 
    0.009746246, 0.1610254, 0.1598007, 0.1104315, 0.04869195, 0.05607904, 
    0.07868095, 0.009524122,
  0.1200111, 0.1262808, 0.09695091, 0.03026757, 0.01018103, 0.07427251, 
    0.0409924, 0.1168923, 0.09594315, 0.0472719, 0.07436942, 0.18002, 
    0.1532064, 0.1518193, 0.2297645, 0.2257252, 0.3312398, 0.4353907, 
    0.2584974, 0.1253154, 0.06125605, 0.09835237, 0.1135672, 0.2139332, 
    0.1658628, 0.133223, 0.1944579, 0.2525282, 0.2583622,
  0.3317819, 0.313054, 0.1764642, 0.08301263, 0.1261638, 0.08753454, 
    0.1989635, 0.2611364, 0.08890219, 0.1525041, 0.2352325, 0.2479221, 
    0.331747, 0.2383548, 0.1271777, 0.3318138, 0.3150129, 0.4687516, 
    0.3774291, 0.1429136, 0.1122082, 0.1998224, 0.1722506, 0.2815055, 
    0.1700779, 0.2028182, 0.2909139, 0.4641633, 0.4211095,
  0.37995, 0.2406861, 0.2136627, 0.1494586, 0.1904661, 0.1591422, 0.2515355, 
    0.2606926, 0.1646158, 0.3071594, 0.2033397, 0.2327683, 0.183519, 
    0.1384087, 0.1048787, 0.1175403, 0.1597858, 0.07582187, 0.1579998, 
    0.1403969, 0.1991325, 0.1688893, 0.2584451, 0.2097147, 0.1109982, 
    0.3175632, 0.1670643, 0.2274173, 0.3110128,
  0.1910687, 0.2718775, 0.3046767, 0.2901209, 0.2945119, 0.2605821, 
    0.2185208, 0.2109933, 0.3129495, 0.2853384, 0.3312885, 0.3283177, 
    0.4166022, 0.3317118, 0.388394, 0.3691134, 0.3229784, 0.2197751, 
    0.1567297, 0.2566472, 0.2297576, 0.3011577, 0.2532668, 0.159999, 
    0.1089566, 0.1429864, 0.1842641, 0.1067442, 0.1745204,
  0.1390322, 0.1334855, 0.1279387, 0.1223919, 0.1168451, 0.1112984, 
    0.1057516, 0.09069144, 0.09243388, 0.09417632, 0.09591876, 0.0976612, 
    0.09940364, 0.1011461, 0.09794988, 0.1011755, 0.1044011, 0.1076268, 
    0.1108524, 0.114078, 0.1173037, 0.1448486, 0.1454273, 0.146006, 
    0.1465847, 0.1471635, 0.1477422, 0.1483209, 0.1434697,
  0.0782954, 0.1083198, 0.1206205, 0.06540996, 0.02057202, 0.01552548, 
    0.03396347, 0.04422864, 0.04683832, 0.07237025, 0.06431613, 0.04424101, 
    0.1215716, 0.1318207, 0.2070855, 0.1941503, 0.1562539, 0.1374178, 
    0.1434425, 0.2000882, 0.3381819, 0.2822495, 0.2376538, 0.1652847, 
    0.1833381, 0.1416635, 0.2054348, 0.1110531, 0.08352374,
  0.2958495, 0.3515985, 0.4592991, 0.3608922, 0.1934476, 0.09557781, 
    0.09707972, 0.2701478, 0.2820952, 0.1825389, 0.2866223, 0.3298482, 
    0.2723016, 0.2827714, 0.3676395, 0.3313674, 0.2742254, 0.3645215, 
    0.3818301, 0.4110717, 0.3840867, 0.3374525, 0.2374161, 0.3651035, 
    0.08000997, 0.1125046, 0.1715677, 0.287037, 0.2644884,
  0.1763907, 0.3111776, 0.4927516, 0.329797, 0.2667077, 0.3331782, 0.1464008, 
    0.487138, 0.375019, 0.2788312, 0.3304305, 0.3344041, 0.3873877, 
    0.4269811, 0.2962211, 0.3268903, 0.3848522, 0.3858978, 0.3556487, 
    0.341063, 0.3888221, 0.3597575, 0.3651175, 0.4463759, 0.3919353, 
    0.3245717, 0.2702482, 0.2217062, 0.2171111,
  0.3923606, 0.40298, 0.4122528, 0.4296345, 0.406813, 0.3038518, 0.3177814, 
    0.2749594, 0.2674017, 0.2822899, 0.2705496, 0.2379189, 0.2876299, 
    0.2520421, 0.2821704, 0.2497412, 0.2086577, 0.2798621, 0.3316686, 
    0.3106461, 0.2893098, 0.2749071, 0.2394107, 0.2659256, 0.1953278, 
    0.3126676, 0.4135563, 0.3783826, 0.3886642,
  0.2311038, 0.2129654, 0.1104519, 0.2126978, 0.2344963, 0.2202015, 
    0.1932876, 0.2044946, 0.174189, 0.09815884, 0.1362834, 0.1164186, 
    0.1294152, 0.11758, 0.2583505, 0.1256795, 0.1472309, 0.2012244, 
    0.1578014, 0.2050315, 0.2556254, 0.2930498, 0.2302797, 0.4677492, 
    0.06908917, 0.1343842, 0.1609184, 0.1703007, 0.1312939,
  0.2232794, 0.07033428, 0.03607691, 0.1150927, 0.150784, 0.1185559, 
    0.296602, 0.2139701, 0.1444827, 0.1069951, 0.0009114144, 0.002121428, 
    0.09495602, 0.05387035, 0.1153874, 0.1112037, 0.1329634, 0.111219, 
    0.2091342, 0.1047846, 0.141139, 0.1401832, 0.2259068, 0.02630455, 
    0.0624913, 0.1301766, 0.1410384, 0.1031232, 0.1305198,
  0.3246144, -0.0008963922, 0.01029923, 0.08223926, 0.1009511, 0.1380702, 
    0.1420197, 0.2133476, 0.2683637, 0.02438805, -1.164603e-09, 0.0001847809, 
    0.09157342, 0.2479823, 0.1471047, 0.05450142, 0.1814075, 0.05302348, 
    0.07162384, 0.119848, 0.1627268, 0.320168, 0.3424256, -2.695207e-05, 
    0.03104746, 0.02665905, 0.05001596, 0.1996048, 0.2535698,
  0.02393292, 6.028822e-05, -0.0002634787, 0.08907054, 0.04723921, 
    0.06478196, 0.1091131, 0.1176975, 0.07207693, 0.1145601, 0.1295495, 
    0.09882487, 0.1861069, 0.06964322, 0.06886394, 0.04283519, 0.05252564, 
    0.05890953, 0.04341341, 0.04611992, 0.09755312, 0.1788553, 4.417846e-05, 
    0.02741843, 3.373239e-05, -8.685169e-07, 0.1065035, 0.04194393, 0.1816189,
  0.06688873, 0.1518477, 0.02587148, 0.02250995, 0.0405599, 0.07350293, 
    0.03381655, 0.04094023, 0.04604079, 0.1882914, 0.058906, 0.03203269, 
    0.02789035, 0.02729173, 0.02833249, 0.03756491, 0.0306266, 0.01685798, 
    0.01605579, 0.02354239, 0.04425302, 0.01155057, 0.003592071, 0.1808695, 
    0.1139638, 0.02232285, 0.05246334, 0.03592869, 0.03447543,
  0.08438178, 0.0466167, 0.01138549, 0.1962216, -0.0001730862, 0.0263171, 
    0.0287478, 0.03214498, 0.01112119, 0.02120876, 0.02373488, 0.04489935, 
    0.02619929, 0.02908201, 0.03839153, 0.06766208, 0.06718807, 0.07853013, 
    0.09492195, 0.1291653, 0.133989, 0.05575075, 0.1129475, 0.05979808, 
    0.03030434, 0.05737741, 0.1085633, 0.1356884, 0.1441508,
  1.581206e-07, 2.629939e-07, 6.237084e-08, 8.451917e-09, 4.51361e-08, 
    0.005758552, 0.1101501, 0.09612012, 0.1969551, 0.016851, 0.02950704, 
    0.06957617, 0.03583556, 0.03556281, 0.03572981, 0.05555573, 0.1391378, 
    0.1741162, 0.0720111, 0.02761328, 0.02031983, 0.06486852, 0.01753142, 
    0.02499252, 0.05524355, 0.07555044, 0.07568679, 0.0004303808, 2.55077e-07,
  5.93797e-07, -4.764716e-10, -4.639898e-11, 2.635669e-10, 5.666581e-08, 
    -1.526605e-09, 0.004614266, 0.3470452, 0.2958517, 0.07349955, 0.06003611, 
    0.07099833, 0.09564172, 0.02561029, 0.03833222, 0.09499618, 0.1506257, 
    0.1634463, 0.003464886, 1.295522e-07, 3.055298e-05, 0.02159577, 
    0.04277012, 0.0201909, 0.02737874, 0.0443453, 0.147912, 0.06088855, 
    -2.352115e-05,
  -1.650904e-05, 0.0004938584, 0.01701522, 0.1066115, -9.046376e-05, 
    -1.090775e-06, 0.01203392, 7.15914e-07, -0.0001281562, 0.02978243, 
    0.1874912, 0.07116355, 0.1528897, 0.3119336, 0.2231491, 0.211173, 
    0.2234685, 0.2621228, 0.185754, 6.55421e-06, 1.584069e-06, 0.004494554, 
    0.1528675, 0.1495135, 0.1370044, 0.08911276, 0.09076115, 0.1938001, 
    0.03127628,
  0.1118897, 0.0892358, 0.06844347, 0.02572111, 0.01012547, 0.06520817, 
    0.02865085, 0.09166484, 0.09095019, 0.03592687, 0.07036236, 0.1930572, 
    0.1781958, 0.1685401, 0.261672, 0.2924677, 0.4225106, 0.5164338, 
    0.3420287, 0.1019594, 0.05840571, 0.08678902, 0.0987473, 0.1982002, 
    0.1463072, 0.1886311, 0.2646654, 0.3275366, 0.3182002,
  0.3330655, 0.2731206, 0.1879663, 0.0579472, 0.08130514, 0.05261457, 
    0.1892007, 0.2470117, 0.07054625, 0.1243072, 0.2425873, 0.2573225, 
    0.3604486, 0.2667712, 0.1506554, 0.3846121, 0.2756642, 0.4542406, 
    0.343271, 0.1146804, 0.08806844, 0.1691904, 0.205982, 0.258557, 
    0.1636648, 0.174629, 0.3327022, 0.4750262, 0.4498554,
  0.496497, 0.2422126, 0.2224076, 0.150168, 0.1863918, 0.2084246, 0.341031, 
    0.2722147, 0.1557501, 0.3282374, 0.285469, 0.2800501, 0.1857401, 
    0.1310423, 0.1449758, 0.1514065, 0.1749934, 0.07875083, 0.1265913, 
    0.134544, 0.1868525, 0.2163383, 0.2699625, 0.2685389, 0.1125857, 
    0.3530452, 0.2181162, 0.257364, 0.4025623,
  0.3313595, 0.4074541, 0.4324322, 0.3473619, 0.3928224, 0.3162906, 
    0.3069598, 0.2754077, 0.3633613, 0.3255531, 0.3597022, 0.4008155, 
    0.5185685, 0.4398034, 0.4630664, 0.4190129, 0.3555679, 0.3328048, 
    0.2813699, 0.260488, 0.2921963, 0.3234585, 0.287611, 0.181284, 0.1167895, 
    0.153757, 0.1452802, 0.1192452, 0.2299224,
  0.1642184, 0.159615, 0.1550115, 0.1504081, 0.1458047, 0.1412012, 0.1365978, 
    0.1300755, 0.1310154, 0.1319552, 0.1328951, 0.1338349, 0.1347747, 
    0.1357146, 0.137502, 0.1402841, 0.1430661, 0.1458482, 0.1486302, 
    0.1514123, 0.1541943, 0.1566108, 0.1574924, 0.1583739, 0.1592554, 
    0.160137, 0.1610185, 0.1619001, 0.1679012,
  0.07852578, 0.1151201, 0.1177414, 0.08001711, 0.02630174, 0.01849694, 
    0.03670844, 0.05059768, 0.0441845, 0.07955635, 0.08736292, 0.06094813, 
    0.132438, 0.1235226, 0.2072541, 0.1819636, 0.1310061, 0.1054347, 
    0.1473177, 0.2010861, 0.3719546, 0.3148987, 0.2303051, 0.1552643, 
    0.1862418, 0.1440856, 0.2216881, 0.08721185, 0.07283626,
  0.2670684, 0.3194022, 0.4460277, 0.2670651, 0.150258, 0.1030974, 
    0.05541357, 0.2680224, 0.2800581, 0.1862259, 0.2968717, 0.3006954, 
    0.2489171, 0.2624879, 0.3404071, 0.3486291, 0.3321801, 0.420656, 
    0.4679423, 0.3946656, 0.3916322, 0.2969935, 0.2749689, 0.3994626, 
    0.06091537, 0.1287108, 0.1739647, 0.2811515, 0.3023556,
  0.1819401, 0.3088763, 0.4622976, 0.2741128, 0.290023, 0.3947661, 0.2336105, 
    0.5271591, 0.3103086, 0.2341161, 0.3041739, 0.3494633, 0.3593244, 
    0.3683781, 0.2233667, 0.2486109, 0.3681618, 0.422908, 0.3687567, 
    0.3090784, 0.3240359, 0.3380107, 0.277262, 0.4420553, 0.3895155, 
    0.3124048, 0.3439249, 0.2530235, 0.2780377,
  0.3773439, 0.4309731, 0.4696349, 0.4694091, 0.4221555, 0.3147838, 
    0.3067359, 0.1979394, 0.265837, 0.271374, 0.2777756, 0.2078345, 
    0.2556323, 0.1930821, 0.2542499, 0.2085685, 0.2235285, 0.2417204, 
    0.3191397, 0.3132904, 0.2616856, 0.2915042, 0.2280437, 0.2614222, 
    0.1650043, 0.3358302, 0.3803647, 0.3745343, 0.3616867,
  0.2040127, 0.1829785, 0.09548566, 0.1717834, 0.2039715, 0.1788937, 
    0.1866284, 0.1882977, 0.1698196, 0.1040956, 0.101473, 0.1067587, 
    0.05321858, 0.1156772, 0.3480175, 0.08730959, 0.1067381, 0.15643, 
    0.1221083, 0.2084232, 0.1936884, 0.2892828, 0.218483, 0.5335205, 
    0.04853464, 0.1101733, 0.146525, 0.153321, 0.1336811,
  0.1650915, 0.05245638, 0.04673729, 0.07467373, 0.1311983, 0.1048238, 
    0.122981, 0.08015405, 0.059578, 0.023935, 0.0001294736, 0.001510213, 
    0.06928956, 0.02707459, 0.05767605, 0.08628445, 0.1086342, 0.09038337, 
    0.1782784, 0.1070519, 0.08817922, 0.09690291, 0.2095736, 0.03753044, 
    0.0980171, 0.1249439, 0.1240938, 0.07631619, 0.07423109,
  0.2841078, 0.005629038, 0.00630046, 0.1682809, 0.06558159, 0.0708387, 
    0.06190715, 0.1824247, 0.159484, 0.01851379, -5.938789e-10, 8.791347e-06, 
    0.05791423, 0.2407992, 0.1772133, 0.09141073, 0.1353224, 0.08613775, 
    0.05643766, 0.04703536, 0.08058462, 0.1692346, 0.3373595, -0.001285838, 
    0.04336174, 0.02619073, 0.02212507, 0.08393694, 0.134503,
  0.2418727, 0.0005620997, 0.0002996615, 0.07456079, 0.04416224, 0.07632751, 
    0.1055122, 0.09827426, 0.05408322, 0.04994595, 0.08883014, 0.06820556, 
    0.1959013, 0.0707382, 0.06011943, 0.06533472, 0.05274458, 0.05352326, 
    0.03960609, 0.02481249, 0.0658442, 0.3099119, 0.1200458, 0.009861331, 
    4.150107e-06, -1.221477e-06, 0.04610145, 0.02960819, 0.2732853,
  0.2057713, 0.140984, 0.01052643, 0.02604453, 0.04701403, 0.1064611, 
    0.1213794, 0.0939533, 0.03471727, 0.1593481, 0.08694078, 0.08460546, 
    0.08438581, 0.04089239, 0.1092739, 0.0574813, 0.05147803, 0.0505928, 
    0.07043161, 0.05437358, 0.0511447, 0.0687331, 0.01179516, 0.1290323, 
    0.06653648, 0.03739606, 0.0607779, 0.06517135, 0.08183042,
  0.07564644, 0.03560017, 0.006054456, 0.181254, -0.0001078119, 0.0266894, 
    0.02591573, 0.0367769, 0.007638947, 0.06223587, 0.01516482, 0.1376392, 
    0.04112073, 0.03366721, 0.04335447, 0.06758612, 0.08712576, 0.1199043, 
    0.1315142, 0.1179023, 0.1436377, 0.06322797, 0.09515437, 0.0619072, 
    0.03776247, 0.06441651, 0.1043639, 0.1451406, 0.1143439,
  1.76609e-07, 7.978431e-08, 5.278467e-08, 6.297369e-09, 4.284627e-08, 
    0.02876776, 0.1028107, 0.08395779, 0.1516508, 0.01342281, 0.03034662, 
    0.06276472, 0.04280103, 0.03841776, 0.0319869, 0.04420527, 0.06836363, 
    0.2097639, 0.2319881, 0.08334727, 0.02648023, 0.07405649, 0.04780807, 
    0.01799269, 0.04933478, 0.1264136, 0.2427943, 0.008206213, -9.470634e-07,
  5.434379e-07, -4.727145e-10, -7.423902e-08, 6.157548e-11, 4.291964e-08, 
    -1.095983e-09, 0.001743388, 0.3584629, 0.2951187, 0.06116539, 0.06993056, 
    0.06915499, 0.1124124, 0.02369954, 0.05699369, 0.08370204, 0.1877768, 
    0.2716845, 0.2319609, 1.482603e-05, 1.965261e-05, 0.01319955, 0.02943879, 
    0.03250615, 0.05093879, 0.06791531, 0.1093515, 0.302552, -0.0001546344,
  -0.0001292783, 3.723031e-05, 0.01172492, 0.1262485, -8.461927e-05, 
    -4.51531e-07, 0.009660374, 6.275904e-07, -0.0001031359, 0.0259018, 
    0.1872663, 0.06336124, 0.173374, 0.3278976, 0.2767965, 0.3459804, 
    0.3783207, 0.3860998, 0.3621732, -2.646918e-05, 1.626671e-06, 
    0.0008240004, 0.1420066, 0.140475, 0.1333592, 0.1187149, 0.1690302, 
    0.378396, 0.05076766,
  0.123516, 0.06876892, 0.07714792, 0.02952908, 0.01027903, 0.06133291, 
    0.01848466, 0.09037982, 0.09740123, 0.03188402, 0.06151954, 0.1775338, 
    0.2222255, 0.2626923, 0.3216738, 0.3598891, 0.5095279, 0.5023623, 
    0.4039457, 0.09598241, 0.0548638, 0.0558785, 0.08508585, 0.1729004, 
    0.1424765, 0.2590086, 0.3420305, 0.4030271, 0.3647362,
  0.3129483, 0.2038944, 0.153076, 0.04505533, 0.05092646, 0.02616898, 
    0.1409092, 0.2064147, 0.05030562, 0.1029407, 0.2033096, 0.2857375, 
    0.3649671, 0.287865, 0.1748247, 0.4940506, 0.2554074, 0.4247097, 
    0.3264714, 0.09864586, 0.09591299, 0.1574681, 0.2075465, 0.2337915, 
    0.1588558, 0.1580573, 0.3745111, 0.4974894, 0.4486132,
  0.5667696, 0.2541797, 0.2474173, 0.156874, 0.2083676, 0.1858958, 0.3596599, 
    0.3008715, 0.1339396, 0.3418681, 0.267608, 0.2983179, 0.1486008, 
    0.1868207, 0.1972731, 0.2471132, 0.2478454, 0.1038075, 0.1149172, 
    0.1712934, 0.2711416, 0.2231023, 0.2549259, 0.2579896, 0.1015571, 
    0.3693063, 0.2301488, 0.3326674, 0.5434728,
  0.481971, 0.4684842, 0.4109285, 0.4124272, 0.3737672, 0.3722179, 0.4754738, 
    0.4405177, 0.4927392, 0.4605145, 0.4082858, 0.4492038, 0.5090842, 
    0.4332976, 0.4395225, 0.4046193, 0.3635748, 0.3383534, 0.3486082, 
    0.3781283, 0.3546233, 0.4090296, 0.2958198, 0.2110851, 0.1309302, 
    0.153422, 0.153973, 0.1388238, 0.4348211,
  0.2157677, 0.2129067, 0.2100456, 0.2071845, 0.2043234, 0.2014624, 
    0.1986013, 0.1826456, 0.1813609, 0.1800762, 0.1787914, 0.1775067, 
    0.176222, 0.1749372, 0.1600944, 0.1630578, 0.1660212, 0.1689846, 
    0.171948, 0.1749115, 0.1778749, 0.1819723, 0.1831546, 0.184337, 
    0.1855194, 0.1867018, 0.1878842, 0.1890666, 0.2180566,
  0.08349716, 0.1126601, 0.1243021, 0.082722, 0.03338293, 0.01861759, 
    0.03859127, 0.0497555, 0.03710808, 0.08571683, 0.1215094, 0.1000878, 
    0.1550826, 0.1013818, 0.2309711, 0.1501079, 0.1314013, 0.09638197, 
    0.1491543, 0.2307328, 0.4010349, 0.352947, 0.2239227, 0.1423846, 
    0.2003408, 0.1639424, 0.2100974, 0.06856304, 0.07225238,
  0.2463093, 0.3025615, 0.4122625, 0.1768219, 0.1166726, 0.09387223, 
    0.03289853, 0.2656706, 0.2724629, 0.1960288, 0.3056551, 0.2784183, 
    0.2251882, 0.2383333, 0.3439958, 0.3725888, 0.3858243, 0.4589153, 
    0.5289141, 0.3994271, 0.3992459, 0.2806065, 0.3135121, 0.4334411, 
    0.05382648, 0.1301562, 0.1858118, 0.2690183, 0.3086577,
  0.1748659, 0.300932, 0.3933959, 0.2843222, 0.2622209, 0.3544689, 0.2309732, 
    0.4585472, 0.2374981, 0.1886514, 0.2813746, 0.3617502, 0.3135364, 
    0.3063202, 0.200058, 0.2180461, 0.322246, 0.4311922, 0.3408347, 
    0.2956034, 0.3149967, 0.302237, 0.2444897, 0.4319316, 0.3169506, 
    0.3112072, 0.3403174, 0.3034102, 0.319305,
  0.3491898, 0.4426516, 0.4900311, 0.4654759, 0.4346734, 0.3194723, 
    0.2841668, 0.1636585, 0.2604268, 0.281687, 0.3123249, 0.2126735, 
    0.2166466, 0.1538766, 0.1780159, 0.1699615, 0.1823543, 0.2083524, 
    0.3001895, 0.2880416, 0.2325668, 0.276078, 0.1840402, 0.253441, 
    0.1371766, 0.307199, 0.3527821, 0.3468159, 0.3416736,
  0.1642302, 0.1213331, 0.07489721, 0.1341355, 0.1291368, 0.1391365, 
    0.1226172, 0.1537916, 0.1365059, 0.08028351, 0.07375767, 0.06287564, 
    0.02956231, 0.0769855, 0.294134, 0.07741578, 0.08851302, 0.1366886, 
    0.1184663, 0.2064733, 0.1700424, 0.2266092, 0.1954857, 0.5534292, 
    0.05075826, 0.09613861, 0.1484762, 0.1690314, 0.145578,
  0.1149964, 0.04989072, 0.04301288, 0.03989091, 0.05530841, 0.0475621, 
    0.04596836, 0.02950365, 0.03014174, 0.006370442, -2.160838e-05, 
    0.0002254515, 0.04826451, 0.01466226, 0.03141842, 0.05277791, 0.09767453, 
    0.0613647, 0.1712305, 0.07895049, 0.04563552, 0.05001119, 0.1122357, 
    0.03178335, 0.07352661, 0.1010593, 0.0781683, 0.04219645, 0.05847781,
  0.1485853, 0.02573799, 0.001691002, 0.05557417, 0.02570395, 0.02031431, 
    0.02389055, 0.1179872, 0.08049332, 0.004319106, -4.22459e-10, 
    -5.436834e-05, 0.02734576, 0.1440936, 0.1244931, 0.04960465, 0.0694199, 
    0.06037394, 0.03391265, 0.01287335, 0.03074058, 0.05571138, 0.2726784, 
    0.004266235, 0.04046459, 0.02094518, 0.001881842, 0.03015602, 0.06756582,
  0.4139042, 0.006972575, 0.0002349132, 0.05513525, 0.01803732, 0.06665941, 
    0.0769439, 0.05815808, 0.01161763, 0.01135268, 0.05970082, 0.02838198, 
    0.1549934, 0.07551435, 0.04617587, 0.02605092, 0.02414469, 0.01012778, 
    0.008836634, 0.006037467, 0.01877677, 0.130116, 0.2951162, 0.004125669, 
    6.388099e-07, -2.52611e-07, -0.0002220678, 0.008420042, 0.1079478,
  0.3029755, 0.08644567, 0.003736852, 0.0321078, 0.03653654, 0.03183645, 
    0.06439963, 0.03180792, 0.02846676, 0.1328605, 0.1432351, 0.1106844, 
    0.03937729, 0.03039056, 0.02352362, 0.01058944, 0.02304516, 0.01903751, 
    0.0301853, 0.03339645, 0.04073627, 0.3519694, 0.05333129, 0.06663053, 
    0.03823366, 0.01978536, 0.01638181, 0.03660234, 0.1355876,
  0.04791786, 0.0212345, 0.005085092, 0.1638921, -7.883459e-05, 0.009283442, 
    0.02283467, 0.01566887, 0.0006915394, 0.01713585, 0.005698514, 0.1147643, 
    0.1192972, 0.07075226, 0.02800272, 0.03891413, 0.0664052, 0.1039608, 
    0.08804407, 0.1259775, 0.1420615, 0.0802729, 0.1276402, 0.05521146, 
    0.02798358, 0.0557706, 0.1233604, 0.1637365, 0.08227985,
  1.639867e-07, 7.097665e-08, 4.738767e-08, 4.02951e-09, 4.216991e-08, 
    0.0826966, 0.1111953, 0.05995415, 0.1231019, 0.013219, 0.03064517, 
    0.03611825, 0.01959195, 0.0112452, 0.007189555, 0.01241491, 0.01732381, 
    0.08967883, 0.4749458, 0.303132, 0.06822872, 0.09682658, 0.008685282, 
    0.005099813, 0.01738778, 0.05275353, 0.2230795, 0.1153061, -4.39038e-07,
  5.098734e-07, -3.784359e-10, -1.06951e-05, -6.161898e-09, 3.447171e-08, 
    -9.311019e-10, -0.0017876, 0.3933712, 0.308703, 0.04532759, 0.1000945, 
    0.05593706, 0.1480552, 0.01895125, 0.03982176, 0.02401138, 0.1282935, 
    0.2353462, 0.5531787, 0.009177232, -1.223636e-05, 0.01124622, 0.0165336, 
    0.02982008, 0.09073, 0.1007989, 0.04675491, 0.2954982, -0.0007839623,
  -0.0003176719, 9.380402e-05, 0.01008804, 0.1335711, -5.270059e-05, 
    -1.126866e-07, 0.008126249, 5.612702e-07, -9.062472e-05, 0.02309189, 
    0.1696773, 0.06081315, 0.3467011, 0.4008149, 0.3815794, 0.5080291, 
    0.4712785, 0.3949598, 0.2753149, -0.0001520671, 1.420445e-06, 
    0.0002983857, 0.1106241, 0.1541678, 0.1483891, 0.09642575, 0.1646553, 
    0.3702347, 0.07955739,
  0.1359358, 0.04035765, 0.0528376, 0.02441473, 0.008445336, 0.04479026, 
    0.01401773, 0.09650066, 0.09640675, 0.03285249, 0.05035539, 0.1510848, 
    0.2609712, 0.3477926, 0.4991021, 0.5446634, 0.6295775, 0.5109337, 
    0.4689406, 0.1026901, 0.04666118, 0.04642961, 0.07226208, 0.1560631, 
    0.1348949, 0.3626712, 0.374121, 0.4840321, 0.4123681,
  0.3087487, 0.1780539, 0.1133687, 0.02861148, 0.02208064, 0.017837, 
    0.09594398, 0.1722654, 0.03131155, 0.0871266, 0.1749143, 0.2875716, 
    0.3893766, 0.3606611, 0.1731593, 0.6066753, 0.2486549, 0.3885383, 
    0.2771605, 0.08439001, 0.08805336, 0.1466809, 0.1979313, 0.2132199, 
    0.1981532, 0.1883592, 0.3830756, 0.4745339, 0.4640319,
  0.6200204, 0.2788228, 0.2068168, 0.211556, 0.259216, 0.1874737, 0.3245934, 
    0.2672449, 0.1049422, 0.3193146, 0.2593443, 0.2976359, 0.1593391, 
    0.1980869, 0.2315977, 0.3628074, 0.276162, 0.1259204, 0.1213318, 
    0.1751347, 0.3472109, 0.2279188, 0.2572161, 0.2399744, 0.1548207, 
    0.3623102, 0.2562665, 0.4277319, 0.7045257,
  0.6499484, 0.606909, 0.3933594, 0.5114208, 0.539441, 0.5147291, 0.6324663, 
    0.596788, 0.5775507, 0.5687795, 0.4798928, 0.4784828, 0.5060946, 
    0.4623311, 0.4288722, 0.4651518, 0.469806, 0.354436, 0.388586, 0.4792831, 
    0.4303123, 0.4886418, 0.2721379, 0.3467212, 0.1871643, 0.1506108, 
    0.1489286, 0.2273822, 0.5389452,
  0.2232485, 0.2196473, 0.2160461, 0.2124448, 0.2088436, 0.2052423, 
    0.2016411, 0.1924573, 0.19261, 0.1927627, 0.1929154, 0.1930681, 
    0.1932208, 0.1933735, 0.1935742, 0.1969726, 0.200371, 0.2037694, 
    0.2071678, 0.2105662, 0.2139646, 0.2253119, 0.225362, 0.2254122, 
    0.2254623, 0.2255124, 0.2255626, 0.2256127, 0.2261295,
  0.08397945, 0.09468019, 0.1136821, 0.07600796, 0.03597293, 0.01652369, 
    0.0374339, 0.04946839, 0.03795253, 0.09256129, 0.1066286, 0.1093779, 
    0.177486, 0.07399303, 0.2187161, 0.1492724, 0.1369403, 0.1247654, 
    0.1576414, 0.2381424, 0.3930561, 0.4063205, 0.2085953, 0.1379774, 
    0.2295996, 0.21259, 0.1988808, 0.06515906, 0.08271325,
  0.2392301, 0.2710469, 0.3678829, 0.1055857, 0.09514095, 0.08701802, 
    0.01636699, 0.2559188, 0.2595045, 0.1989647, 0.3062661, 0.278218, 
    0.1815902, 0.2090592, 0.372875, 0.3892459, 0.438808, 0.4676288, 
    0.4639089, 0.3719917, 0.3929717, 0.296132, 0.3204163, 0.4423927, 
    0.06733252, 0.1625599, 0.2215933, 0.2820893, 0.31912,
  0.2000558, 0.3120754, 0.3272939, 0.2649697, 0.2240829, 0.2538508, 0.221178, 
    0.3650373, 0.212019, 0.1601664, 0.2649999, 0.3441007, 0.2916641, 
    0.2766863, 0.1747494, 0.2076586, 0.2981153, 0.4087931, 0.3098434, 
    0.2631446, 0.2831788, 0.2702039, 0.2179528, 0.3528067, 0.2836391, 
    0.3254575, 0.3533736, 0.359868, 0.3200445,
  0.3175897, 0.4144691, 0.4516474, 0.4040198, 0.4305831, 0.3177034, 
    0.2515394, 0.1444848, 0.2389386, 0.2739635, 0.2648466, 0.1963522, 
    0.1959454, 0.1287942, 0.1387709, 0.1323014, 0.1295705, 0.1760993, 
    0.2638776, 0.244974, 0.1906036, 0.2295698, 0.1441402, 0.2311143, 
    0.132739, 0.2652619, 0.3129576, 0.3133283, 0.3407738,
  0.1502744, 0.07182356, 0.05002172, 0.09820139, 0.08380937, 0.1064751, 
    0.06956878, 0.0950264, 0.1039208, 0.05206832, 0.04925603, 0.03439236, 
    0.01253558, 0.04257361, 0.2344521, 0.05909288, 0.07231484, 0.1355672, 
    0.1152589, 0.1777185, 0.1537821, 0.1906682, 0.1416756, 0.5521268, 
    0.04267567, 0.07494661, 0.1326454, 0.1549032, 0.1170317,
  0.06405929, 0.04122926, 0.03188509, 0.03048116, 0.02346807, 0.01492425, 
    0.0151618, 0.01268215, 0.03864424, 0.002282487, -6.990377e-06, 
    -1.793721e-05, 0.03699724, 0.0102252, 0.01963039, 0.03415019, 0.09231026, 
    0.04639887, 0.1596441, 0.06644743, 0.02670041, 0.02658931, 0.04215565, 
    0.02903945, 0.04333415, 0.08578038, 0.0567908, 0.02509683, 0.02844921,
  0.06461665, 0.03001664, 0.0001929872, 0.01779891, 0.00886385, 0.006742476, 
    0.009375894, 0.07036747, 0.02559226, 0.001695377, -2.945334e-10, 
    -4.363656e-05, 0.006525387, 0.1004722, 0.0528871, 0.0192329, 0.02887271, 
    0.01311567, 0.01493062, 0.002973307, 0.01046445, 0.01953551, 0.1193166, 
    0.04279113, 0.01643964, 0.02970719, 0.0001651755, 0.01096772, 0.02022195,
  0.2018451, 0.06012417, 0.0001859101, 0.03914383, 0.006878107, 0.02086684, 
    0.04055375, 0.03149709, 0.0008534391, 0.001641342, 0.03271124, 
    0.005190252, 0.1298129, 0.04436664, 0.02876727, 0.008163332, 0.01058662, 
    0.0009676201, 0.0006690058, 0.0002234411, 0.003437308, 0.04001389, 
    0.2271173, 0.001013824, 9.317949e-08, 2.130199e-09, -0.002859869, 
    0.0002561941, 0.03648899,
  0.1127304, 0.07176763, 0.001545658, 0.0210014, 0.01676702, 0.009683507, 
    0.008236515, 0.005021572, 0.03393627, 0.0924153, 0.046, 0.02767202, 
    0.0153359, 0.005675589, 0.005410677, 0.001818988, 0.004029708, 
    0.003141825, 0.00915978, 0.01336003, 0.0227872, 0.2317209, 0.3561842, 
    0.04096536, 0.02742546, 0.001589634, 0.001173723, 0.007868723, 0.06434429,
  0.02789117, 0.02201011, 0.003004251, 0.1542622, -3.263538e-05, 
    0.0009980025, 0.03296485, 0.003839831, -0.002084055, 0.003498819, 
    0.001745478, 0.0210054, 0.02576323, 0.01497989, 0.01344026, 0.02263597, 
    0.02004371, 0.05240919, 0.03937458, 0.06847515, 0.1102782, 0.07191533, 
    0.1848269, 0.05413629, 0.006544027, 0.03160719, 0.08854365, 0.1044357, 
    0.06169613,
  1.54347e-07, 6.585739e-08, 4.465458e-08, 1.53781e-09, 4.145599e-08, 
    0.1095573, 0.09369701, 0.03807708, 0.1259628, 0.008785757, 0.01741312, 
    0.01846429, 0.005354896, 0.0007628291, 0.0007740529, 0.001277231, 
    0.003782979, 0.03253074, 0.2704875, 0.4807252, 0.1006134, 0.07788739, 
    0.0008788736, -0.0008863828, 0.00345199, 0.01434318, 0.0886322, 
    0.08511404, -5.127382e-08,
  4.865198e-07, -4.448522e-09, 0.0001170188, -3.136618e-08, 2.968125e-08, 
    -7.809237e-10, -0.003195308, 0.3816747, 0.3149649, 0.03944853, 0.0714955, 
    0.04766507, 0.06088017, 0.006441122, 0.00429628, 0.002642074, 0.03873057, 
    0.1690964, 0.3287258, 0.2674595, -1.697373e-05, 0.003837343, 0.009792316, 
    0.003723222, 0.01838882, 0.01635253, 0.005543944, 0.1766454, 0.003299479,
  -0.0004871464, 1.748297e-05, 0.0061805, 0.1533363, -4.343741e-05, 
    1.414712e-09, 0.006725254, 4.388496e-07, -8.253905e-05, 0.01982849, 
    0.1762733, 0.0835808, 0.4029107, 0.5398378, 0.4825345, 0.5538755, 
    0.3952184, 0.3143402, 0.3653571, -0.0001738996, 1.287233e-06, 
    0.0001186529, 0.08524115, 0.2383464, 0.173801, 0.109747, 0.1026209, 
    0.2175819, 0.07788102,
  0.1267636, 0.024497, 0.04283953, 0.01921435, 0.00460605, 0.02680516, 
    0.009365958, 0.1047008, 0.0787802, 0.03723836, 0.05606608, 0.1318594, 
    0.3733104, 0.4325558, 0.6896156, 0.704008, 0.6598687, 0.4946731, 
    0.3637418, 0.1035069, 0.03693135, 0.02759521, 0.06595303, 0.1435242, 
    0.1273105, 0.3965905, 0.3792161, 0.5020563, 0.4197465,
  0.2661173, 0.1662714, 0.08813128, 0.02202296, 0.01985196, 0.01386089, 
    0.07361067, 0.1360692, 0.02396361, 0.07727742, 0.1567933, 0.3089274, 
    0.4501532, 0.3965072, 0.2362633, 0.6806774, 0.2301728, 0.3756022, 
    0.2622066, 0.07060278, 0.0703942, 0.1293595, 0.2057526, 0.201638, 
    0.2621663, 0.208579, 0.3934357, 0.3914557, 0.4025229,
  0.6361969, 0.320728, 0.184459, 0.2522253, 0.3237232, 0.2474345, 0.3295867, 
    0.219651, 0.07014702, 0.271516, 0.2337313, 0.2925618, 0.1684213, 
    0.2133414, 0.2506035, 0.4030626, 0.2710906, 0.1658458, 0.2101368, 
    0.2068581, 0.3893789, 0.2447891, 0.219108, 0.2316979, 0.256508, 
    0.3538164, 0.2387829, 0.4081771, 0.7163323,
  0.6640461, 0.5878845, 0.4051805, 0.6236284, 0.6575892, 0.6214832, 
    0.5981843, 0.5750192, 0.5653905, 0.5468103, 0.4576463, 0.5482981, 
    0.5711424, 0.5231987, 0.4967948, 0.5013248, 0.5173043, 0.5202816, 
    0.52888, 0.5872384, 0.5383393, 0.547001, 0.2034039, 0.3781995, 0.2591447, 
    0.1473026, 0.1868518, 0.3915804, 0.5327128,
  0.1200811, 0.1160422, 0.1120033, 0.1079644, 0.1039255, 0.0998866, 
    0.0958477, 0.1026325, 0.1045213, 0.1064102, 0.1082991, 0.1101879, 
    0.1120768, 0.1139657, 0.125542, 0.1311807, 0.1368195, 0.1424582, 
    0.1480969, 0.1537356, 0.1593743, 0.1853548, 0.1818661, 0.1783774, 
    0.1748887, 0.1714, 0.1679114, 0.1644227, 0.1233122,
  0.08360814, 0.05772583, 0.0985506, 0.0649704, 0.03612576, 0.01623433, 
    0.02796021, 0.0428253, 0.02983061, 0.05083635, 0.03206352, 0.07065942, 
    0.1797609, 0.04931138, 0.2162351, 0.1487639, 0.1756874, 0.1897732, 
    0.2270315, 0.257445, 0.4540962, 0.4558477, 0.1787338, 0.1057413, 
    0.2923242, 0.2724985, 0.188257, 0.07568422, 0.08499543,
  0.2347103, 0.2426831, 0.3054936, 0.07456808, 0.06629381, 0.07864482, 
    0.008795464, 0.2133384, 0.236952, 0.1936702, 0.2984614, 0.2929691, 
    0.1391865, 0.1793493, 0.3969692, 0.432392, 0.4452255, 0.4948171, 
    0.400525, 0.342833, 0.3524344, 0.3369048, 0.3482977, 0.4758162, 
    0.06435632, 0.2151398, 0.307997, 0.3759548, 0.3578872,
  0.2660184, 0.3319994, 0.243092, 0.2207148, 0.1834518, 0.1957237, 0.2121835, 
    0.2933171, 0.1858492, 0.1484647, 0.2425016, 0.2992357, 0.2659169, 
    0.251716, 0.1358969, 0.191474, 0.2616846, 0.3628935, 0.2779585, 
    0.2195469, 0.2349035, 0.223751, 0.2072462, 0.3004831, 0.2711661, 
    0.3916283, 0.3776195, 0.4587819, 0.4006128,
  0.2880872, 0.3645189, 0.3739842, 0.3462655, 0.4129733, 0.3109035, 
    0.2116716, 0.1143586, 0.1931645, 0.2342248, 0.1931014, 0.1531505, 
    0.1476846, 0.08560296, 0.102591, 0.1097973, 0.0941404, 0.1363498, 
    0.201375, 0.2178779, 0.1518597, 0.1612921, 0.1171847, 0.1949451, 
    0.1116688, 0.234977, 0.289897, 0.2847106, 0.323849,
  0.1162435, 0.03741594, 0.04020609, 0.06205801, 0.05510078, 0.06546092, 
    0.04569121, 0.05290297, 0.07396163, 0.03441157, 0.04363761, 0.02060049, 
    0.00713977, 0.0312268, 0.1676329, 0.03965136, 0.05362372, 0.1229886, 
    0.08530233, 0.1437739, 0.1227296, 0.1442506, 0.1013372, 0.536672, 
    0.03053105, 0.05695266, 0.1026362, 0.1129393, 0.08771997,
  0.0233154, 0.01364893, 0.02555631, 0.007538101, 0.007388877, 0.006263459, 
    0.007789666, 0.006811851, 0.02054726, 0.001299975, -2.099076e-05, 
    -5.791535e-05, 0.0321454, 0.008285201, 0.01384225, 0.0229847, 0.0761375, 
    0.03381535, 0.1138149, 0.04674558, 0.01617715, 0.01255697, 0.02031544, 
    0.02524826, 0.03654753, 0.07287959, 0.03658905, 0.01262995, 0.01055616,
  0.0303767, 0.0305446, 6.004132e-06, 0.005659726, 0.002582669, 0.002876311, 
    0.003620746, 0.03657987, 0.008855238, 0.0009405608, -2.096707e-10, 
    -1.996264e-05, 0.001676313, 0.05496396, 0.02205509, 0.005235036, 
    0.01327098, 0.003114238, 0.00778426, 0.0004457895, 0.004754735, 
    0.00708185, 0.0448487, 0.03322171, 0.007153343, 0.03820553, 5.014545e-05, 
    0.005960157, 0.008564564,
  0.09726654, 0.07584259, 0.0007775322, 0.03079676, 0.002057372, 0.00784904, 
    0.01650919, 0.01329033, 0.00010893, -0.001087387, 0.01762101, 
    0.0004127026, 0.09676189, 0.01824692, 0.01168643, 0.002665912, 
    0.003602843, 0.0004054161, 0.0002779912, 7.585337e-05, 0.001433294, 
    0.0158565, 0.1012014, 0.0004853466, -2.964945e-07, 1.893002e-08, 
    -0.001492736, 1.43126e-05, 0.01496144,
  0.03999783, 0.05698816, 0.0007019923, 0.01172426, 0.002194336, 0.001961957, 
    0.002401889, 0.001166089, 0.02956918, 0.07401447, 0.0123916, 0.00554206, 
    0.002954651, 0.00204097, 0.003080835, 0.0007571859, 0.0008186882, 
    0.0004176315, 0.001320459, 0.00161278, 0.002824394, 0.0777131, 0.2061549, 
    0.03451915, 0.02215542, 0.0002413713, 0.0001566345, 0.00066204, 0.01241263,
  0.02080987, 0.02917074, 0.002006221, 0.1532293, -1.620985e-06, 
    5.349335e-05, 0.04504694, 0.0001703748, -0.002001885, 0.0009616798, 
    0.0002445064, 0.006294259, 0.006224622, 0.003068494, 0.005430043, 
    0.01083407, 0.008657827, 0.0131487, 0.02988728, 0.03385105, 0.05951716, 
    0.02807068, 0.2092848, 0.03767897, 0.0004480894, 0.01068458, 0.02231238, 
    0.04963952, 0.05867331,
  1.501621e-07, 6.227508e-08, 4.290424e-08, 7.844168e-10, 4.038037e-08, 
    0.01200036, 0.05779286, 0.01849827, 0.1332177, 0.003156791, 0.002639866, 
    0.006302902, 0.0005429381, 4.526089e-06, 4.52183e-05, 6.813916e-05, 
    0.001247887, 0.01471319, 0.1453475, 0.3467221, 0.02584041, 0.06270715, 
    0.0002794519, -0.002696885, 0.0007342873, 0.004103048, 0.03089235, 
    0.06251338, 1.101433e-07,
  4.698148e-07, -3.132223e-07, 0.0002767594, -1.241543e-07, 2.641673e-08, 
    -6.785248e-10, -0.001365272, 0.3550223, 0.3088551, 0.03232703, 0.0795111, 
    0.02133249, 0.02361759, 0.001065574, 0.0006377498, 0.0005569693, 
    0.01473139, 0.07424743, 0.145372, 0.2903568, 1.074006e-05, 0.001288867, 
    0.005936213, 0.0007497424, 0.005178608, 0.006162548, 0.001171968, 
    0.08091333, 0.006742094,
  -0.0005887075, 1.024346e-05, 0.002160454, 0.1717376, -4.494232e-05, 
    2.483771e-08, 0.004707202, 4.706955e-07, -6.483342e-05, 0.01520379, 
    0.196753, 0.09747232, 0.5287007, 0.6320807, 0.6243804, 0.3925393, 
    0.272512, 0.2191657, 0.2646734, -0.000613716, 1.184922e-06, 3.86709e-05, 
    0.07021581, 0.2659445, 0.1426411, 0.1168954, 0.05043345, 0.1157602, 
    0.06686284,
  0.1282435, 0.02269769, 0.04068715, 0.01417057, 0.002028594, 0.01133061, 
    0.005652801, 0.09462227, 0.07091412, 0.04220041, 0.04888555, 0.1264987, 
    0.6274477, 0.5038415, 0.7889193, 0.671948, 0.6614916, 0.428477, 
    0.2990535, 0.1023355, 0.024392, 0.01633787, 0.05677654, 0.1285886, 
    0.1242203, 0.450987, 0.3693551, 0.5066249, 0.4175797,
  0.1956001, 0.14782, 0.07155818, 0.01459715, 0.0128968, 0.009879913, 
    0.05931268, 0.1114599, 0.01442217, 0.06274643, 0.1431481, 0.3303479, 
    0.4714952, 0.3778697, 0.3583522, 0.7067556, 0.2192705, 0.341822, 
    0.239728, 0.06410912, 0.05265344, 0.119773, 0.2183615, 0.1768363, 
    0.2907936, 0.1969324, 0.3365478, 0.3162823, 0.3028432,
  0.5979961, 0.3532441, 0.1649766, 0.2149337, 0.3455572, 0.2488898, 
    0.3200896, 0.1808263, 0.05440015, 0.2304734, 0.1883279, 0.2735039, 
    0.161642, 0.2320882, 0.3727695, 0.3785012, 0.2634764, 0.2899865, 
    0.2919892, 0.2589802, 0.3931771, 0.3034964, 0.1936868, 0.1897642, 
    0.3536792, 0.3402502, 0.2024314, 0.3588312, 0.6670461,
  0.5407155, 0.4519178, 0.4975023, 0.589817, 0.6187246, 0.623868, 0.5444843, 
    0.5016699, 0.5268529, 0.4974583, 0.4967321, 0.6231439, 0.6733866, 
    0.5689744, 0.5347598, 0.5369877, 0.576857, 0.5872586, 0.5527424, 
    0.5196217, 0.5992894, 0.5213636, 0.1556297, 0.3033219, 0.281722, 
    0.175845, 0.1944402, 0.4735162, 0.434123,
  0.03526216, 0.03352587, 0.03178957, 0.03005327, 0.02831697, 0.02658067, 
    0.02484437, 0.01848728, 0.0226525, 0.02681772, 0.03098294, 0.03514816, 
    0.03931338, 0.0434786, 0.04788874, 0.04964246, 0.05139618, 0.05314989, 
    0.0549036, 0.05665732, 0.05841104, 0.06376018, 0.05957755, 0.05539491, 
    0.05121228, 0.04702965, 0.04284701, 0.03866438, 0.03665121,
  0.06743748, 0.05211816, 0.06984687, 0.05106279, 0.02419188, 0.02051468, 
    0.02575105, 0.05660721, 0.008769364, 0.00882257, 0.01983142, 0.06720608, 
    0.1595159, 0.02207967, 0.2312839, 0.2454449, 0.2002462, 0.2146919, 
    0.2318533, 0.3043006, 0.489147, 0.5188637, 0.1105591, 0.07735156, 
    0.3012301, 0.3599666, 0.1617505, 0.07191543, 0.08265244,
  0.2091282, 0.2043533, 0.2434098, 0.05408188, 0.03986508, 0.07359525, 
    0.004264153, 0.1565253, 0.2363753, 0.1793556, 0.2446803, 0.2807811, 
    0.1033059, 0.1573431, 0.3893532, 0.4270184, 0.4237675, 0.4138163, 
    0.3249751, 0.3192123, 0.3115044, 0.3285317, 0.3420495, 0.4879681, 
    0.05316578, 0.2686034, 0.3622423, 0.4667179, 0.3849453,
  0.3110683, 0.3137497, 0.1799081, 0.1758564, 0.1389531, 0.1504959, 
    0.2225314, 0.2406644, 0.1586812, 0.1188455, 0.2176105, 0.2497294, 
    0.2263502, 0.2197512, 0.109191, 0.1621632, 0.2243974, 0.3140047, 
    0.2426093, 0.1654528, 0.1836343, 0.1755183, 0.1740591, 0.2539314, 
    0.2621957, 0.4190674, 0.4218733, 0.4989216, 0.4236468,
  0.2469431, 0.2905945, 0.3017129, 0.3082385, 0.375931, 0.2641644, 0.1661657, 
    0.08270784, 0.1453496, 0.1759304, 0.1337195, 0.1037056, 0.09723265, 
    0.05444298, 0.05937598, 0.08428872, 0.06045028, 0.09905908, 0.1384218, 
    0.1571793, 0.1156687, 0.1192163, 0.09122994, 0.1562932, 0.08893543, 
    0.1987508, 0.2526004, 0.2289788, 0.2824515,
  0.07818455, 0.02185335, 0.02880314, 0.03666565, 0.03436575, 0.03720627, 
    0.02329814, 0.02952051, 0.0463324, 0.0231009, 0.03765719, 0.0107711, 
    0.003710956, 0.0233059, 0.1220917, 0.02579503, 0.03970509, 0.103487, 
    0.06321043, 0.1113158, 0.09124792, 0.1048418, 0.066045, 0.5048783, 
    0.02563305, 0.04003458, 0.07808771, 0.0704811, 0.05930728,
  0.01200804, 0.004259807, 0.02067907, 0.003255332, 0.002935835, 0.003359696, 
    0.005195982, 0.00469897, 0.008289221, 0.0008824443, -2.66113e-05, 
    -3.356137e-05, 0.0259612, 0.005023316, 0.008407537, 0.01468982, 
    0.05236106, 0.02086589, 0.07768732, 0.024061, 0.01019531, 0.005695479, 
    0.01238254, 0.0139512, 0.03060425, 0.03715118, 0.01403897, 0.005691668, 
    0.005747661,
  0.01765648, 0.01993892, -3.272754e-06, 0.002848399, -0.0006310969, 
    0.001103155, 0.001473325, 0.01938906, 0.004383745, 0.0006112394, 
    -1.946074e-10, -6.363587e-06, 0.0008651583, 0.02418051, 0.0105325, 
    0.002352965, 0.007503755, 0.001408625, 0.003604766, 0.0001535073, 
    0.002006879, 0.003489055, 0.02309251, 0.02419768, 0.004610726, 0.0433674, 
    2.710995e-05, 0.002522657, 0.00481145,
  0.05460936, 0.06172686, 0.001033819, 0.02159004, 0.00022172, 0.001916688, 
    0.006562949, 0.004011713, 6.195206e-05, -0.0009128869, 0.01191112, 
    0.0001687032, 0.0503599, 0.006158267, 0.004116661, 0.000872585, 
    0.001280698, 0.0002320074, 0.0001571417, 3.579858e-05, 0.000802712, 
    0.008446322, 0.05857161, 0.0004857443, -6.005466e-06, 1.625375e-08, 
    -0.0009383007, -2.929012e-06, 0.008226463,
  0.01977927, 0.04633877, 0.0003686173, 0.005759589, 0.0001740354, 
    0.0008264721, 0.00124574, 0.000598037, 0.02982387, 0.08634491, 
    0.004460125, 0.002465642, 0.001081535, 0.0008526587, 0.001743376, 
    0.0004619703, 0.0004121624, 0.000201135, 0.0006413727, 0.0003664576, 
    0.0004141021, 0.0315707, 0.1131526, 0.0426797, 0.03236528, 0.0001251614, 
    6.811701e-05, 0.0002900444, 0.004716944,
  0.01548436, 0.02712905, 0.001149497, 0.1543195, -1.287033e-06, 
    1.729794e-05, 0.03385627, 2.324899e-05, -0.0007468487, 0.0004661131, 
    3.472393e-05, 0.003146798, 0.002877575, 0.0008405857, 0.002569191, 
    0.004890042, 0.005153025, 0.00562129, 0.02253017, 0.014443, 0.02434824, 
    0.009424506, 0.1759592, 0.02761297, 6.646368e-05, 0.0061615, 0.009788066, 
    0.02384447, 0.04758951,
  1.446696e-07, 6.002873e-08, 4.166937e-08, 2.344516e-10, 3.959362e-08, 
    0.001794746, 0.02258612, 0.006489732, 0.1092729, 0.0008022526, 
    0.0003803015, 0.001850667, 0.0001549071, 9.032431e-06, 2.145473e-05, 
    1.323346e-05, 0.0004961777, 0.007605376, 0.0845972, 0.2033971, 
    0.01169694, 0.05026156, 0.0001479447, -0.002140018, 0.0001795015, 
    0.001672076, 0.01343279, 0.04804289, 1.224542e-07,
  4.582824e-07, -6.372488e-08, 0.00188747, -3.523749e-07, 2.445274e-08, 
    -6.109302e-10, -0.002177437, 0.3146548, 0.2910803, 0.02303137, 0.1182993, 
    0.01500872, 0.009776256, 0.0001428798, 0.000205568, 0.0001779457, 
    0.006834011, 0.03550488, 0.06967308, 0.1828368, 1.158911e-06, 
    0.000547717, 0.003656767, 0.0001363191, 0.002603912, 0.003545587, 
    0.0005514267, 0.03974522, 0.006021539,
  -0.0006274686, -4.504906e-05, 0.000602383, 0.1764154, -3.608215e-05, 
    2.366978e-08, 0.002760394, 5.275979e-07, -4.374327e-05, 0.01084726, 
    0.2135888, 0.1684307, 0.502865, 0.6494609, 0.593051, 0.2768794, 
    0.1857406, 0.1944892, 0.1861219, 0.002222847, 1.115744e-06, 2.275607e-05, 
    0.05900783, 0.2288266, 0.09247181, 0.06286318, 0.01457696, 0.05816987, 
    0.07038491,
  0.09452061, 0.01802212, 0.02782783, 0.008306365, 0.0007718506, 0.00420839, 
    0.003033729, 0.08589595, 0.06413515, 0.044914, 0.04901785, 0.1131469, 
    0.6745132, 0.5330821, 0.7329865, 0.5698771, 0.5504106, 0.3468291, 
    0.2541621, 0.09014024, 0.01456472, 0.008521781, 0.04353098, 0.1147494, 
    0.122897, 0.4699104, 0.3511157, 0.4561478, 0.4017934,
  0.1410323, 0.1268056, 0.05517234, 0.01002346, 0.009530043, 0.01026633, 
    0.05093365, 0.096348, 0.01101775, 0.05402579, 0.1397086, 0.3090389, 
    0.4679868, 0.3493474, 0.4590001, 0.6817364, 0.1980792, 0.3001798, 
    0.1924937, 0.0579862, 0.03894854, 0.1074325, 0.2676236, 0.1435528, 
    0.3328658, 0.1875371, 0.29026, 0.2568581, 0.2189206,
  0.564106, 0.3468174, 0.1482068, 0.225695, 0.3394805, 0.2948329, 0.2707237, 
    0.149493, 0.04672392, 0.1980128, 0.1566073, 0.2342812, 0.147704, 
    0.2934976, 0.3923379, 0.3699422, 0.2418933, 0.3711045, 0.3280913, 
    0.2970388, 0.3233047, 0.3256559, 0.1636762, 0.1864112, 0.4436279, 
    0.2903619, 0.1742227, 0.3245826, 0.6323336,
  0.4850056, 0.4129018, 0.478561, 0.5374393, 0.5624758, 0.5458484, 0.5676073, 
    0.4757782, 0.4825101, 0.49969, 0.5369585, 0.6503433, 0.6841354, 
    0.6073442, 0.5765366, 0.5598023, 0.5898811, 0.5572487, 0.4977491, 
    0.4855828, 0.5802202, 0.454467, 0.129184, 0.2349582, 0.2525159, 
    0.1765293, 0.1922513, 0.4263946, 0.3849387,
  0.01526833, 0.01406171, 0.01285508, 0.01164845, 0.01044183, 0.0092352, 
    0.008028573, 0.003112674, 0.004187748, 0.005262822, 0.006337896, 
    0.007412971, 0.008488045, 0.009563119, 0.01051431, 0.0117378, 0.01296128, 
    0.01418477, 0.01540825, 0.01663174, 0.01785522, 0.01321806, 0.01212613, 
    0.0110342, 0.009942266, 0.008850333, 0.007758401, 0.006666468, 0.01623364,
  0.06677447, 0.06787933, 0.0173575, 0.01943078, 0.04620567, 0.02093542, 
    0.02537923, 0.05028959, 0.01181858, 0.007412223, 0.01559533, 0.06594155, 
    0.1167285, 0.01219562, 0.2407819, 0.3072168, 0.1894041, 0.2208325, 
    0.2059418, 0.2813375, 0.5249989, 0.5837263, 0.06853685, 0.04621614, 
    0.3031895, 0.4413087, 0.1561419, 0.05352951, 0.06916965,
  0.1812392, 0.158418, 0.1747584, 0.04264985, 0.02207367, 0.07156203, 
    0.003930942, 0.08609995, 0.1955622, 0.1661914, 0.2254488, 0.2004969, 
    0.07751093, 0.1362744, 0.3788669, 0.396354, 0.3706061, 0.3466962, 
    0.2614997, 0.2761045, 0.2864866, 0.321546, 0.3339368, 0.4797568, 
    0.06628794, 0.2985058, 0.3477225, 0.4890465, 0.338562,
  0.2988267, 0.2668107, 0.1338565, 0.1321964, 0.1056453, 0.1153379, 
    0.1962769, 0.2028276, 0.1254189, 0.09197925, 0.1807782, 0.1999684, 
    0.1741772, 0.1782386, 0.08213787, 0.1322847, 0.1773375, 0.2547836, 
    0.1858215, 0.1244698, 0.1393783, 0.1281643, 0.1285977, 0.2064318, 
    0.2376469, 0.4229119, 0.3917542, 0.4873369, 0.3979493,
  0.2066316, 0.2159642, 0.2459358, 0.2607522, 0.3132561, 0.2024707, 
    0.1265039, 0.05773469, 0.1078831, 0.1290519, 0.08853227, 0.06452905, 
    0.06178242, 0.02979719, 0.0321389, 0.0520305, 0.03543006, 0.06650765, 
    0.08857227, 0.09932669, 0.07557569, 0.08172154, 0.06146336, 0.1328204, 
    0.05929116, 0.1652865, 0.2119553, 0.1811784, 0.2391918,
  0.05504747, 0.01307051, 0.02210695, 0.02027103, 0.02024311, 0.02079626, 
    0.01232096, 0.01700278, 0.02691691, 0.01401614, 0.02362197, 0.005070991, 
    0.002074574, 0.01432124, 0.08925016, 0.01630593, 0.02590489, 0.07992509, 
    0.042945, 0.08417981, 0.06212853, 0.06856014, 0.03942013, 0.4658651, 
    0.01983483, 0.02549707, 0.05458238, 0.03969472, 0.034131,
  0.007853253, 0.002370907, 0.01524169, 0.002090935, 0.001720502, 
    0.002443014, 0.0039254, 0.003606022, 0.004217152, 0.0006509767, 
    -0.000135359, -3.570765e-05, 0.01938878, 0.002565125, 0.003720509, 
    0.008813673, 0.03308174, 0.01063627, 0.049539, 0.01093349, 0.004637254, 
    0.002460384, 0.008157451, 0.007634442, 0.02373758, 0.01428714, 
    0.006030383, 0.002939808, 0.003744578,
  0.01195962, 0.01385023, -9.118279e-06, 0.001859253, -0.001637633, 
    0.000502547, 0.0008005553, 0.007687861, 0.002680974, 0.0004422574, 
    -1.555545e-10, -2.705153e-06, 0.0005890247, 0.0102943, 0.005250502, 
    0.001193647, 0.003084831, 0.0009211275, 0.001155187, 8.730194e-05, 
    0.001061118, 0.002108805, 0.01476921, 0.01737374, 0.005104272, 
    0.03883436, 1.822549e-05, 0.001282612, 0.003220113,
  0.03627963, 0.04039166, 0.0007687969, 0.01376281, 3.984366e-05, 
    0.0008104832, 0.002304132, 0.001505326, 3.990295e-05, -0.000636706, 
    0.007352556, 0.0001109853, 0.02086418, 0.002012577, 0.001260744, 
    0.0003458872, 0.0005139756, 0.0001551589, 0.0001051806, 2.144395e-05, 
    0.000532279, 0.005446594, 0.03920673, 0.00263506, -2.912292e-06, 
    1.375048e-08, -0.0005013579, -3.577451e-06, 0.005460892,
  0.0125234, 0.04482412, 0.0008991595, 0.002867925, 7.301978e-05, 
    0.0005183042, 0.0007842759, 0.0003816663, 0.02301423, 0.08554646, 
    0.002409194, 0.001461742, 0.0005770823, 0.0003964727, 0.0007674192, 
    0.0003938203, 0.0002645569, 0.0001265148, 0.0003929389, 0.00019973, 
    0.0001841228, 0.017914, 0.07498595, 0.04461396, 0.03643906, 7.825563e-05, 
    3.93878e-05, 0.000174984, 0.002797695,
  0.008544073, 0.01462737, 0.0003735835, 0.1404911, -6.754573e-07, 
    7.646559e-06, 0.01744634, 1.083658e-05, -0.0002770678, 0.000277877, 
    2.00648e-05, 0.001947054, 0.001629194, 0.0004136024, 0.0009610803, 
    0.001717274, 0.002876024, 0.002881897, 0.01293298, 0.005802046, 
    0.009495152, 0.003137445, 0.1439755, 0.02712319, 3.61717e-05, 
    0.002841251, 0.005388966, 0.01219415, 0.03235703,
  1.41313e-07, 5.856698e-08, 4.076848e-08, -9.936861e-11, 3.894311e-08, 
    0.000766537, 0.005345596, 0.001855493, 0.0627906, 5.808123e-05, 
    0.0001571209, 0.0004253162, 6.92673e-05, 6.789853e-06, 1.306085e-05, 
    6.62751e-06, 0.0002933473, 0.003446375, 0.04743901, 0.1087493, 
    0.00555301, 0.03610016, 9.594543e-05, -0.001610257, 0.000102149, 
    0.0009465283, 0.007568378, 0.02568934, 1.196714e-07,
  4.503448e-07, -4.614503e-08, 0.002859742, -1.106416e-06, 2.350534e-08, 
    -5.616189e-10, -0.00236923, 0.2797909, 0.2588464, 0.01432315, 0.09523126, 
    0.01167229, 0.003438157, 7.849517e-05, 0.0001095444, 8.874367e-05, 
    0.004035821, 0.02112753, 0.04090783, 0.1197861, -2.877344e-06, 
    0.001146065, 0.002568084, 7.721694e-05, 0.001666142, 0.002421541, 
    0.0003334702, 0.02319975, 0.005669937,
  -0.0005920147, -5.178625e-05, 7.890502e-05, 0.1687139, -2.830939e-05, 
    2.303192e-08, 0.001485478, 5.160566e-07, -2.910436e-05, 0.007036031, 
    0.2043313, 0.2688566, 0.4560128, 0.629004, 0.4971142, 0.1778607, 
    0.1078891, 0.1516558, 0.1256683, 0.002135725, 1.064528e-06, 9.275943e-06, 
    0.03983757, 0.1682503, 0.05259111, 0.02461923, 0.005350448, 0.03516424, 
    0.06364521,
  0.06040238, 0.01213474, 0.01843243, 0.004572055, 0.0003496899, 0.00208611, 
    0.001290586, 0.08602288, 0.05405074, 0.04014672, 0.04366211, 0.09757269, 
    0.6146411, 0.5037696, 0.6432669, 0.4467222, 0.3632903, 0.2234817, 
    0.2025354, 0.0767806, 0.008444263, 0.004392619, 0.03383607, 0.09577776, 
    0.1191397, 0.4350183, 0.2881255, 0.3416326, 0.3149029,
  0.09731352, 0.1024018, 0.03614258, 0.006418859, 0.009912139, 0.01419965, 
    0.04067331, 0.07599058, 0.01046783, 0.04902865, 0.1349236, 0.2734333, 
    0.4584492, 0.2994792, 0.5148062, 0.5812787, 0.1722222, 0.2624623, 
    0.125572, 0.05032167, 0.03196347, 0.09928955, 0.3412441, 0.117151, 
    0.4103026, 0.1757605, 0.227824, 0.1966601, 0.139442,
  0.4841968, 0.3038802, 0.1244194, 0.2401953, 0.3471741, 0.3851778, 
    0.2208313, 0.1144587, 0.03874893, 0.1689823, 0.1239232, 0.2025056, 
    0.1324593, 0.3289906, 0.3729301, 0.3240189, 0.1995348, 0.3716137, 
    0.3645328, 0.357943, 0.2514188, 0.3406934, 0.132898, 0.1810737, 
    0.4131429, 0.25218, 0.1583688, 0.2962404, 0.5485451,
  0.4255754, 0.3448168, 0.4022624, 0.4864803, 0.4931755, 0.4691181, 0.539049, 
    0.4028753, 0.4329841, 0.492965, 0.4975249, 0.5844173, 0.6003786, 
    0.4994689, 0.4977238, 0.514726, 0.4757157, 0.4723196, 0.4313899, 
    0.4078559, 0.5145769, 0.3976443, 0.1067, 0.1886759, 0.2237862, 0.1692589, 
    0.1858351, 0.3762613, 0.3392276,
  0.007301806, 0.006589465, 0.005877124, 0.005164783, 0.004452442, 
    0.003740101, 0.00302776, -0.0001993982, 0.0007906981, 0.001780794, 
    0.002770891, 0.003760987, 0.004751083, 0.00574118, 0.002664645, 
    0.004601967, 0.006539289, 0.008476611, 0.01041393, 0.01235125, 
    0.01428858, 0.02062868, 0.01841361, 0.01619853, 0.01398345, 0.01176837, 
    0.009553296, 0.007338218, 0.007871678,
  0.05158073, 0.04500922, 0.004680179, 0.01009208, 0.05184742, 0.02083061, 
    0.04317346, 0.02783657, 0.00944898, 0.007763642, 0.009922258, 0.05485279, 
    0.09640738, 0.006391765, 0.2912247, 0.246132, 0.1620731, 0.2193674, 
    0.1869417, 0.2756042, 0.5581102, 0.5909317, 0.05408606, 0.03817494, 
    0.2737066, 0.441405, 0.1329037, 0.03115784, 0.05294662,
  0.1519927, 0.1289391, 0.1335251, 0.03628453, 0.01608553, 0.06662814, 
    0.003928299, 0.06121745, 0.1414287, 0.1673863, 0.214429, 0.1668365, 
    0.05956238, 0.1087744, 0.3401344, 0.3679282, 0.3184523, 0.2978626, 
    0.219438, 0.2545007, 0.2680943, 0.2863398, 0.3129737, 0.464628, 0.051253, 
    0.3210358, 0.2868886, 0.3978671, 0.272347,
  0.2529148, 0.2336919, 0.1103052, 0.1065153, 0.08483194, 0.09355507, 
    0.1834408, 0.1790807, 0.09135379, 0.07761973, 0.1492888, 0.1703673, 
    0.1412501, 0.1465999, 0.06711388, 0.1070486, 0.1462146, 0.2102991, 
    0.1490897, 0.09790044, 0.1109086, 0.1029005, 0.09892856, 0.1682205, 
    0.2088782, 0.4121154, 0.3602477, 0.4502492, 0.3466206,
  0.1753377, 0.1746063, 0.2082091, 0.2276252, 0.2628733, 0.1695005, 
    0.1040292, 0.04349551, 0.08533756, 0.09645341, 0.06398246, 0.04604333, 
    0.0401755, 0.01942388, 0.01991959, 0.03604907, 0.02334775, 0.03874798, 
    0.06309018, 0.06998668, 0.05329138, 0.0598235, 0.04415398, 0.1321623, 
    0.03733394, 0.1310166, 0.1716798, 0.1470147, 0.200378,
  0.04044852, 0.008298518, 0.01777443, 0.0118882, 0.01341169, 0.01286342, 
    0.007326629, 0.01032017, 0.01760624, 0.008762678, 0.01451953, 
    0.003277812, 0.001643335, 0.008646008, 0.07416151, 0.01073637, 
    0.01302938, 0.05921159, 0.0281323, 0.05992584, 0.03982181, 0.04702172, 
    0.02244586, 0.4291695, 0.01171576, 0.01655655, 0.03753416, 0.02465782, 
    0.0195884,
  0.005932534, 0.00167635, 0.01125967, 0.001514389, 0.001252051, 0.002002005, 
    0.003212505, 0.002979581, 0.002456087, 0.0005147787, 0.0002751502, 
    -2.82963e-05, 0.01815999, 0.001191842, 0.002108373, 0.005251199, 
    0.02188817, 0.005824946, 0.03150332, 0.00558211, 0.002718287, 
    0.001431121, 0.00573822, 0.005158748, 0.02005724, 0.00677101, 
    0.003288096, 0.0017741, 0.002677485,
  0.009064477, 0.01089688, -1.202744e-05, 0.00137643, -0.001533171, 
    0.0003194922, 0.0005532496, 0.004084882, 0.001901606, 0.0003501388, 
    -1.28406e-10, -1.350882e-06, 0.0004469695, 0.005070751, 0.002910489, 
    0.0008682965, 0.00182177, 0.0006929421, 0.0005996515, 6.078636e-05, 
    0.0007114864, 0.001487558, 0.01078089, 0.01387605, 0.004751025, 
    0.03257624, 1.391375e-05, 0.0008396239, 0.002423778,
  0.027124, 0.0262618, 0.0004187788, 0.00793237, 2.334531e-05, 0.0005286753, 
    0.001147284, 0.0006945761, 2.988063e-05, -0.0004673136, 0.004148235, 
    8.386106e-05, 0.01011271, 0.0007238845, 0.0005183396, 0.0002141945, 
    0.000293512, 0.0001167149, 7.950114e-05, 1.5237e-05, 0.0003987657, 
    0.004013161, 0.02951471, 0.008949095, -1.063434e-06, 1.248205e-08, 
    -0.0003020743, -3.255571e-06, 0.004108042,
  0.009152206, 0.05561602, 0.001004544, 0.001431444, 4.579874e-05, 
    0.0003815625, 0.0005647694, 0.0002812726, 0.01839539, 0.08957382, 
    0.001590371, 0.0008624283, 0.0003716322, 0.0002140953, 0.0004682275, 
    0.0002485169, 0.0001947307, 9.186214e-05, 0.0002805199, 0.000135134, 
    0.0001178073, 0.01231723, 0.0556647, 0.04446673, 0.03009915, 
    5.724787e-05, 2.758111e-05, 0.0001266583, 0.001981516,
  0.005812005, 0.007116769, 0.0001522732, 0.1161918, -3.711244e-07, 
    4.79501e-06, 0.01045248, 7.157124e-06, -0.0001703752, 0.0001967781, 
    1.636068e-05, 0.001390557, 0.001015371, 0.0002775355, 0.0004034846, 
    0.0008144737, 0.001740563, 0.001562563, 0.006503909, 0.002658331, 
    0.004195514, 0.001369442, 0.1220829, 0.03148673, 2.902157e-05, 
    0.001287672, 0.002572183, 0.006335869, 0.01758985,
  1.357788e-07, 5.732783e-08, 4.009624e-08, -1.715439e-10, 3.796318e-08, 
    0.0004338358, 0.003264035, 0.0004385923, 0.03722546, -2.00851e-05, 
    9.385769e-05, 0.0002240618, 4.564009e-05, 5.664925e-06, 9.756909e-06, 
    4.448149e-06, 0.0002137459, 0.001812053, 0.02943499, 0.06741379, 
    0.003468408, 0.02673478, 7.071713e-05, -0.001299047, 7.112812e-05, 
    0.0006453972, 0.005098443, 0.01613803, 1.183398e-07,
  4.447035e-07, -1.059134e-07, 0.001512766, -7.86425e-07, 2.321858e-08, 
    -5.338973e-10, -0.002203383, 0.2524789, 0.2341042, 0.009701973, 
    0.06139953, 0.007585925, 0.001860036, 5.111613e-05, 7.093271e-05, 
    5.820319e-05, 0.002793437, 0.01507534, 0.02804185, 0.09045304, 
    -2.050106e-06, 0.009179479, 0.004916001, 5.321756e-05, 0.001217954, 
    0.001845936, 0.0002380185, 0.01613617, 0.004738485,
  -0.0005277481, -5.637774e-05, -8.881655e-05, 0.1533505, -2.332664e-05, 
    2.367042e-08, 0.0008706359, 5.073044e-07, -2.067402e-05, 0.004469397, 
    0.1869761, 0.2548399, 0.3750954, 0.5885293, 0.3841216, 0.1186306, 
    0.06303149, 0.09501154, 0.08345018, 0.002058067, 9.611608e-07, 
    8.392659e-05, 0.02209953, 0.1143285, 0.02754658, 0.01144632, 0.002949264, 
    0.02594968, 0.04968501,
  0.04146407, 0.008778753, 0.01340348, 0.00287809, 0.0002042777, 0.001205211, 
    0.0006867717, 0.08066388, 0.04513579, 0.03382052, 0.04747418, 0.08456401, 
    0.5028737, 0.4287893, 0.5470661, 0.3229718, 0.2570368, 0.1411711, 
    0.1331078, 0.06745587, 0.00566555, 0.002739939, 0.02860044, 0.07569589, 
    0.1225563, 0.3977433, 0.2212357, 0.2543198, 0.2154174,
  0.05866003, 0.08641016, 0.02485221, 0.004417872, 0.01316616, 0.01937711, 
    0.03629835, 0.0599131, 0.01242234, 0.05088361, 0.1306782, 0.2457418, 
    0.4347366, 0.2478078, 0.4789941, 0.4284888, 0.1528166, 0.2342352, 
    0.0843948, 0.04373321, 0.02860577, 0.09571487, 0.3572923, 0.09507848, 
    0.3985349, 0.1675981, 0.1803598, 0.1445638, 0.09158504,
  0.3826483, 0.2414675, 0.1111231, 0.2682442, 0.3284228, 0.4519345, 
    0.1811569, 0.08979918, 0.03197144, 0.1404792, 0.09801087, 0.1785798, 
    0.1122127, 0.368901, 0.3751721, 0.271846, 0.1675269, 0.3537527, 
    0.3597673, 0.4942658, 0.1913673, 0.3470334, 0.1047874, 0.162408, 
    0.3690342, 0.2257134, 0.1437556, 0.2600336, 0.4422283,
  0.3407692, 0.3047169, 0.346143, 0.4237717, 0.4120035, 0.409349, 0.4619511, 
    0.3341182, 0.3948003, 0.4015776, 0.4129427, 0.4860184, 0.473844, 
    0.3996458, 0.4045362, 0.4127926, 0.3917949, 0.3848046, 0.3494167, 
    0.3434191, 0.4269061, 0.3543073, 0.09380339, 0.1602956, 0.1937211, 
    0.1626247, 0.1748837, 0.3448317, 0.2910016,
  0.006030517, 0.005746993, 0.005463469, 0.005179945, 0.004896421, 
    0.004612897, 0.004329373, 0.0008422141, 0.001424568, 0.002006922, 
    0.002589277, 0.003171631, 0.003753985, 0.004336339, 0.004055295, 
    0.005693711, 0.007332128, 0.008970545, 0.01060896, 0.01224738, 0.0138858, 
    0.01612719, 0.01418995, 0.0122527, 0.01031545, 0.008378207, 0.006440959, 
    0.004503713, 0.006257336,
  0.01315673, 0.01630084, 0.004122925, 0.0121777, 0.02028319, 0.1052789, 
    0.06342374, 0.02748396, 0.002084313, 0.007978473, 0.01005963, 0.04727972, 
    0.09228095, 0.004419802, 0.2673807, 0.1549338, 0.1390872, 0.254449, 
    0.186403, 0.2783056, 0.5237392, 0.5448208, 0.05710712, 0.04495587, 
    0.2508533, 0.425148, 0.1430862, 0.02895029, 0.04292064,
  0.1538011, 0.1248109, 0.12542, 0.03306207, 0.01553982, 0.0647819, 
    0.003854091, 0.05648961, 0.1241504, 0.1556782, 0.2145611, 0.1601202, 
    0.05539513, 0.1013601, 0.30837, 0.3349928, 0.3112874, 0.2749675, 
    0.1995324, 0.2442417, 0.2606224, 0.2814255, 0.2984984, 0.4597895, 
    0.04941702, 0.3194396, 0.2720214, 0.3577707, 0.2518033,
  0.2323648, 0.213414, 0.09942394, 0.09359533, 0.07513611, 0.08209456, 
    0.1951218, 0.1677753, 0.07702138, 0.06689075, 0.1281411, 0.1497625, 
    0.1220068, 0.1281664, 0.05880786, 0.09210838, 0.1263536, 0.1809399, 
    0.1294241, 0.08223215, 0.09238556, 0.08717739, 0.0805877, 0.1431282, 
    0.1951904, 0.400959, 0.3417438, 0.4245615, 0.3117474,
  0.1505049, 0.1476961, 0.1758342, 0.1912211, 0.2220207, 0.1460175, 
    0.09158278, 0.03764451, 0.07354876, 0.0825175, 0.05341945, 0.03792933, 
    0.02966522, 0.01495722, 0.01455471, 0.02805818, 0.01749073, 0.02539748, 
    0.04946633, 0.05378533, 0.0420731, 0.04684505, 0.03587883, 0.1846058, 
    0.02909709, 0.1034039, 0.1424025, 0.1260125, 0.1744389,
  0.03234378, 0.006596302, 0.01368224, 0.008623922, 0.01053948, 0.009255153, 
    0.005472914, 0.007582396, 0.01332956, 0.006260622, 0.01073526, 
    0.002729488, 0.001408928, 0.005861625, 0.08326817, 0.007897099, 
    0.006777454, 0.04537721, 0.02121783, 0.04598406, 0.02775312, 0.03268286, 
    0.01502821, 0.4206078, 0.007353112, 0.01237004, 0.0287776, 0.01768154, 
    0.01398674,
  0.004985985, 0.001373237, 0.01204993, 0.00124345, 0.001045684, 0.001758834, 
    0.002815539, 0.002638672, 0.001890751, 0.0003834508, 0.0008092728, 
    -1.91528e-05, 0.03205072, 0.0007671913, 0.001475256, 0.003582589, 
    0.01346074, 0.004017139, 0.02172799, 0.003540233, 0.002143309, 
    0.001105925, 0.004597149, 0.004157795, 0.02788489, 0.004662691, 
    0.002235123, 0.00134368, 0.002193173,
  0.007632053, 0.009635728, -2.102565e-05, 0.00113597, -0.001555847, 
    0.0002497855, 0.0004536623, 0.002950194, 0.001548247, 0.0003040503, 
    -1.082984e-10, -6.893479e-07, 0.0003797626, 0.00329695, 0.001836504, 
    0.0007123187, 0.001364288, 0.0005731905, 0.0004297128, 4.953667e-05, 
    0.0005694975, 0.001218451, 0.008861399, 0.01180895, 0.009534176, 
    0.03093634, 1.199802e-05, 0.0006547166, 0.002033854,
  0.0225358, 0.02024436, 0.0002982775, 0.009913038, 1.846334e-05, 
    0.0004181925, 0.0007729676, 0.0004679791, 2.553979e-05, -0.0004083033, 
    0.002978405, 7.226398e-05, 0.006821919, 0.0004856005, 0.0003419002, 
    0.00016284, 0.0002226152, 9.809399e-05, 6.687365e-05, 1.258468e-05, 
    0.0003378107, 0.003345018, 0.02463944, 0.02065998, -5.72796e-07, 
    1.355658e-08, -0.0002537902, -2.965327e-06, 0.003444923,
  0.007495322, 0.1000469, 0.007841782, 0.00104704, 3.618715e-05, 
    0.0003167362, 0.0004546724, 0.0002318723, 0.02204502, 0.09222147, 
    0.001221654, 0.0006486317, 0.0002949859, 0.000147232, 0.0003480147, 
    0.000209634, 0.0001619161, 7.591108e-05, 0.0002310913, 0.0001089283, 
    9.204829e-05, 0.009698396, 0.04506382, 0.07492201, 0.05333252, 
    4.784439e-05, 2.286548e-05, 0.0001045895, 0.00159349,
  0.0445649, 0.004807863, 6.856181e-06, 0.1064679, -2.388912e-07, 
    3.718495e-06, 0.02026708, 5.849749e-06, -0.002230432, 0.0001650783, 
    1.463534e-05, 0.001123334, 0.000759629, 0.0002190363, 0.0002546156, 
    0.0005526759, 0.001067943, 0.001129223, 0.003836085, 0.001714139, 
    0.002680828, 0.0009206738, 0.1745558, 0.04901984, 2.473296e-05, 
    0.0007626578, 0.001445705, 0.00402355, 0.04730679,
  1.346646e-07, 5.68587e-08, 3.956616e-08, -1.842919e-10, 3.787334e-08, 
    0.0003275725, 0.001576493, 0.0001236474, 0.08358395, -0.0006840831, 
    7.13686e-05, 0.0001659536, 3.698286e-05, 5.049866e-06, 8.380248e-06, 
    3.618789e-06, 0.0001805315, 0.001339206, 0.02034061, 0.04865915, 
    0.002594612, 0.02294326, 5.78114e-05, -0.00174514, 5.893843e-05, 
    0.0005271143, 0.004058548, 0.01262403, 1.184646e-07,
  4.40731e-07, -5.543109e-07, 0.0009552256, -5.528197e-07, 2.371748e-08, 
    -5.195758e-10, -0.002164425, 0.2401588, 0.2474296, 0.007061253, 
    0.04557889, 0.003802082, 0.001308369, 4.107733e-05, 5.459756e-05, 
    4.690782e-05, 0.002230953, 0.01214405, 0.02218018, 0.07570424, 
    -1.393215e-06, 0.051671, 0.0561174, 4.282341e-05, 0.0009923133, 
    0.001541795, 0.000198877, 0.01287513, 0.003978719,
  -0.0005443579, -5.289087e-05, -0.0003959713, 0.1571751, -2.136776e-05, 
    2.42575e-08, 0.0006228199, 4.925461e-07, -1.662668e-05, 0.002875646, 
    0.1932767, 0.2112363, 0.2892685, 0.4549776, 0.2749645, 0.08174684, 
    0.04345909, 0.06729043, 0.0579255, 0.001455344, 5.679489e-07, 
    0.0008369734, 0.03049195, 0.0840178, 0.0176721, 0.007536475, 0.002148522, 
    0.01783584, 0.04139098,
  0.03426034, 0.0137964, 0.01128204, 0.002613914, 0.0001410874, 0.0008700647, 
    0.000520778, 0.07692616, 0.05991899, 0.04175999, 0.1143258, 0.1012701, 
    0.4017895, 0.3646603, 0.441189, 0.2349328, 0.1929144, 0.09998474, 
    0.09307356, 0.06653016, 0.008074711, 0.002110883, 0.0345467, 0.09693899, 
    0.1190683, 0.3520847, 0.1698614, 0.1944967, 0.1583402,
  0.03687258, 0.08766023, 0.02796907, 0.0105904, 0.04805257, 0.03849158, 
    0.05155611, 0.08382114, 0.04211374, 0.07674708, 0.1504181, 0.2655444, 
    0.4291697, 0.2207209, 0.4140976, 0.3147385, 0.1580278, 0.2246396, 
    0.08376734, 0.05328149, 0.04618392, 0.1024559, 0.3185391, 0.09255984, 
    0.3414399, 0.1561779, 0.1417878, 0.107942, 0.06283557,
  0.297838, 0.1854385, 0.123129, 0.2629025, 0.2943343, 0.5262829, 0.1641528, 
    0.08501172, 0.03122984, 0.1293643, 0.09547542, 0.178781, 0.1130918, 
    0.3772413, 0.386584, 0.2521979, 0.1575834, 0.340663, 0.3242236, 
    0.5281329, 0.1548383, 0.34569, 0.08618345, 0.1466389, 0.3284837, 
    0.2094824, 0.1415147, 0.2213221, 0.3522151,
  0.2869428, 0.2705804, 0.2969197, 0.3672748, 0.3529845, 0.3619412, 
    0.4123618, 0.2860667, 0.3510319, 0.3281116, 0.3459038, 0.4100188, 
    0.3961231, 0.3305266, 0.3288443, 0.3448489, 0.3426966, 0.3395096, 
    0.3019188, 0.2870085, 0.377228, 0.3272761, 0.0851128, 0.1424526, 
    0.1759765, 0.1616799, 0.1653738, 0.322729, 0.250118,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3.304549e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 7.397156e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -7.776899e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.001311019, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -9.953089e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0.003724629, 0, 0, 0, 2.74305e-05, 0, 0, 0, 5.257033e-06, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 4.142155e-05, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0001409479, 0.0002028111, 0, 
    0.001499262, 0.0001671886, 0.0002866296, -1.456187e-05, 0, 0, 0, 0, 
    0.004406724, 0, 0, 0, 0, -3.162182e-06, 0,
  0, 0, 0, 0, 0, 0, -0.0001792046, 0, 0, -2.223314e-05, -4.948355e-06, 
    -1.990618e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -4.299484e-05, 0, 0.000316019, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -3.765766e-06, 2.326148e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0.005536182, 0, 0, -3.652606e-05, 0.002081734, 0, 
    4.624165e-05, 0.0012426, 0.0004588696, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0001284299, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0003264929, 0.0005709807, 1.145682e-05, 
    0.002133867, 0.001307737, 0.0004818797, 0.001110239, 0, 0.0007508649, 
    -3.668315e-06, -8.351467e-07, 0.007701748, 6.724415e-05, -3.178334e-07, 
    0, 0.0004436756, 7.730328e-06, 0.004361155,
  0, 0, 0, 0, 0, 0, 0.0005996231, -3.780832e-07, 0, -0.0001708506, 
    -7.505884e-05, -1.919966e-05, 0, -1.274635e-05, 0, 0, 0, 0, 0, 0, 0, 
    0.0002550754, 0, -1.288199e-05, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -8.732542e-06, -4.455276e-05, 0.001082908, 0, 
    0.0007340096, -7.313337e-06, 0.0004886498, 0.00259362, -4.380831e-06, 0, 
    0, 0, 0, 0, 0, 0, 0.0001929127, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -1.538317e-06, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -0.0001481485, 0.0003187897, -1.346809e-05, 0, 0, 0, 0, 
    -1.72096e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0.007508911, 0, -5.577214e-06, -5.56094e-05, 0.005643562, 0, 
    9.860314e-05, 0.006746626, 0.001830018, -2.458648e-05, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.000129561, 0, 0, 0, 0, 0,
  -7.917817e-06, -1.227245e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0005300812, 
    0.0008827217, -4.822146e-05, 0.004057602, 0.001817226, 0.002040703, 
    0.005593573, 0.005355057, 0.002424941, -9.199588e-05, 0.0001356112, 
    0.01207872, 0.000114598, -1.650468e-06, 0, 0.002817814, 0.0001092851, 
    0.008052548,
  0, 0, 0, 0, 0, 0, 0.002813574, -1.995693e-05, -4.497698e-05, 0.0003167441, 
    -0.0001448739, -0.0001683019, 6.585693e-05, 0.0001808968, 0, 0, 0, 0, 0, 
    0, -1.315078e-05, 0.0005250791, 0, -7.945183e-05, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -5.347989e-05, -0.0002024675, 0.003692323, 0, 0.01054096, 
    -6.25521e-05, 0.001740642, 0.004631435, 0.0006853461, 0, 0, 0, 0, 0, 0, 
    0, 0.001567923, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.462447e-05, -3.225035e-05, 
    -4.525334e-10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0003132753, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0.002107496, 0.0004470313, 0.0005177587, 0, 0, 0, 0, 
    -2.067763e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0.009483919, 0, -3.216952e-05, -7.535047e-05, 0.01109623, 0, 
    0.001478271, 0.01801215, 0.005368839, -3.302236e-05, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.0001680588, 0, 0, 0, 0, 0,
  0.001336893, 0.002384237, -4.212142e-06, -2.480496e-06, 0, 0, 0, 
    0.0001171919, 0, 0, 0, -0.0004924404, 0.002834129, 0.0006062714, 
    0.007454579, 0.004004705, 0.005317218, 0.01513781, 0.01285087, 
    0.01057123, 0.0004697243, 0.0007077801, 0.01732193, 0.003504835, 
    -3.954097e-06, -2.900555e-05, 0.006211355, 0.000397121, 0.01267898,
  0, 0, 0, 0, 0, 0, 0.005121784, -0.0001571707, -7.831419e-05, 0.002702977, 
    0.0001819023, -0.000397217, 0.0005743127, 0.0006341203, 0, 0, 0, 0, 0, 0, 
    -6.434934e-05, 0.001821695, 0, 0.0001732864, -2.967143e-11, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0.0001243431, 0.0008893317, 0.006925838, 0, 0.02456839, 
    0.001797317, 0.006305302, 0.00986966, 0.0008490715, 0, 0, 0, 0, 0, 0, 
    -4.185141e-05, 0.002589069, -6.173724e-05, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001859774, 0.002532947, 6.99085e-05, 
    -4.951944e-06, -4.18717e-05, 0, 0, 0, 0, 0, 0, -9.662086e-06, 
    0.0006374117, -2.973677e-05, 0.004732923, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.023473e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.000278982, -2.580431e-05, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -4.992336e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 8.142883e-05, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -5.06416e-08, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.00147794, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0.009570234, 0.002069654, 0.006799331, 0, 0, 0, 0, 
    0.001451626, -5.074075e-06, -1.666716e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0,
  0, -6.262029e-06, 0, 0, 0, 0.01454605, 0, -8.432538e-05, -0.0002534013, 
    0.01572421, 2.581624e-05, 0.006926895, 0.03216372, 0.007613408, 
    0.001196315, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002270795, 0, 0, 0, 0, 0,
  0.004674089, 0.006932403, 9.001642e-05, -3.472694e-05, 0, -1.188203e-05, 0, 
    0.0007171815, 0, 0, 0, 0.005231637, 0.009201746, 0.004367336, 0.01206532, 
    0.008322548, 0.01307393, 0.02874839, 0.0201867, 0.02565956, 0.002767293, 
    0.004653561, 0.02453566, 0.007830152, -1.368633e-05, -4.096375e-05, 
    0.01070916, 0.003844445, 0.02346979,
  0, 0, 0, 0, 0, 0.0003727683, 0.02922405, -0.0001640122, 0.0002605611, 
    0.005843909, 0.004652539, 8.427067e-05, 0.001872297, 0.004797274, 
    9.764454e-05, 0, 0, 0, -1.468673e-08, 0, -0.0003448326, 0.01091358, 
    -5.948958e-06, 0.0007882839, -5.61284e-06, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0.001959874, 0.001852271, 0.00873722, 0.0002395745, 
    0.03731093, 0.004519033, 0.01224527, 0.01393964, 0.005299149, 0, 0, 0, 0, 
    0, 0, 0.001676562, 0.005134747, 0.0002452342, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0.002213508, -1.12519e-05, 0.00823541, 0.013747, 
    0.004443977, -0.0001829939, 0.0001091054, 0.001220764, 0.000170672, 0, 0, 
    0, 0, 9.598994e-06, 0.001291662, -5.226551e-05, 0.008579751, 0, 
    8.492551e-05, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, -2.739777e-05, 0.0001963397, -8.405982e-05, 
    0.001158407, 0, -0.0001272488, -9.33483e-05, 0, 0, 0, 0, 0, 
    -4.400938e-06, 0.002969042, 0.001718197, 0.004095128, -0.0001133639, 
    0.00177, -3.841392e-09, 0, 0.001245724,
  0, -6.644782e-05, 0, 0, 0, -2.061698e-05, 0, 0, 0, -1.878505e-05, 
    -4.912081e-06, -4.930709e-05, 0, 0, 0, 0.0002016717, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, -2.464759e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.001146291, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0005717142, 0, 
    -3.484401e-06, 4.572875e-05, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -5.252848e-05, 0.002545451, 
    0.0001248476, -6.557962e-05, 0.001027197, 0, 0, 0, 0, -1.241109e-05, 
    0.003161028, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.34073e-06, -9.612618e-08, 
    0.01033895, 0, 0, 0, 0, 0, -4.697615e-07, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0.01980515, 0.005463761, 0.009142965, 0, 0, 8.784213e-05, 
    0.0001310355, 0.005184997, 0.0003053266, -3.902416e-05, 0, 0, 0, 0, 0, 0, 
    0, 0, -1.369034e-08, 0, 0, 0, 0,
  0, 6.180784e-06, 0, 0, 0, 0.02063347, -3.103803e-06, -9.242928e-05, 
    0.000836546, 0.02520403, 1.019498e-06, 0.01229699, 0.04952792, 
    0.01321484, 0.002904749, -3.309563e-06, 0, 0, 0, 0, 0, -2.797373e-05, 
    -6.090294e-08, 0.0005202969, 0, 0, 0, 0, 0,
  0.008289454, 0.0110069, 2.759479e-05, 0.001739517, 0, 6.559515e-05, 
    0.000200859, 0.002618325, -3.873834e-05, -8.812211e-06, 4.306621e-07, 
    0.01031664, 0.02208038, 0.0100124, 0.0146865, 0.02026351, 0.02702035, 
    0.05273103, 0.02682408, 0.04287529, 0.01183497, 0.01771812, 0.03485927, 
    0.01208379, 0.0001224194, -2.517798e-07, 0.01844166, 0.01372994, 
    0.03243214,
  0, 0, 0, -9.92722e-10, -8.692593e-07, 0.001398805, 0.0724159, 0.002858388, 
    0.001156392, 0.02157481, 0.01292486, 0.005634544, 0.007044317, 
    0.02324247, 0.0004706559, 0, 0, 0, -4.772965e-05, 0, -3.167496e-05, 
    0.02113503, 0.0004294256, 0.001411471, -3.653967e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0.01358942, 0.004002441, 0.01363089, 0.0008014104, 
    0.04239978, 0.009120496, 0.02922448, 0.02376681, 0.02376383, 0.000146351, 
    0, 0, 0, 0, -1.02503e-05, 0.002490466, 0.01605566, 0.006885165, 0, 0, 0, 
    0, 0,
  0, 0, 0, -1.343327e-10, 0, 0, -1.678351e-10, -2.467592e-07, 0.003318746, 
    2.434718e-05, 0.01512498, 0.02628683, 0.01148302, 0.001898528, 
    0.005976528, 0.004704235, 0.000103431, 0, 0, 0, 0, 2.587327e-05, 
    0.003802098, -4.084435e-05, 0.01508746, -5.09648e-06, 0.003915021, 
    -6.013477e-06, 0,
  -6.259682e-05, -1.415495e-05, 8.180382e-05, 0.0004066682, 0.001174048, 
    -3.261762e-05, 0, 0, -0.0002601964, 0.01145511, 0.008003554, 0.01054175, 
    -0.0001255473, 0.009389894, 0.003178949, -5.951984e-06, 0.0003647356, 0, 
    0, 0, 0.0005263283, 0.006682093, 0.002866116, 0.006788748, 0.001417548, 
    0.00315884, 0.0006679969, -3.51169e-07, 0.004293205,
  5.541941e-05, -0.0001263121, 0.003008289, 0, 0, -0.000168312, 
    -5.548661e-05, 0, 0, 0.0004192867, -4.782166e-05, 0.004536358, 
    -5.151101e-05, 0.0003426692, -4.518401e-05, 0.003009316, -0.0001575986, 
    0, 0, 0, 7.223123e-05, 4.494044e-05, -3.50832e-05, -2.327108e-06, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -5.028679e-09, 2.931763e-08, 0, 5.907725e-10, 
    0, 0, 0, 0, 0, 0, -3.591023e-06, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.898473e-09, 1.237189e-07, 
    4.14432e-07, -4.165202e-10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0.003844227, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002987092, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.00261012, 0,
  0, 0, -5.572049e-06, 0.0003995509, 0, -8.099038e-06, 0, 0, 0, 0, 0, 0, 0, 
    0, -3.768579e-05, 0, 0, 0, 0.00476088, 6.603153e-05, -3.034671e-05, 
    0.006966325, -2.941264e-07, 0, 0.001374895, 0.001638276, 0.0003729905, 
    0.0006544045, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.008073164, 0.01395371, 
    0.0122365, 0.004657384, 0.005940538, 0, 0, 0, 0, -8.973612e-05, 
    0.005451042, -9.094698e-06, 0, 0,
  0, 0, 0, 0, 0, 0, -3.360113e-06, 0, 0, 0, 0, 0, 0, 0, 0.00033436, 
    0.007359319, 0.02083879, 0.000298249, -1.767262e-08, 0, 0, 0, 
    -8.732157e-08, -1.813373e-09, 0, -1.018004e-05, 0, 0, 0,
  2.680633e-07, -2.280568e-09, 0, 0, 0, -6.866236e-06, 0.04248492, 
    0.01268951, 0.01328574, 0, 0.0001276861, 0.0003862284, 0.0009824735, 
    0.01060671, 0.0006219893, -6.373235e-05, 0, 0, 0, 1.306376e-07, 0, 
    -1.635645e-09, 2.090346e-08, 0, -2.6859e-05, 5.454172e-09, 0, 0, 0,
  -2.357044e-09, 0.001461975, 0.0001069484, 0, 0, 0.0397763, 0.0008985173, 
    0.004179223, 0.009909909, 0.04315565, 0.004765333, 0.02786676, 
    0.07600684, 0.02475824, 0.005063667, -2.419823e-05, 0, -1.300911e-07, 0, 
    -2.456395e-07, 0.0003739936, 0.0004182456, -2.242515e-05, 0.01231015, 
    -1.294105e-06, 0, -7.923767e-06, 0, 0,
  0.02135233, 0.01912989, 0.002261188, 0.005615908, 0, -1.471553e-05, 
    0.000466752, 0.01216478, 0.0006145011, 0.0001842776, 0.0003306283, 
    0.02400938, 0.04901005, 0.02544281, 0.02996717, 0.0519166, 0.05389896, 
    0.07647538, 0.04287825, 0.06664182, 0.03476495, 0.06535684, 0.0608172, 
    0.02425157, 0.002125872, 0.004546729, 0.02812391, 0.03209441, 0.04445796,
  0, -1.874642e-07, 0, 0.0002345633, 0.0004460297, 0.01045888, 0.1131899, 
    0.0796807, 0.02056959, 0.13424, 0.02851774, 0.02791097, 0.04669183, 
    0.06430186, 0.005214353, 0.0001357061, -3.380981e-09, 0, 0.001839814, 
    6.239612e-06, 0.006619763, 0.04793481, 0.001955726, 0.004407904, 
    0.0002301237, 0, 0, 0, 0,
  0, 0, 0, 0, -6.524264e-09, 4.396855e-09, 0.08259246, 0.009121002, 
    0.02375734, 0.01837235, 0.08228625, 0.01527679, 0.08733953, 0.05291534, 
    0.05193381, 0.006472963, -4.523436e-05, 0, 0, 0, 1.014326e-06, 
    0.01092432, 0.03750905, 0.01442527, -2.696887e-05, 0.00144685, 0, 0, 0,
  0, -7.086202e-06, 0, 3.142625e-07, -6.433844e-10, 0, -1.940673e-07, 
    -5.076038e-05, 0.005449301, 0.00278661, 0.02976443, 0.04575851, 
    0.01821931, 0.0109873, 0.02883829, 0.00685322, 0.005897025, 
    -2.293478e-05, 1.764445e-06, 0, -2.33696e-05, 0.002317676, 0.007111168, 
    0.004499816, 0.02227736, 0.003542014, 0.01303509, 0.002348113, 0,
  0.0004535955, -6.394247e-05, 0.005022265, 0.002414867, 0.005091988, 
    -4.731597e-05, 0, 0, 0.01351955, 0.0233358, 0.02124802, 0.0201611, 
    0.001739988, 0.04509094, 0.01122006, 2.987908e-05, 0.0007682983, 
    -3.523877e-06, 0.003251411, -2.62944e-05, 0.002504099, 0.01263889, 
    0.01213107, 0.0117402, 0.01525427, 0.01555066, 0.007070671, 9.587759e-05, 
    0.008830003,
  0.0009196003, 0.003610704, 0.006722202, 0, 0, 0.001310323, 0.0001003922, 0, 
    0, 0.004996229, 0.000833871, 0.02872721, 0.009794442, 0.00482068, 
    0.003757741, 0.009100131, 0.00715574, 0, 0, 0, 0.00220031, 0.0004896531, 
    0.00245683, -2.372447e-05, 0.0002302959, 0.0005379948, -4.53133e-05, 0, 0,
  0, 0, 0, 0, 0, 0, 0.002162455, 0, 0, 0, 9.336148e-09, 1.547096e-08, 
    -0.0001166451, -0.0001074879, 0, 0, 0, 0, 0, -8.662677e-05, 0.0008817705, 
    -1.728536e-05, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3.837988e-11, -1.655783e-09, 
    2.379938e-07, 2.559478e-07, 0, 0, 2.453433e-09, -1.439317e-10, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0.001131341, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, -3.002754e-05, 0.007838336, 0, 4.780838e-05, 0, 0, 0, 0, 0, 0, 0, 
    -9.281848e-06, 0, 0.003654681, 0, 0, 0, 0, 0, 0, -2.471161e-06, 
    0.0005585153, 0, 0, 0.003963839, 0,
  -1.759534e-05, 0, -1.085765e-05, 0.01180865, 0, 0.001385811, -2.308302e-05, 
    0, 0, 0, 0, 0, 0, 1.278087e-05, -0.0001176223, 0, 0, -7.603237e-05, 
    0.01112767, 0.001116808, 0.007069221, 0.008505846, 0.00221176, 0, 
    0.003143449, 0.005610232, 0.005131502, 0.006644465, -5.988514e-05,
  0, 0.0006208092, 0, 0, 0.007095178, -2.268293e-05, -2.535537e-08, 
    -1.706842e-09, 0, 0, 0, 0, 0, -9.32865e-11, 5.285583e-07, 0.02535327, 
    0.03879215, 0.04001778, 0.02091275, 0.008254429, 0.0008232347, 
    2.624112e-05, 0, 0.0005317514, -0.0001968321, 0.006653407, -0.0001066114, 
    -1.635043e-10, -1.469334e-05,
  3.491621e-07, -2.348227e-08, 0, 0, 1.053754e-08, 5.625227e-08, 
    2.541026e-05, 3.27451e-08, 9.606359e-08, 4.910433e-07, 8.665261e-08, 
    3.244603e-07, 9.815503e-07, -1.226558e-07, 0.002237148, 0.02031091, 
    0.03213, 0.006729029, 4.083345e-05, 6.500465e-06, 0, 0, 4.680188e-05, 
    1.407636e-05, 5.302121e-05, 0.0001194547, 2.525526e-07, -3.176194e-08, 0,
  4.196027e-05, 0.0007824645, 0, 0, 0, -1.811336e-05, 0.06693203, 0.02161211, 
    0.03386589, 0.004668963, 0.004172014, 0.04533813, 0.01197225, 0.02948149, 
    0.02229525, -2.587405e-05, -3.321124e-12, -1.095312e-09, 5.395279e-08, 
    0.0005218142, 0.0002054188, 1.092298e-07, -1.322425e-05, -1.999745e-05, 
    0.001182201, -5.282764e-05, 1.11094e-05, -1.605554e-06, 9.533804e-06,
  2.008484e-05, 0.01150605, 0.003619328, -3.554218e-06, 0, 0.06479231, 
    0.00140867, 0.03846778, 0.07732544, 0.09578491, 0.1349769, 0.1650334, 
    0.2309377, 0.08936402, 0.06482057, 0.002469472, -2.779443e-05, 
    -7.615253e-06, 6.326775e-05, 0.0008634938, 0.0008341963, 0.003656212, 
    0.005434915, 0.05006442, 0.00108868, -2.101804e-10, 0.0004289402, 
    0.0135436, -2.210466e-07,
  0.1085113, 0.0462448, 0.02106875, 0.01133608, -0.0003324538, 0.004075763, 
    0.05695664, 0.4376762, 0.3045285, 0.155822, 0.2278366, 0.1897102, 
    0.2451996, 0.1815838, 0.1801092, 0.2020406, 0.09989878, 0.1194179, 
    0.112225, 0.1265262, 0.1187095, 0.2770516, 0.1282605, 0.0848323, 
    0.0271461, 0.008566303, 0.04480879, 0.07848062, 0.06833235,
  -2.100613e-08, 5.404039e-05, 0.002149213, 0.01324818, 0.02266627, 
    0.1087798, 0.2650246, 0.2762249, 0.3419448, 0.3220634, 0.2538406, 
    0.152956, 0.3444712, 0.3137313, 0.09260428, 0.0002917164, -6.548918e-05, 
    -1.683771e-07, 0.01353745, 0.001449322, 0.04176468, 0.1700991, 
    0.08330962, 0.02951318, 0.005000202, 2.818439e-05, 1.536588e-06, 
    -1.099925e-05, -2.630571e-09,
  0, 0, -1.801047e-09, 6.197139e-09, 4.313172e-08, 5.296974e-06, 0.0958974, 
    0.02568438, 0.04696335, 0.1465935, 0.1728704, 0.1404321, 0.2224196, 
    0.1145518, 0.1574249, 0.01358107, 0.0003157331, 0.0005496058, 
    0.000255367, 0.000389851, -0.0004017521, 0.07610944, 0.1083692, 
    0.04065051, -1.700917e-05, 0.002293741, -1.598642e-07, -7.11769e-08, 0,
  1.64215e-07, -3.7922e-05, -3.515158e-08, 5.274786e-06, 3.393724e-07, 
    6.921226e-08, -2.379973e-06, 0.0007728606, 0.02900562, 0.02898898, 
    0.09907199, 0.1634849, 0.04459911, 0.04320022, 0.09335726, 0.02018435, 
    0.03195043, 0.0002494831, 4.52768e-05, -2.805962e-07, 0.001404786, 
    0.004136387, 0.01308151, 0.01251211, 0.04143108, 0.00412366, 0.02307442, 
    0.004835872, 1.015691e-06,
  0.004817833, 0.001466917, 0.0329572, 0.007557849, 0.008988601, 0.004439468, 
    0.0003818473, 5.707696e-06, 0.03269875, 0.04844164, 0.05521877, 
    0.03982623, 0.02304566, 0.09738136, 0.06594928, 0.01159832, 0.002730931, 
    0.0009636034, 0.00977392, 0.0002554241, 0.004707641, 0.0305669, 
    0.02139337, 0.01952155, 0.02357862, 0.03334093, 0.01736954, 0.004427945, 
    0.01242901,
  0.006248, 0.006602046, 0.0148462, 0, -2.319807e-06, 0.005102154, 
    0.005560953, 0, 0, 0.01822768, 0.009978306, 0.05445928, 0.01872464, 
    0.009715192, 0.01486216, 0.01525131, 0.01407491, -1.548117e-05, 0, 
    -1.703092e-06, 0.006878066, 0.002872576, 0.009712783, 0.002584942, 
    0.01546248, 0.007874371, 5.589144e-05, 0.0002820354, 0,
  0, 0, 0, 0, 0, 0, 0.007695911, -0.000144586, 0, 0.001865294, 0.004083153, 
    0.0004119349, 0.0008283443, 0.0007815849, 0, -1.398555e-05, 
    -3.648466e-06, 0, -7.179699e-06, -8.662677e-05, 0.008547327, 
    -0.0005427463, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.065335e-09, 4.453072e-08, 0.0003630721, 
    -0.0003529459, -1.910196e-08, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0.003387537, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, -4.322415e-06, 0.0008418779, 0.01770718, -8.101541e-06, 0.001713551, 
    0, -8.819572e-06, 0, 0, 0, 0, -2.382343e-05, 8.156036e-05, 0, 
    0.005449108, 1.383775e-05, 0, 0, 0, -5.587958e-06, 0, 0.0006037121, 
    0.002499716, -2.05553e-05, 0.0002411634, 0.007031661, 0,
  1.445625e-05, -5.528191e-08, -4.869031e-05, 0.02461677, -3.064023e-05, 
    0.009247381, 0.001182981, 0, 0, 0, 0, -9.10536e-06, 3.547126e-05, 
    0.002122973, 0.003022506, 3.452778e-05, 0.001407566, 0.00772771, 
    0.02837292, 0.007382915, 0.03716985, 0.02021425, 0.005037869, 
    0.002940356, 0.00612743, 0.008044433, 0.0166729, 0.02622486, 0.002338784,
  1.422251e-05, 0.001008015, 0, -3.504052e-06, 0.01594759, 0.001372472, 
    2.638683e-05, -3.340556e-06, -1.479111e-10, 0, -7.41966e-13, 
    -1.998323e-09, 0, -2.590912e-08, 5.993666e-05, 0.04577648, 0.08642297, 
    0.08504912, 0.04402977, 0.01100489, 0.006100169, 0.004644585, 
    -1.2028e-05, 0.001147616, -0.000206166, 0.008843996, 0.006679348, 
    0.001215233, -7.215612e-05,
  2.627122e-05, 0.0004223532, 1.808674e-08, -7.507042e-09, 1.567064e-06, 
    -1.681034e-08, -5.441294e-05, -3.099161e-05, -2.369807e-09, 
    -8.110791e-09, 1.204108e-08, 1.861083e-07, 6.479294e-07, 3.680818e-07, 
    0.005204255, 0.04612865, 0.07003355, 0.02250561, 0.003642045, 
    5.603737e-06, 6.88355e-05, 3.332739e-05, -6.931517e-05, 0.01889183, 
    0.009673898, -2.358872e-05, 0.007216202, 7.938199e-05, 9.403087e-05,
  0.004648967, 0.003721067, 2.157023e-06, 9.123691e-08, 1.212406e-06, 
    0.002411068, 0.09314236, 0.05895509, 0.07072681, 0.0103225, 0.002877953, 
    0.03656054, 0.02428925, 0.03454594, 0.02457944, 0.0007676451, 
    2.11411e-07, -1.64435e-08, 7.649357e-07, 0.01119347, 0.0012021, 
    6.451433e-05, 0.001695847, 0.001854958, 0.0419034, 0.04284737, 
    0.01860088, 2.666707e-05, 7.116076e-05,
  0.08214649, 0.3008662, 0.2281179, 0.0001099518, 5.08023e-05, 0.1881109, 
    0.1326342, 0.2646042, 0.4094155, 0.3527321, 0.3461715, 0.2071249, 
    0.2409277, 0.07769839, 0.05525686, 0.00413458, 0.001235031, 0.0001160051, 
    5.874947e-05, 0.03910004, 0.03806615, 0.03165842, 0.1126411, 0.209888, 
    0.02497765, 0.0001053504, 0.008771579, 0.05970509, 0.0201473,
  0.4325725, 0.3566338, 0.2900557, 0.01935619, 0.001843409, 0.0544444, 
    0.1093676, 0.3292532, 0.1653044, 0.07647513, 0.1568196, 0.1317706, 
    0.1842445, 0.1464996, 0.1654013, 0.1852072, 0.1069816, 0.1410632, 
    0.1349824, 0.1662247, 0.1712683, 0.3175635, 0.2875664, 0.1403468, 
    0.06888334, 0.07975212, 0.1615964, 0.2176418, 0.2717985,
  1.896029e-05, 0.002759917, 0.003484778, 0.005982502, 0.02236372, 
    0.07774913, 0.2517695, 0.2059575, 0.3270203, 0.2281503, 0.201826, 
    0.1307552, 0.2825445, 0.3054706, 0.2526327, 0.1197579, 0.01043284, 
    4.674159e-06, 0.01442342, 0.003893395, 0.04001063, 0.1967951, 0.1275568, 
    0.08166529, 0.07084208, 0.009828597, 0.0001232918, 0.002583616, 
    3.905703e-05,
  4.341488e-06, 0, 0, -2.417797e-09, 1.933045e-07, 1.394256e-05, 0.08353089, 
    0.05144641, 0.1004989, 0.1051253, 0.1557251, 0.112081, 0.2391766, 
    0.1657033, 0.2255542, 0.05077263, 0.07019242, 0.02721978, 0.008370291, 
    0.004726426, 0.02957031, 0.204219, 0.3377766, 0.1564461, 0.07406028, 
    0.1048903, 0.02395801, -2.855469e-06, -0.000124555,
  0.01568588, 0.00339105, 0.0001998201, 0.0002275859, -1.720796e-05, 
    -5.891257e-05, 4.519315e-06, 0.05489721, 0.07576043, 0.1017299, 
    0.2175533, 0.2290247, 0.07016724, 0.1481574, 0.1656155, 0.1353191, 
    0.1401992, 0.05690609, 0.03628066, 0.0009269874, 0.007542076, 0.05332682, 
    0.05095465, 0.08928492, 0.1896924, 0.06483819, 0.101844, 0.0408181, 
    0.009527181,
  0.008680499, 0.01062081, 0.07078166, 0.01125937, 0.01180104, 0.01882291, 
    0.001137817, 0.0002298349, 0.04942827, 0.08343315, 0.1298685, 0.1853018, 
    0.1068373, 0.2364315, 0.1813587, 0.1313021, 0.05126804, 0.0560573, 
    0.05104323, 0.00319844, 0.01623312, 0.04557758, 0.04076744, 0.03340047, 
    0.02933988, 0.06491302, 0.04764775, 0.029208, 0.02035202,
  0.0160387, 0.008369292, 0.0199488, 0, -0.0002264575, 0.02458193, 
    0.01114465, -0.0003099657, 0.00331592, 0.04977356, 0.06377792, 
    0.09345688, 0.04399346, 0.03718682, 0.0593368, 0.04202861, 0.01997279, 
    0.001540074, 0.0004406938, -4.083898e-05, 0.01879591, 0.01139085, 
    0.02297767, 0.008789419, 0.02632609, 0.01272036, 0.005092022, 
    0.006391515, -6.308713e-05,
  0, -1.270207e-05, 0.001379762, -0.0002770561, 0.0009035292, 0.003907763, 
    0.01256845, 0.002517218, -2.361037e-07, 0.006214858, 0.00647116, 
    0.002255222, 0.001096791, 0.002874945, -4.872314e-05, -1.965856e-05, 
    0.0001356947, -3.204709e-05, 0.0001313901, -0.0001361278, 0.01875028, 
    0.001596373, 0.0009408633, -7.510161e-05, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, -0.0001379214, -4.165209e-05, -6.021709e-05, 
    1.237761e-09, 1.197277e-06, 8.480544e-07, 0.001386237, 0.003845043, 
    -2.879415e-09, -4.57221e-07, -2.18572e-05, 4.976862e-06, -3.768616e-06, 
    0.004619523, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, -1.042715e-05, 0.00561272, -1.586611e-05, 0, 0, 0, 0, 
    -5.929327e-05, 3.412312e-06, 0.001085394, 0, 0, 0, -8.458986e-06, 0, 0, 
    0, 0, 0, -8.274244e-06, 0, 0, 0, 0, 0, 0,
  -2.418455e-09, 0, 0.001754406, 0.003987315, 0.03333492, 0.0007039567, 
    0.007211696, 0.0009727411, 0.0006612338, -1.794329e-05, -7.882827e-07, 
    0.0005661712, 0, -0.0001355504, 7.938858e-06, -7.472316e-06, 0.008251427, 
    0.000541592, 0, -6.250252e-05, 0.0001337319, 1.024875e-05, 0.001597296, 
    0.003120999, 0.003190766, 0.0009896512, 0.004845298, 0.01339992, 
    -3.877654e-09,
  0.006067787, -9.546709e-05, 0.0005048527, 0.0405437, 0.006257299, 
    0.01645462, 0.009803605, -1.825056e-05, -2.253162e-06, -8.659812e-07, 
    5.01465e-05, 0.001573865, 0.004737416, 0.003836934, 0.01338839, 
    0.00342878, 0.007852229, 0.02016805, 0.05624932, 0.02246739, 0.07106271, 
    0.0474896, 0.02165969, 0.008914732, 0.01710297, 0.03222182, 0.04540347, 
    0.03745731, 0.0170643,
  0.0006475855, 0.009726916, 4.098185e-05, 0.001600488, 0.02082318, 
    0.01523781, 0.0004403828, 0.0005057291, 8.827946e-07, 7.825714e-09, 
    -9.169877e-12, -1.99461e-09, 6.339299e-09, -1.031084e-06, 0.0006092073, 
    0.06179627, 0.14207, 0.1645541, 0.1001791, 0.04437264, 0.02656266, 
    0.03053017, 0.001909212, 0.003244685, 0.007515389, 0.0263441, 0.04138116, 
    0.03594866, 0.003180921,
  6.550464e-06, 4.584802e-05, 8.235525e-06, -3.976429e-09, 4.765681e-05, 
    -2.801723e-07, -2.027079e-07, 3.226275e-05, -1.230912e-08, 9.907009e-07, 
    1.945618e-07, 1.038934e-07, 1.161658e-06, 1.62131e-06, 0.01921596, 
    0.04424536, 0.04658468, 0.01291308, 0.008459629, -3.26391e-07, 
    1.681906e-05, 9.517532e-06, 1.791866e-06, 0.01043975, 0.01401709, 
    0.003819734, 0.0001640613, 0.0001530689, 4.659928e-06,
  2.656542e-05, 8.895672e-05, 1.544733e-06, -6.394137e-10, 3.786401e-06, 
    0.001976029, 0.0827168, 0.04270872, 0.05772259, 0.006663411, 
    0.0005424599, 0.02167353, 0.005831842, 0.02778886, 0.01708084, 
    0.001743179, 4.433317e-05, 5.107179e-07, 1.730863e-08, 0.0001850657, 
    3.671911e-05, -3.247088e-05, 8.219492e-05, 0.001067606, 0.03304515, 
    0.02760871, 0.007209179, 0.0001695368, 2.028608e-06,
  0.07012687, 0.2338197, 0.1500881, 5.409351e-06, 4.258653e-05, 0.1141487, 
    0.07034616, 0.1879713, 0.3472611, 0.3147277, 0.2076651, 0.1692883, 
    0.2250724, 0.0639842, 0.03407567, 0.001328845, 2.165552e-05, 
    1.371677e-05, 1.01614e-05, 0.005144835, 0.003432952, 0.002281169, 
    0.08009159, 0.1475393, 0.008518527, 0.0001841226, 0.003219998, 
    0.05087754, 0.001445003,
  0.3853228, 0.3019428, 0.2175017, 0.06826893, 0.000173099, 0.0397064, 
    0.04791077, 0.181775, 0.08552528, 0.02501617, 0.06211946, 0.06880611, 
    0.1541009, 0.1132483, 0.128957, 0.1245331, 0.08326483, 0.1218138, 
    0.1246595, 0.1541875, 0.1822221, 0.2790709, 0.2232225, 0.1064464, 
    0.04255237, 0.04558682, 0.1130354, 0.1886563, 0.2392087,
  3.271583e-06, 0.0003082929, 0.001162048, 0.003780696, 0.02920303, 
    0.06270522, 0.2177714, 0.1530884, 0.3175968, 0.1728104, 0.2016787, 
    0.1167823, 0.2467051, 0.2594109, 0.2226393, 0.09570458, 0.0007261072, 
    1.947827e-06, 0.01027395, 0.004654961, 0.04184646, 0.1499065, 0.07436997, 
    0.05318338, 0.03092011, 0.008237129, 4.006067e-05, 0.0006508024, 
    0.0002112031,
  -1.432315e-06, 0, 0, -1.128312e-09, 9.366114e-08, 5.247733e-06, 0.08791962, 
    0.1426025, 0.1670861, 0.06018672, 0.1376353, 0.08085811, 0.2251043, 
    0.1451082, 0.2378957, 0.05224228, 0.1365461, 0.02144681, 0.002322813, 
    0.005274509, 0.03047964, 0.1403536, 0.2602745, 0.1155992, 0.05177399, 
    0.09679691, 0.03316842, -1.132404e-07, 0.0005016949,
  0.04974744, 0.01530914, 0.004951439, 0.0036803, 0.001531387, 0.003315777, 
    0.0003990073, 0.1076733, 0.1385527, 0.1500604, 0.2152308, 0.2110184, 
    0.04524145, 0.1439078, 0.1483066, 0.1529273, 0.1476022, 0.105281, 
    0.04299196, 0.003403055, 0.08753918, 0.06549691, 0.06628104, 0.08553093, 
    0.1888411, 0.09348751, 0.1441559, 0.0666917, 0.03876536,
  0.06484488, 0.06119414, 0.142735, 0.04741398, 0.04409773, 0.1093111, 
    0.06880006, 0.0001373861, 0.0725157, 0.1811228, 0.1776627, 0.2330535, 
    0.1552602, 0.2552498, 0.1979658, 0.1362723, 0.09057381, 0.08437435, 
    0.1497578, 0.006693043, 0.0978765, 0.1222321, 0.09471164, 0.07490569, 
    0.08738112, 0.1374682, 0.1712273, 0.1135632, 0.133173,
  0.049851, 0.01243119, 0.04061975, 0.01187318, 0.006854673, 0.08128558, 
    0.06890246, 0.02540107, 0.03533799, 0.1088048, 0.1779453, 0.1668856, 
    0.06166665, 0.06249697, 0.1387254, 0.08768903, 0.07536785, 0.03060231, 
    0.004850545, 0.03321957, 0.04184879, 0.0751302, 0.0967228, 0.07399602, 
    0.05585032, 0.0242987, 0.02934182, 0.04398473, 0.01912065,
  0, 0.0001149338, 0.001823708, 0.006042243, 0.009374836, 0.006465342, 
    0.01710053, 0.007859873, 0.0212658, 0.0347636, 0.03429709, 0.05384485, 
    0.06062831, 0.06656369, 0.03108173, 0.02326404, 0.01700622, 0.02225563, 
    0.03284104, 0.01776111, 0.0488692, 0.02390637, 0.02193468, 0.004872754, 
    -7.017882e-05, -2.336087e-05, -2.101469e-06, 0.007532853, 2.590614e-05,
  -3.918674e-08, 0, 0, 0, -5.790786e-05, 0, 0, -0.0004740427, -2.678653e-05, 
    -2.055532e-05, 1.807645e-06, -6.888662e-06, -5.121472e-05, 0.002234011, 
    0.004995116, -8.027742e-05, 0.002349736, 0.001269283, 0.002959954, 
    -4.786591e-05, 0.007115882, -0.000318518, 3.820553e-05, -6.056871e-08, 
    -1.170955e-05, 0, 0, -3.62369e-07, 1.308431e-06,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.836605e-07, -2.157704e-05, 0, 0, 0, 
    0, 0, 0, 0, -1.405658e-05, 0, 0, 0, 0, 0, 0, 0,
  0, -3.875256e-06, -8.678374e-06, 0.001325072, 0.008339694, 0.004447701, 
    0.001984823, 1.370227e-05, 0, 0, 0.001983746, 0.0006553981, 0.003263999, 
    0.002510664, -2.32454e-05, 0, -5.084624e-05, -4.106812e-08, 
    -6.882015e-06, 0.003703995, 0, -9.843371e-06, -3.590302e-05, 
    0.0007570133, -0.0001790229, 0, 0, -5.250899e-06, 0,
  0.003466818, -5.222123e-06, 0.003855148, 0.008183463, 0.06615169, 
    0.01762894, 0.01520747, 0.005486659, 0.00342645, 8.105245e-05, 
    0.0004132777, 0.003183819, -4.589723e-05, 0.001603402, 0.001255176, 
    1.012329e-05, 0.01054831, 0.01455438, 0.0001367782, 0.004437262, 
    0.005631061, 0.007784175, 0.0102379, 0.009536568, 0.008018293, 0.0137145, 
    0.03082861, 0.04432604, 0.0007522773,
  0.07219977, 0.00955693, 0.03160876, 0.09431819, 0.02053902, 0.03776002, 
    0.04881765, 0.03456041, 0.01974793, 0.01112947, 0.01476937, 0.01834178, 
    0.02810865, 0.009454425, 0.04009528, 0.02625208, 0.02196862, 0.04750324, 
    0.1205995, 0.09069753, 0.1312719, 0.1154728, 0.09698512, 0.04246081, 
    0.0757505, 0.1381023, 0.1452252, 0.119034, 0.1215907,
  0.00295888, 0.006796498, 0.007932193, 0.02067163, 0.05602093, 0.02119742, 
    0.002079967, 0.01076495, 0.006508003, -1.267394e-05, 2.619358e-08, 
    -1.926484e-09, 6.156594e-06, -3.305236e-05, 0.002890982, 0.06941951, 
    0.1814841, 0.2188005, 0.1451136, 0.06049886, 0.03283334, 0.01230485, 
    0.001563557, 0.002199227, 0.007845594, 0.02450023, 0.05029375, 
    0.03277577, 0.01203221,
  1.492897e-06, 6.275356e-06, 2.655981e-06, -2.230524e-09, 0.0002925864, 
    1.433654e-07, 3.558844e-06, 0.001798947, -3.136181e-08, 2.43231e-06, 
    1.063534e-06, 5.060823e-08, 7.297171e-07, 0.000190473, 0.04363481, 
    0.05088966, 0.03640136, 0.005589369, 0.0002312896, -5.612523e-08, 
    5.811676e-07, 4.490354e-06, 4.372871e-06, 5.524453e-05, 0.01092264, 
    0.004077906, 0.0004529745, 0.000246456, -0.0001216587,
  7.051596e-07, 1.647738e-05, 1.901145e-07, -1.526947e-12, -1.090427e-06, 
    0.002888352, 0.07958864, 0.04516567, 0.05587007, 0.00912834, 
    0.0003152495, 0.01655482, 0.001478536, 0.0297779, 0.01824346, 0.00366199, 
    0.0002925493, 1.010496e-07, -2.170495e-09, 5.678385e-06, 3.351051e-06, 
    -5.372509e-08, 0.0002510091, 0.001123074, 0.03223293, 0.01014273, 
    0.0001041855, 1.10563e-06, 2.268433e-07,
  0.02467112, 0.1816158, 0.0890198, 1.385104e-06, 2.090483e-05, 0.09563157, 
    0.05230907, 0.1284567, 0.3086419, 0.2719301, 0.1522348, 0.1470608, 
    0.2334601, 0.06679279, 0.03843493, 0.001258336, 1.39058e-05, 
    8.982443e-06, 1.287871e-05, 8.71075e-05, 0.001908464, 0.00114607, 
    0.04987723, 0.1173578, 0.007038019, 0.0001627981, 0.003269571, 
    0.03415628, 9.835316e-05,
  0.3581684, 0.2809675, 0.1710068, 0.04614966, 0.0006705035, 0.01810937, 
    0.02845406, 0.09438039, 0.04852975, 0.01635948, 0.02281255, 0.05038037, 
    0.1352117, 0.09495256, 0.1177825, 0.08964523, 0.07079289, 0.1158654, 
    0.1082277, 0.1665669, 0.1783729, 0.2410467, 0.2176924, 0.09702566, 
    0.03970262, 0.03868335, 0.1004839, 0.1741434, 0.2570384,
  9.902624e-07, 1.062042e-05, 2.700388e-06, 0.0006454575, 0.02446574, 
    0.06419645, 0.1877237, 0.1112413, 0.2835271, 0.1301817, 0.1722854, 
    0.09941962, 0.2000351, 0.2162204, 0.2057168, 0.0771635, 0.0005535032, 
    2.26265e-06, 0.01185837, 0.003428041, 0.04243299, 0.1275738, 0.05568698, 
    0.04029749, 0.02754497, 0.00237848, 5.072799e-05, 0.0004025477, 
    0.002990805,
  -9.295927e-08, 0, 0, -8.544571e-10, 3.474111e-09, 5.037682e-07, 0.0858729, 
    0.189135, 0.1710823, 0.04372998, 0.1219191, 0.06297999, 0.2160537, 
    0.1308263, 0.2159775, 0.03822838, 0.0923508, 0.009528956, 0.0001918825, 
    0.01185798, 0.03490575, 0.09530704, 0.235194, 0.1031964, 0.04559395, 
    0.081923, 0.01957957, -5.189726e-08, -1.868104e-05,
  0.04464616, 0.01054397, 0.002844852, 0.02368381, 0.002272695, 0.003003204, 
    0.001293668, 0.1441082, 0.1676855, 0.1769001, 0.1718703, 0.2030913, 
    0.04733939, 0.139954, 0.1438629, 0.1311554, 0.1193305, 0.0939194, 
    0.0452668, 0.0009688221, 0.1164281, 0.04013453, 0.05341073, 0.0706104, 
    0.1646621, 0.08633193, 0.1263539, 0.05310449, 0.03004432,
  0.1142134, 0.1622889, 0.223729, 0.145722, 0.05480841, 0.1145195, 
    0.06046147, 0.02457617, 0.148078, 0.1961028, 0.1503361, 0.2046764, 
    0.1322602, 0.2211368, 0.1437851, 0.1325023, 0.09007862, 0.1184549, 
    0.1864888, 0.05172839, 0.09412978, 0.09286273, 0.09933863, 0.1301535, 
    0.1354787, 0.1850059, 0.2124377, 0.1429024, 0.185743,
  0.1504328, 0.09050486, 0.09277894, 0.05421025, 0.08818185, 0.1867451, 
    0.1660201, 0.07088253, 0.08815653, 0.1681575, 0.2162486, 0.2090548, 
    0.09852442, 0.07367986, 0.1652885, 0.09319168, 0.09603782, 0.0950163, 
    0.07510688, 0.1025449, 0.1536895, 0.1843062, 0.1451585, 0.1195626, 
    0.144497, 0.1124721, 0.09828819, 0.1237037, 0.06870542,
  0.02590693, 0.01399397, 0.02932544, 0.0373815, 0.06982265, 0.06746519, 
    0.08970191, 0.07529428, 0.06286485, 0.09482803, 0.1231228, 0.140382, 
    0.09922478, 0.1211416, 0.1490302, 0.06960588, 0.1054536, 0.08147027, 
    0.05239247, 0.08362442, 0.139203, 0.1425005, 0.08563933, 0.03534657, 
    0.07890543, 0.000166788, 1.540354e-05, 0.05986828, 0.04632514,
  0.02180598, 0.01446398, 0.02609337, 0.01331014, 0.004853562, 0.01767511, 
    0.001259215, -0.00041048, 0.001625058, 6.626453e-05, 1.599786e-05, 
    -0.0001778062, -0.0007108346, 0.02021411, 0.01643613, 0.01872229, 
    0.02323901, 0.04402227, 0.02765061, 0.05438154, 0.139253, 0.1455802, 
    0.07012052, 4.623936e-05, -0.0009241656, -0.0002964838, -0.0003235211, 
    -0.002314421, 0.02705524,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0003153392, -0.0001521938, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.836605e-07, -2.157704e-05, 
    0.0002169559, 0, 0, 0, 0, 0, 0, -2.728458e-05, 2.353558e-05, 0, 0, 0, 
    0.0001265367, 0, 0,
  0.00219188, 1.592413e-05, 4.031841e-05, 0.002093346, 0.01182481, 
    0.01133506, 0.01006185, 0.001942888, 0, 0.000473987, 0.004692862, 
    0.005656148, 0.006341174, 0.00492952, 0.0005183928, 0.0001232959, 
    0.006756111, 0.00137009, 0.004326542, 0.01189534, 0.0002969278, 
    0.003448277, 0.005039493, 0.004203418, 0.003518921, -6.696288e-05, 
    0.000807436, 0.002415128, 0.007359247,
  0.08859549, 0.0424505, 0.03066622, 0.04693598, 0.1565614, 0.08799631, 
    0.05664311, 0.03560745, 0.02687847, 0.02941191, 0.017885, 0.006925193, 
    0.00794463, 0.01759817, 0.01303024, 0.03347801, 0.04938801, 0.04559971, 
    0.02825918, 0.01949943, 0.03855577, 0.05540705, 0.06184979, 0.03815606, 
    0.04882422, 0.0597747, 0.05632798, 0.09117483, 0.07577156,
  0.1855311, 0.08607762, 0.06803539, 0.1204345, 0.0454897, 0.08120312, 
    0.0828459, 0.07296913, 0.04952103, 0.03703471, 0.04291699, 0.03246029, 
    0.0477737, 0.01831761, 0.0905696, 0.08764263, 0.03817698, 0.07618017, 
    0.1360875, 0.1148627, 0.1922611, 0.1603687, 0.1602837, 0.07849666, 
    0.1295517, 0.197167, 0.1514216, 0.1360361, 0.1991769,
  0.0009784648, 0.006568023, 0.02212667, 0.01314746, 0.0551776, 0.01938061, 
    0.004318592, 0.009134052, 0.005972612, 0.0007596262, 4.508812e-08, 
    -3.271409e-08, 0.008884535, -0.0001053274, 0.006810193, 0.07569404, 
    0.2039043, 0.2178712, 0.1384157, 0.04313642, 0.01919251, 0.007520194, 
    0.0003356379, 0.001167997, 0.01519579, 0.02723871, 0.05034837, 
    0.03753092, 0.007033097,
  4.446331e-07, 6.319552e-07, 4.204844e-07, -1.208938e-10, 0.0004735179, 
    -1.767341e-06, -8.77128e-06, 0.004334808, -3.816161e-08, 1.220975e-05, 
    2.08324e-06, 1.922841e-05, 2.403893e-07, 0.0009013843, 0.06978057, 
    0.04791668, 0.04537585, 0.01060177, -7.863334e-05, -1.196807e-08, 
    1.308578e-08, 1.260516e-06, 1.656143e-06, 8.257241e-06, 0.00451676, 
    0.005582752, 0.002678143, 0.007788516, 0.0001434078,
  2.795889e-07, 2.186048e-06, 4.324117e-08, 0, 4.309368e-08, 0.003444125, 
    0.09376086, 0.05370708, 0.04370677, 0.007970089, 0.0005339879, 
    0.02299544, 0.001625699, 0.03308867, 0.01301774, 0.008024122, 
    0.0001593896, 1.290796e-07, -9.864354e-11, 1.737195e-06, 1.104364e-07, 
    2.066592e-07, 2.995974e-07, 0.001180016, 0.02583735, 0.003321777, 
    7.390807e-06, 4.645823e-07, 4.819899e-08,
  0.001584168, 0.1405804, 0.05292914, 7.971639e-07, 2.312501e-05, 0.08157754, 
    0.03180255, 0.08016952, 0.2431233, 0.2255629, 0.1058985, 0.1326173, 
    0.2356227, 0.0706301, 0.03470429, 0.002445801, 0.0001000245, -6.5266e-07, 
    1.470383e-05, 1.19724e-05, 9.914165e-05, 0.005303054, 0.04729792, 
    0.07071956, 0.007390378, 0.0001268838, 0.001405551, 0.003621301, 
    8.934071e-05,
  0.3169554, 0.2387117, 0.1147659, 0.05500266, 0.003642801, 0.008906828, 
    0.02745701, 0.05670026, 0.03106802, 0.01349237, 0.01004244, 0.04230182, 
    0.1164128, 0.07824267, 0.101243, 0.06639237, 0.0547494, 0.116356, 
    0.08382718, 0.1813763, 0.1479806, 0.2044238, 0.1942728, 0.07841239, 
    0.03316635, 0.03455572, 0.07838293, 0.1643463, 0.2724577,
  4.010082e-05, 1.790472e-06, 2.467227e-06, 1.942248e-05, 0.02571383, 
    0.0557284, 0.1847547, 0.07419129, 0.2707236, 0.09959286, 0.1340957, 
    0.07648363, 0.1369473, 0.1847183, 0.171201, 0.08054604, 0.007517723, 
    1.576806e-06, 0.013083, 0.01310161, 0.04073687, 0.1014413, 0.03592078, 
    0.02775335, 0.0203435, 0.001158077, 0.0001619925, 0.0003143296, 
    0.001618689,
  1.618085e-07, 5.273046e-10, 0, -5.277618e-10, -1.17473e-09, -1.751475e-07, 
    0.09024672, 0.1671999, 0.1733543, 0.04652827, 0.1073386, 0.05859586, 
    0.2002904, 0.1209125, 0.2064133, 0.04777608, 0.06190138, 0.00395081, 
    0.000137155, 0.0127534, 0.03176682, 0.06969528, 0.2016317, 0.07815364, 
    0.03807906, 0.05999334, 0.007017369, -4.151788e-08, -5.917049e-05,
  0.03632131, 0.006302655, 0.002347096, 0.02090609, 0.004313191, 0.001515863, 
    0.01275419, 0.1679573, 0.1689108, 0.1474949, 0.1404979, 0.1798579, 
    0.04130894, 0.147412, 0.1282564, 0.1243294, 0.0995095, 0.08555195, 
    0.0477514, 4.573553e-05, 0.0932894, 0.03911631, 0.04664296, 0.05736546, 
    0.1430687, 0.07659721, 0.1129086, 0.04545881, 0.01831231,
  0.1238665, 0.1891055, 0.2410987, 0.1144926, 0.03808185, 0.1137848, 
    0.05319764, 0.05322061, 0.1739704, 0.1753722, 0.1114125, 0.1729735, 
    0.1178476, 0.1998287, 0.1210396, 0.1269123, 0.102433, 0.1334116, 
    0.1918374, 0.05392273, 0.07564683, 0.07105338, 0.07942414, 0.1310203, 
    0.1163551, 0.1629614, 0.1669424, 0.1505738, 0.1618602,
  0.1506517, 0.1147176, 0.1359498, 0.1106717, 0.1257213, 0.1895895, 
    0.2080422, 0.1173279, 0.1107208, 0.1934015, 0.2176313, 0.1846142, 
    0.07706314, 0.06909782, 0.1594257, 0.117247, 0.1267039, 0.1702503, 
    0.2013586, 0.1363599, 0.160458, 0.1536727, 0.1527099, 0.1381723, 
    0.1795421, 0.2572791, 0.1353887, 0.1592427, 0.1681805,
  0.1282476, 0.1571618, 0.08643093, 0.1085945, 0.1464364, 0.1370142, 
    0.1896173, 0.1370616, 0.1419986, 0.1762782, 0.1672233, 0.180633, 
    0.1367884, 0.1885402, 0.203871, 0.1491699, 0.1453161, 0.1646828, 
    0.1596915, 0.1920078, 0.1657503, 0.1474129, 0.1199509, 0.06439377, 
    0.1231981, 0.00995142, 0.001639425, 0.1580565, 0.1513014,
  0.06204029, 0.09640746, 0.1322977, 0.153333, 0.1466272, 0.08735581, 
    0.04816258, 0.0275104, 0.02649868, 0.0114658, 0.001440481, -0.0002716768, 
    6.008682e-05, 0.03360104, 0.05316504, 0.05064588, 0.08791273, 0.1843432, 
    0.2103958, 0.1664833, 0.2277043, 0.2517357, 0.1725407, 0.08683624, 
    0.04515295, 0.002578149, -0.003543657, 0.03883754, 0.06334755,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.993262e-05, 7.908513e-05, 0, 0, 0, 
    0, 0, 0, 0, 0.001748716, 0.0002997036, 0, 0, 0, 0, 0,
  -1.334777e-05, 0, 0, 0, -4.230684e-05, 0, 0, 0, 0, 0, 0, 0, -2.836605e-07, 
    -2.293873e-05, 0.0008725686, 0, -3.347696e-05, 0, 0.0005026205, 
    -3.413355e-05, 0.00236628, 0.0004666095, 0.003756893, 0.0008439255, 
    0.00213898, 0.0002762444, 0.002613856, -2.293116e-05, -8.819324e-05,
  0.06387129, 0.03744086, 0.01505878, 0.02468867, 0.04926442, 0.04591222, 
    0.04422037, 0.02608167, 0.005919452, 0.007430786, 0.01945295, 0.01722981, 
    0.01572477, 0.02649583, 0.01282682, 0.01798112, 0.03000758, 0.03766213, 
    0.02079231, 0.02452638, 0.007854312, 0.01547929, 0.01472932, 0.0169892, 
    0.02891977, 0.0100879, 0.008609506, 0.02816574, 0.06546111,
  0.1401121, 0.1485988, 0.2011769, 0.1656045, 0.2316011, 0.1832992, 
    0.1198148, 0.08708934, 0.09347472, 0.1002861, 0.08794041, 0.1087655, 
    0.09705735, 0.1018402, 0.1072363, 0.1667572, 0.1121437, 0.07868312, 
    0.06232598, 0.0440468, 0.08713796, 0.1264777, 0.1491769, 0.09784448, 
    0.1185313, 0.1177369, 0.1238968, 0.136321, 0.1250567,
  0.2076756, 0.1199425, 0.08673082, 0.1320727, 0.03821911, 0.08116246, 
    0.09381893, 0.107976, 0.07263242, 0.06532297, 0.06946559, 0.08718114, 
    0.0695636, 0.08286224, 0.1172996, 0.1432523, 0.05977245, 0.0714907, 
    0.1231119, 0.1395575, 0.1803603, 0.1717964, 0.1640073, 0.09853108, 
    0.1024214, 0.1532096, 0.113758, 0.1252577, 0.2165498,
  0.000851689, 0.003744225, 0.01783255, 0.006793121, 0.05200113, 0.0261917, 
    0.01008845, 0.008227023, 0.004055921, 0.0003748105, -8.039414e-07, 
    -3.603304e-06, 0.01564733, 0.001797124, 0.02398394, 0.08097906, 0.227835, 
    0.2188081, 0.1296157, 0.03573687, 0.01410984, 0.006549288, -4.203796e-06, 
    0.001637241, 0.02609968, 0.0337755, 0.05934023, 0.04017241, 0.007051605,
  1.605825e-08, 1.837677e-07, 1.428796e-07, -3.854203e-07, 0.0004217345, 
    -6.282602e-06, -1.566542e-07, 0.002748835, 4.546958e-07, 0.0003467842, 
    3.29654e-05, 0.001223963, 4.160976e-06, -9.917736e-05, 0.07277064, 
    0.04643121, 0.0575349, 0.00943295, 0.0008545056, -5.655378e-10, 
    -2.857627e-10, 1.416559e-07, 1.61238e-07, 1.41207e-06, 0.0007997651, 
    0.007531092, 0.00135642, 9.477943e-05, 1.079757e-06,
  2.538866e-07, 3.809014e-07, -1.441453e-10, 0, 5.687679e-09, 0.002970306, 
    0.09482662, 0.06738225, 0.0368566, 0.007851988, 0.0002494977, 0.01428512, 
    0.001969182, 0.03421782, 0.01185569, 0.01133313, 0.0001768768, 
    4.87656e-08, 0, 4.697181e-07, 1.380223e-08, 2.461425e-07, 3.147405e-06, 
    0.001188769, 0.02093852, 0.001291129, 2.658007e-06, 1.67074e-07, 
    7.283752e-09,
  0.0002468254, 0.09547417, 0.03811819, 9.890217e-07, 2.606209e-05, 
    0.06775271, 0.0203317, 0.05354485, 0.1744438, 0.1972036, 0.07390346, 
    0.116371, 0.2297007, 0.05738484, 0.03031389, 0.002632621, 0.0001689065, 
    -7.85503e-06, 1.496302e-05, -6.031786e-06, -2.240393e-06, 0.00260532, 
    0.04076302, 0.04371031, 0.00826731, 0.0001739373, 0.0001285507, 
    3.833535e-05, 5.116113e-05,
  0.2569163, 0.1858953, 0.08601162, 0.06500633, 0.007615411, 0.006556301, 
    0.02058421, 0.02566647, 0.01926595, 0.009879406, 0.004390826, 0.03021004, 
    0.08450677, 0.05770649, 0.07629155, 0.05880272, 0.05128465, 0.1283383, 
    0.0861384, 0.2055704, 0.117869, 0.1403747, 0.1853325, 0.06668681, 
    0.02838324, 0.03131027, 0.05581719, 0.1631663, 0.2642154,
  5.457253e-05, 6.594873e-07, 1.26261e-06, 0.000111693, 0.02995181, 
    0.06718527, 0.1434504, 0.04717198, 0.2537084, 0.07127898, 0.09944449, 
    0.05426554, 0.07972039, 0.147395, 0.1080184, 0.06941085, 0.002124121, 
    4.953631e-06, 0.01231254, 0.005066324, 0.04090304, 0.0821825, 0.02292719, 
    0.01565103, 0.01287687, 0.00104263, 0.0001492881, 0.0004043088, 
    0.002247859,
  5.455981e-08, 1.054644e-08, 0, -2.034245e-10, -8.022681e-09, -1.778434e-06, 
    0.07598353, 0.1553873, 0.1787207, 0.03283763, 0.1075158, 0.04941948, 
    0.1860665, 0.1043773, 0.185928, 0.05770743, 0.04458763, 0.000595333, 
    2.327211e-05, 0.03476439, 0.03158109, 0.04263001, 0.1600291, 0.05095854, 
    0.02721916, 0.03909492, 0.001762497, -1.301223e-08, 4.679164e-05,
  0.02841202, 0.004028032, 0.003405007, 0.01453081, 0.005950952, 0.008714706, 
    0.04591374, 0.1673337, 0.1672309, 0.1319243, 0.113909, 0.1383449, 
    0.03286061, 0.1439708, 0.1345724, 0.1192362, 0.08923292, 0.06942811, 
    0.02303398, -5.653035e-05, 0.07592843, 0.03108354, 0.03886355, 0.0450643, 
    0.1270815, 0.06860638, 0.09852476, 0.04453362, 0.01086378,
  0.1371746, 0.1714211, 0.2298229, 0.0956253, 0.03317374, 0.09709904, 
    0.03893775, 0.04613007, 0.1750493, 0.1586193, 0.0854223, 0.1520251, 
    0.1127267, 0.1886907, 0.1100594, 0.1276356, 0.09476382, 0.131595, 
    0.1857243, 0.04072513, 0.06575086, 0.06117101, 0.06765237, 0.101163, 
    0.1044516, 0.1425513, 0.161313, 0.1419825, 0.1387887,
  0.1468083, 0.1856361, 0.136139, 0.09615777, 0.0996404, 0.1699299, 0.202547, 
    0.108549, 0.1206708, 0.2078427, 0.2084323, 0.1550053, 0.05846531, 
    0.06208904, 0.1449372, 0.1393841, 0.192157, 0.254431, 0.273761, 
    0.1194875, 0.1526662, 0.1321741, 0.1467485, 0.1630929, 0.1764269, 
    0.2565807, 0.1568309, 0.1778304, 0.1974453,
  0.1389959, 0.2152244, 0.1558729, 0.1615019, 0.1847592, 0.1669433, 
    0.2076151, 0.1682362, 0.1828181, 0.1784826, 0.1933544, 0.1926535, 
    0.1328327, 0.2125054, 0.2413388, 0.1644421, 0.2413562, 0.2012062, 
    0.1870332, 0.2120475, 0.1843492, 0.1537821, 0.1378784, 0.1177923, 
    0.1361265, 0.05012825, 0.01713576, 0.1374873, 0.140156,
  0.1081229, 0.151534, 0.1868734, 0.2110244, 0.2032295, 0.1978665, 0.1534675, 
    0.09595997, 0.1083698, 0.09414028, 0.07282874, 0.06642291, 0.04086667, 
    0.09871119, 0.08002459, 0.093623, 0.172338, 0.2483867, 0.2599845, 
    0.2079366, 0.2684833, 0.3402557, 0.2132493, 0.1531239, 0.08666507, 
    0.06057866, 0.06245756, 0.09326711, 0.1334103,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.000482158, 0.0001384062, 
    -7.969163e-07, 0, -4.85819e-05, 0.0002108449, -3.42015e-05, 
    -2.112095e-05, -1.073684e-05, 0.002558581, 0.00619718, -4.854861e-06, 0, 
    0, 0, 0,
  0.001356642, -0.0001026964, 1.310063e-05, 0.0001161233, -0.0001498248, 0, 
    0.0002690508, 0, 0, 0, -1.118149e-05, 0.0003290201, -0.000333059, 
    0.005257697, 0.02252178, 0.01024908, 0.005467386, -0.0003889739, 
    0.0002419555, 0.00296553, 0.009455111, 0.00541629, 0.004391161, 
    0.003229167, 0.007976079, 0.009351482, 0.007248433, 0.002445339, 
    0.004747775,
  0.133703, 0.1462498, 0.08394995, 0.06822267, 0.1023678, 0.0992393, 
    0.09273267, 0.05719241, 0.04171326, 0.04255757, 0.0517507, 0.08852085, 
    0.1216791, 0.1842649, 0.1772086, 0.1981282, 0.1939828, 0.1607423, 
    0.1051507, 0.08657446, 0.04533099, 0.06959888, 0.04009296, 0.04270184, 
    0.08799163, 0.09310177, 0.04340118, 0.1247484, 0.1295905,
  0.178103, 0.1636641, 0.2609028, 0.2056588, 0.2532019, 0.2039151, 0.155758, 
    0.1367549, 0.1499815, 0.1313671, 0.1958559, 0.2041779, 0.1770911, 
    0.1894412, 0.1323076, 0.193153, 0.1798278, 0.1463838, 0.1290306, 
    0.08883574, 0.1490006, 0.1691555, 0.1815037, 0.1547218, 0.170147, 
    0.1745899, 0.1873254, 0.194648, 0.1821398,
  0.1875777, 0.09355817, 0.08521312, 0.1398061, 0.04091824, 0.07930177, 
    0.09839524, 0.0956085, 0.07341524, 0.07155742, 0.07473328, 0.104131, 
    0.08076432, 0.08576316, 0.1480787, 0.1285243, 0.06004424, 0.0750655, 
    0.1108811, 0.1501911, 0.1776635, 0.171041, 0.162128, 0.0918562, 
    0.08842801, 0.1180291, 0.09270169, 0.1123543, 0.1969022,
  -0.0001285053, 0.001814848, 0.009746457, 0.003757958, 0.0532731, 
    0.05033613, 0.01497834, 0.005725484, 0.000103585, 0.0004598757, 
    -2.108455e-07, -5.214726e-05, 0.01535549, 0.008412579, 0.03512368, 
    0.09534463, 0.2134842, 0.2284479, 0.143394, 0.0204659, 0.01037927, 
    0.003195692, -2.460447e-05, 0.001458059, 0.03027743, 0.04252614, 
    0.06859583, 0.04783738, 0.01128008,
  -1.112125e-09, 7.880824e-08, 9.289308e-08, 5.731947e-05, 0.0001625785, 
    0.0004578552, -7.947238e-07, 0.01141576, -1.06894e-07, 0.002273543, 
    0.003175259, 0.004452673, 0.0003438549, -3.693676e-06, 0.06081765, 
    0.06300183, 0.05761967, 0.004559205, 0.0009148599, -2.030163e-09, 0, 
    8.927714e-08, 2.109469e-08, 4.989337e-07, -0.0002681274, 0.009666793, 
    8.753004e-05, 2.240184e-06, 4.66662e-08,
  2.241278e-08, 7.37649e-07, 3.225881e-09, 0, -9.459775e-08, 0.001789936, 
    0.1028586, 0.07099337, 0.03577879, 0.01227197, 0.0005866317, 0.01191707, 
    0.009371212, 0.05016289, 0.009079091, 0.02045565, 0.0001366152, 0, 0, 
    6.857646e-08, 1.696573e-08, 4.09535e-09, 2.005771e-06, 0.00141133, 
    0.0160988, 0.001448795, 8.285057e-07, 3.209124e-08, 4.975672e-08,
  0.0002044692, 0.07170243, 0.03024481, 7.950854e-07, 3.241443e-05, 
    0.05906838, 0.01500041, 0.0289051, 0.1053515, 0.192396, 0.05460459, 
    0.1101911, 0.2381854, 0.04409798, 0.0264452, 0.003276108, 7.734526e-05, 
    -6.460619e-06, 0.0002539087, -2.05322e-05, 7.293159e-06, 0.01889559, 
    0.05044261, 0.03001054, 0.01013892, 0.0004439093, 0.0006053608, 
    2.92763e-05, 1.406978e-05,
  0.2217822, 0.1570399, 0.07096089, 0.06648095, 0.01361104, 0.004975711, 
    0.02256962, 0.01068957, 0.01333328, 0.007366071, 0.004246215, 0.02152722, 
    0.06823659, 0.046235, 0.06194878, 0.05023946, 0.0536126, 0.1442405, 
    0.09201535, 0.2214925, 0.1211825, 0.08936206, 0.1879727, 0.06226075, 
    0.02243328, 0.03208057, 0.05130965, 0.1546624, 0.2728208,
  4.412255e-05, 2.181394e-06, 7.954981e-07, 0.0004215809, 0.02916111, 
    0.09539408, 0.1515747, 0.03104207, 0.2158485, 0.05744778, 0.08102802, 
    0.04693834, 0.05916672, 0.1222953, 0.06299733, 0.05403076, 0.0001866344, 
    8.760041e-06, 0.006450207, 0.005814093, 0.04416227, 0.08109468, 
    0.01536536, 0.01256095, 0.008914374, 0.001037332, 9.163213e-05, 
    0.000275336, 0.005622492,
  -6.187917e-07, -2.440313e-06, 0, -2.410709e-10, -1.785791e-07, 
    -1.222857e-05, 0.06013826, 0.1596482, 0.1953526, 0.04595547, 0.1042621, 
    0.04906548, 0.1777353, 0.08367115, 0.1396319, 0.04941888, 0.03633561, 
    0.0001237678, 2.420604e-05, 0.02113173, 0.02643377, 0.02427157, 
    0.1238295, 0.03266077, 0.01666916, 0.02294747, 0.0003900131, 
    1.155398e-11, 0.0009308343,
  0.02278162, 0.001850324, 0.004602012, 0.01323461, 0.01403702, 0.00953544, 
    0.07993784, 0.1588127, 0.147423, 0.1148753, 0.1077595, 0.1369526, 
    0.04313091, 0.2013638, 0.1416219, 0.111425, 0.07937799, 0.08274814, 
    0.02180673, -6.396867e-05, 0.06052408, 0.02714517, 0.02985324, 0.0397543, 
    0.1099507, 0.05734412, 0.07604366, 0.0427665, 0.007712962,
  0.1540866, 0.1606477, 0.2181268, 0.080225, 0.02759353, 0.08061472, 
    0.02905936, 0.04599835, 0.1889156, 0.1453148, 0.08207435, 0.1311611, 
    0.1334213, 0.1818099, 0.1006613, 0.1190767, 0.09126863, 0.1271632, 
    0.2012076, 0.03349272, 0.0506764, 0.06807429, 0.0751626, 0.09706635, 
    0.1065661, 0.1428534, 0.1584353, 0.1406533, 0.1226292,
  0.1445243, 0.1545726, 0.1255022, 0.08527251, 0.07529252, 0.1570741, 
    0.1878532, 0.09091399, 0.09991471, 0.1797481, 0.1790022, 0.1420621, 
    0.06017789, 0.05908702, 0.1459581, 0.1638345, 0.2311812, 0.2936259, 
    0.3355277, 0.1096969, 0.1398648, 0.135156, 0.1496128, 0.1607532, 
    0.170334, 0.2747067, 0.1495072, 0.1886462, 0.2071912,
  0.1268812, 0.2012011, 0.1392934, 0.1525978, 0.1711459, 0.15973, 0.2114098, 
    0.1953841, 0.1696711, 0.1663709, 0.1883589, 0.1913684, 0.1250798, 
    0.2140096, 0.253071, 0.1703241, 0.235108, 0.2088194, 0.1862125, 
    0.1976585, 0.1748889, 0.1603085, 0.1265702, 0.1742431, 0.1288743, 
    0.1986677, 0.06195154, 0.1201416, 0.1207182,
  0.102147, 0.137795, 0.1659739, 0.1981845, 0.1887754, 0.1908862, 0.1491942, 
    0.09878998, 0.1302686, 0.1417583, 0.144904, 0.1271281, 0.09021419, 
    0.1128195, 0.115675, 0.1620933, 0.2326723, 0.2687944, 0.2863483, 
    0.2321388, 0.2519051, 0.3438681, 0.2314355, 0.1454409, 0.14521, 
    0.07865024, 0.1138152, 0.1023227, 0.1449046,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001799436, 0.0128057, 0.01034228, 
    0.00933532, -0.0002862941, 0.001269458, 7.890412e-05, 0.001449603, 
    -5.231797e-05, 0.003371444, 0.01362712, -0.0001076101, -3.748744e-10, 
    0.0007285339, -0.0004302296, 0,
  0.07162977, 0.04030817, 0.01772689, 0.01800392, -0.0006574473, 
    -0.0004776852, 0.007987594, 0, 0, -9.365026e-05, 0.001024009, 
    0.000729482, 0.001015045, 0.08806648, 0.1171118, 0.07892657, 0.08824035, 
    0.05072432, 0.03212797, 0.08550607, 0.07239144, 0.0793874, 0.08455093, 
    0.03042771, 0.0158127, 0.02367738, 0.03395574, 0.03032882, 0.1069617,
  0.1712406, 0.1884786, 0.1624165, 0.1558997, 0.1842764, 0.1702321, 
    0.1292107, 0.1066727, 0.0795626, 0.1000601, 0.114928, 0.1885117, 
    0.2419624, 0.2827087, 0.2381145, 0.2531826, 0.2902946, 0.3089127, 
    0.2161618, 0.1894322, 0.1591697, 0.1549802, 0.1332884, 0.1704474, 
    0.2635792, 0.1398603, 0.08632907, 0.1634435, 0.1725378,
  0.1860928, 0.1621898, 0.2709104, 0.1857636, 0.2228702, 0.1845163, 
    0.1623035, 0.1644168, 0.184971, 0.1855112, 0.2412766, 0.2334599, 
    0.1754842, 0.1574722, 0.1150096, 0.1910029, 0.1591818, 0.1570769, 
    0.1253235, 0.1116968, 0.185611, 0.2176929, 0.2458822, 0.1777485, 
    0.1858024, 0.1839159, 0.1997076, 0.210364, 0.2041084,
  0.1654272, 0.09225521, 0.08129415, 0.1355266, 0.0461178, 0.08312849, 
    0.09337474, 0.09877626, 0.06526222, 0.06117442, 0.06257648, 0.09613647, 
    0.06428276, 0.0926654, 0.1296632, 0.1222781, 0.05680185, 0.07430189, 
    0.103834, 0.1531168, 0.1762572, 0.1731362, 0.1801289, 0.1134622, 
    0.09686318, 0.09031353, 0.08052898, 0.09897292, 0.1655766,
  0.001058812, 0.0006707094, 0.003664174, 0.003985768, 0.05607901, 
    0.06319878, 0.01843318, 0.0007543781, 0.0001038884, 1.958866e-05, 
    5.964937e-07, 0.005435558, 0.01274551, 0.01758948, 0.04450521, 
    0.09464758, 0.1833073, 0.2424455, 0.1426039, 0.02012748, 0.02245681, 
    -0.0003190432, 3.203147e-05, 4.233596e-06, 0.02981356, 0.04393893, 
    0.0646824, 0.04765339, 0.01737149,
  9.213101e-09, 1.407436e-08, 5.798447e-07, 0.0001487687, 6.660502e-05, 
    0.01026213, 2.904413e-06, 0.006001037, 3.595926e-09, 0.0115017, 
    0.01896615, 0.003240274, 0.0003671399, -3.998871e-06, 0.06613611, 
    0.1012632, 0.05645439, 0.006636452, 0.0006822808, -1.898502e-09, 
    -6.365204e-11, 2.96021e-09, 1.041506e-08, 1.589267e-07, -8.239398e-05, 
    0.02202738, -6.191104e-05, 3.093899e-08, 3.175101e-08,
  7.02784e-08, 7.84934e-06, 3.989992e-09, 0, -1.008151e-07, 0.001085361, 
    0.08582573, 0.07361233, 0.03240933, 0.01699484, 0.004170999, 0.008400944, 
    0.0156376, 0.05585547, 0.01071467, 0.02120776, 0.0002258764, 
    1.266259e-10, 0, 1.243387e-08, 1.965145e-09, 2.289475e-08, 2.910809e-06, 
    0.001131613, 0.01252501, 0.000890343, 6.485858e-08, 2.917498e-09, 
    2.2357e-08,
  0.0003012415, 0.05801704, 0.02571464, 0.0004917164, 4.466785e-05, 
    0.05898765, 0.01139758, 0.02350813, 0.07048304, 0.1908719, 0.03651645, 
    0.1019041, 0.2399182, 0.04335141, 0.0228864, 0.007283413, 0.0002462178, 
    -1.729922e-05, 0.00311017, -5.57798e-05, 7.227006e-05, 0.01461005, 
    0.05706897, 0.02587972, 0.01075923, 0.001806811, 0.004434372, 
    -7.072609e-06, 3.305945e-06,
  0.2019075, 0.1482958, 0.07408375, 0.08380881, 0.02417377, 0.005197414, 
    0.03187495, 0.00654373, 0.0118336, 0.005268767, 0.00382173, 0.01325846, 
    0.06209654, 0.0405141, 0.05135964, 0.03932149, 0.06093659, 0.1451319, 
    0.1371982, 0.2289765, 0.1188889, 0.07311256, 0.1812506, 0.0564962, 
    0.02001216, 0.03446456, 0.05556928, 0.1595235, 0.2798659,
  6.003928e-05, 1.060504e-05, 7.743916e-07, 0.005040352, 0.03054437, 
    0.1454993, 0.1802717, 0.02090038, 0.1926671, 0.05612781, 0.0966886, 
    0.05918847, 0.0507524, 0.1099001, 0.04180097, 0.04870478, 0.009509766, 
    4.090642e-06, 0.001551719, 0.01064191, 0.02878202, 0.07993772, 
    0.01273887, 0.01240318, 0.006805297, 0.0008191365, 0.00535341, 
    0.000348129, 0.005946639,
  -1.962861e-05, 0.0006007634, 0, 0, 2.476229e-05, -5.366491e-05, 0.05042451, 
    0.1652818, 0.1966401, 0.02409424, 0.09926073, 0.05765029, 0.1693253, 
    0.08435694, 0.1233256, 0.0472253, 0.02590376, 0.01136232, -5.083079e-05, 
    0.03606799, 0.02086786, 0.01054188, 0.1015102, 0.02124282, 0.01149604, 
    0.01340787, 0.0004888545, -7.945798e-12, 0.003274761,
  0.02085904, 0.00171153, 0.004664184, 0.01338483, 0.0203114, 0.0115284, 
    0.07758157, 0.1346869, 0.1329095, 0.1155173, 0.1097036, 0.106127, 
    0.0424862, 0.1357251, 0.1388306, 0.1130834, 0.08828077, 0.05157277, 
    0.009960981, -8.038198e-05, 0.07741358, 0.01885184, 0.02874692, 
    0.03231518, 0.1005077, 0.04782296, 0.06183993, 0.02891446, 0.009256858,
  0.1431949, 0.1601147, 0.2098718, 0.07491256, 0.02697419, 0.06475917, 
    0.02153644, 0.04550003, 0.1707435, 0.1357649, 0.0633378, 0.1193339, 
    0.1006361, 0.1725885, 0.09593873, 0.09922243, 0.1061353, 0.1172133, 
    0.1992673, 0.0267479, 0.04594487, 0.07451351, 0.06077011, 0.06561487, 
    0.1090933, 0.1316832, 0.1479721, 0.1296142, 0.1342798,
  0.1342691, 0.132188, 0.1108546, 0.08368643, 0.06119545, 0.1609914, 
    0.1773577, 0.08315071, 0.08254956, 0.14637, 0.1580804, 0.1348382, 
    0.06287862, 0.06328337, 0.1371981, 0.1665766, 0.2184974, 0.290979, 
    0.3359351, 0.1143601, 0.1388383, 0.127339, 0.1563338, 0.1615815, 
    0.1660404, 0.2812089, 0.1505094, 0.1915263, 0.1853652,
  0.1087644, 0.1938175, 0.1357653, 0.1597863, 0.1700865, 0.1427202, 
    0.2056438, 0.1901794, 0.1544207, 0.1642298, 0.1959253, 0.1913959, 
    0.1328776, 0.2197287, 0.251227, 0.1623314, 0.2400279, 0.2127936, 
    0.178388, 0.1832069, 0.1735522, 0.167495, 0.1328852, 0.1801143, 
    0.1368645, 0.2380912, 0.1270901, 0.1179842, 0.113458,
  0.1027507, 0.1250752, 0.1520067, 0.1776017, 0.1720491, 0.1986331, 0.158751, 
    0.1046683, 0.145614, 0.1688675, 0.1779909, 0.1446738, 0.1240711, 0.15238, 
    0.1697334, 0.20682, 0.2499582, 0.2714207, 0.2867538, 0.2312132, 
    0.2443483, 0.3499393, 0.2199229, 0.1439791, 0.1373112, 0.09596201, 
    0.1277471, 0.09219852, 0.1340705,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.03332121, 0.1184072, 0.06843257, 
    0.02708741, 0.02831076, 0.002466685, 0.001056557, 0.003718227, 
    -0.0001029599, 0.006795402, 0.04456135, 0.01712619, -0.001054848, 
    0.01700797, 0.001876559, 0,
  0.1285457, 0.1023411, 0.06992848, 0.0336344, 0.0001279088, -0.0003496654, 
    0.0403861, -0.0003853344, -0.0002126315, -0.0005196201, 0.003455972, 
    0.0005928643, 0.01900156, 0.191209, 0.2720087, 0.1781342, 0.1603565, 
    0.1317966, 0.1014738, 0.1141452, 0.1368278, 0.2126581, 0.2305853, 
    0.129781, 0.109234, 0.1202965, 0.1616558, 0.1692626, 0.1757429,
  0.2365556, 0.2535794, 0.2206833, 0.2377189, 0.2362337, 0.2111986, 
    0.1690224, 0.1825833, 0.145473, 0.1994276, 0.2044309, 0.2546673, 
    0.3175204, 0.2914281, 0.2319584, 0.2405411, 0.289104, 0.2983037, 
    0.2263283, 0.255728, 0.2415948, 0.2761262, 0.2548287, 0.2380145, 
    0.3384202, 0.2217624, 0.1746603, 0.2020528, 0.2491726,
  0.1915738, 0.166275, 0.2622193, 0.1773296, 0.2087158, 0.1749095, 0.1607241, 
    0.1789225, 0.2024852, 0.1903051, 0.2599516, 0.2347578, 0.1777043, 
    0.1460726, 0.1304543, 0.1846882, 0.1376527, 0.165915, 0.1153729, 
    0.1193477, 0.1877159, 0.1952846, 0.2548242, 0.1895226, 0.1850451, 
    0.1896624, 0.2013567, 0.2198292, 0.2060748,
  0.156422, 0.09278309, 0.07984107, 0.1315152, 0.05044409, 0.07361719, 
    0.08749896, 0.09589904, 0.06047997, 0.05745699, 0.06946189, 0.09648982, 
    0.05718882, 0.08377025, 0.1298012, 0.1068119, 0.05850139, 0.08186298, 
    0.1011056, 0.1313044, 0.1742921, 0.1730019, 0.182771, 0.130916, 
    0.09628837, 0.08836496, 0.07981194, 0.1012122, 0.1449559,
  0.002566205, 0.0002297178, 0.01137084, 0.005931052, 0.054239, 0.06113814, 
    0.01412264, -0.0001155666, -5.070028e-05, -6.417094e-07, 1.461859e-05, 
    0.02766427, 0.01435086, 0.03183668, 0.05063938, 0.09306829, 0.183465, 
    0.2566057, 0.1542875, 0.02481067, 0.01821542, 0.002190336, 0.0002331793, 
    8.348526e-06, 0.03469757, 0.05143866, 0.06006831, 0.04461844, 0.01878879,
  4.622352e-08, 9.303853e-10, 4.410588e-07, 9.782142e-05, 0.007908602, 
    0.01372626, -0.0005002172, 0.000377414, 1.15317e-09, 0.01571669, 
    0.01588566, 0.001437109, 9.616751e-05, -3.595454e-05, 0.08500145, 
    0.08728958, 0.0546056, 0.0007120126, 0.0002924456, -1.032102e-09, 
    -1.029353e-09, 1.018124e-09, -1.191144e-10, 1.63404e-07, 0.0008652475, 
    0.03432064, -0.0002183658, 2.898725e-09, 8.688734e-09,
  3.846313e-08, 4.572717e-05, 1.373997e-07, 8.708621e-09, 1.790457e-06, 
    0.001268937, 0.07336453, 0.07127085, 0.04533052, 0.01992764, 0.002667482, 
    0.001937354, 0.02180749, 0.07290422, 0.009627135, 0.02596963, 
    0.000310622, 4.947714e-07, -2.28328e-09, 4.660976e-09, 1.540922e-09, 
    1.268564e-07, 1.24374e-06, 0.001593773, 0.007364663, 0.0003303463, 
    6.375486e-10, -1.797142e-11, -1.085738e-10,
  0.007076075, 0.04717007, 0.02405337, 0.002885543, 0.0001895075, 0.05384678, 
    0.008875756, 0.01975288, 0.06603106, 0.1982546, 0.02680321, 0.1012947, 
    0.2537824, 0.04401201, 0.02081874, 0.008801778, 0.00274194, 0.004263752, 
    0.004847189, 3.847068e-06, 0.001114954, 0.002144339, 0.05448474, 
    0.02008878, 0.01816271, 0.008770139, 0.002871604, 0.000487713, 
    0.0002769291,
  0.1918379, 0.1422478, 0.07884296, 0.09125938, 0.03435541, 0.01050243, 
    0.03177283, 0.006415821, 0.007585032, 0.004243419, 0.00381737, 
    0.009166666, 0.0567013, 0.03481212, 0.05107887, 0.03648127, 0.06176543, 
    0.1505156, 0.2006493, 0.241164, 0.1228752, 0.07473692, 0.1837123, 
    0.06155129, 0.01442597, 0.03609988, 0.06504381, 0.1546896, 0.2726784,
  2.407564e-05, 3.088258e-05, 1.30023e-06, 0.01476863, 0.02795191, 0.1150069, 
    0.1745123, 0.01853013, 0.1765424, 0.0562791, 0.1096622, 0.07016823, 
    0.04790654, 0.09103113, 0.03213925, 0.03828485, 0.005924825, 
    9.181412e-07, 0.01074436, 0.003603587, 0.02935685, 0.07796448, 
    0.01153414, 0.01145164, 0.005646443, 0.001103769, 0.003341827, 
    0.001143678, 0.002189261,
  0.0003400126, 0.0005893063, 0, -9.202081e-12, 0.002005395, -9.400792e-05, 
    0.05310802, 0.1737932, 0.1944852, 0.02170485, 0.08731809, 0.06461789, 
    0.1803318, 0.07950541, 0.1220507, 0.03912338, 0.02778197, 0.004460567, 
    0.001047889, 0.02700902, 0.01790538, 0.009295228, 0.07989172, 0.01569335, 
    0.007018531, 0.006766085, 0.0005245837, -6.595894e-10, 0.03239554,
  0.01810617, 0.003138228, 0.003774496, 0.01492893, 0.02297018, 0.005569462, 
    0.08830569, 0.1211449, 0.1206424, 0.1076058, 0.1068299, 0.08682351, 
    0.04420445, 0.122929, 0.1325039, 0.09957206, 0.1209214, 0.06601947, 
    0.0142958, -0.000106939, 0.1053626, 0.0164126, 0.03049696, 0.02704195, 
    0.09483238, 0.04456904, 0.05932554, 0.03223852, 0.004671313,
  0.1173427, 0.1551363, 0.2025681, 0.06540856, 0.03026966, 0.05767735, 
    0.01373123, 0.0434647, 0.1677216, 0.1336309, 0.05506882, 0.09298462, 
    0.08235466, 0.1640914, 0.09700636, 0.09615269, 0.1054811, 0.1203556, 
    0.2068833, 0.01965287, 0.04935798, 0.08137714, 0.06134, 0.08270053, 
    0.1071002, 0.124927, 0.1371018, 0.1324867, 0.1135508,
  0.1464902, 0.1304628, 0.09535763, 0.07851053, 0.04454798, 0.1373561, 
    0.1618258, 0.07260823, 0.08203655, 0.1188205, 0.1513343, 0.1374413, 
    0.06417658, 0.07327573, 0.1314939, 0.1507186, 0.2022548, 0.2680443, 
    0.3408399, 0.1093605, 0.1415598, 0.1102128, 0.1463336, 0.1766636, 
    0.1581092, 0.2780216, 0.1335924, 0.202264, 0.2013936,
  0.1103399, 0.2184615, 0.1414735, 0.1836568, 0.1812464, 0.154319, 0.2303817, 
    0.2145239, 0.153956, 0.178456, 0.1896828, 0.2068586, 0.1710266, 
    0.2285627, 0.2647161, 0.1457676, 0.2323886, 0.234037, 0.1703846, 
    0.1834315, 0.1624309, 0.1475297, 0.1313817, 0.1777305, 0.1183693, 
    0.2224576, 0.1275457, 0.1346667, 0.1011318,
  0.1094159, 0.1178132, 0.1445477, 0.1827884, 0.1635803, 0.2143556, 
    0.1584407, 0.1189652, 0.1429236, 0.176653, 0.2079305, 0.1699072, 
    0.194417, 0.2477104, 0.2482799, 0.2703875, 0.2753343, 0.2811076, 
    0.294699, 0.2342487, 0.2488222, 0.3403764, 0.2107281, 0.1287469, 
    0.1346617, 0.1039385, 0.1190189, 0.08450733, 0.1265623,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.148971, 0.1723804, 0.0844778, 
    0.04964517, 0.05292442, 0.05463426, 0.006399156, 0.004462239, 
    0.0001089079, 0.01510676, 0.1061639, 0.1162736, 0.06940673, 0.1229824, 
    0.02267737, 0,
  0.1585617, 0.1996179, 0.150939, 0.1066768, 0.006085228, 0.004065847, 
    0.0827236, -0.001946322, 0.0004515365, -0.0008931037, 0.008094128, 
    0.002495418, 0.06202308, 0.2920738, 0.3082966, 0.2151535, 0.2021408, 
    0.1614096, 0.1734288, 0.2022113, 0.2383447, 0.294945, 0.2989367, 
    0.2777916, 0.2058662, 0.2159697, 0.2718331, 0.2383337, 0.2046002,
  0.264072, 0.27091, 0.2615291, 0.296027, 0.2597614, 0.2427839, 0.2270873, 
    0.2527595, 0.2080368, 0.2662989, 0.2559929, 0.3237484, 0.3163439, 
    0.2634869, 0.2108353, 0.2307135, 0.2691549, 0.2946722, 0.2330071, 
    0.2561299, 0.2537715, 0.2828852, 0.2580715, 0.2377197, 0.3370475, 
    0.22607, 0.1774762, 0.2487735, 0.3067431,
  0.184648, 0.1746886, 0.233007, 0.1639636, 0.189186, 0.1665909, 0.1538823, 
    0.1984403, 0.2032695, 0.2173854, 0.2698255, 0.2333178, 0.1649715, 
    0.1259935, 0.1364912, 0.1765081, 0.1334372, 0.1702183, 0.1226313, 
    0.1052057, 0.1668134, 0.1848304, 0.2486989, 0.1862321, 0.1717681, 
    0.181191, 0.2054214, 0.2201177, 0.2127713,
  0.1449547, 0.08670107, 0.07052939, 0.1253004, 0.05289426, 0.06821783, 
    0.0970152, 0.08726713, 0.05315667, 0.05983989, 0.06061874, 0.08962691, 
    0.06177117, 0.09237883, 0.1477444, 0.1318981, 0.06820136, 0.07604346, 
    0.09815227, 0.129091, 0.1586607, 0.1586953, 0.1534029, 0.1280171, 
    0.0964584, 0.1034053, 0.06967869, 0.1016511, 0.1437422,
  0.003290896, 4.320557e-05, 0.02936066, 0.008194701, 0.05525963, 0.0737804, 
    0.01762158, 0.002267953, -5.886091e-05, 7.459972e-05, 0.001695437, 
    0.05299119, 0.01937605, 0.04506058, 0.04038374, 0.08350358, 0.1815071, 
    0.2589796, 0.1634376, 0.02117102, 0.03691405, 0.01148763, 0.0001964653, 
    1.424666e-05, 0.05414817, 0.05852062, 0.0598763, 0.0376269, 0.02218452,
  2.693287e-08, -3.648364e-10, -8.11738e-07, 7.379237e-05, 0.01960601, 
    0.01575286, 0.001487972, 9.952015e-05, 2.804529e-08, 0.01261066, 
    0.008846251, 5.713696e-05, 0.0009772746, 0.007540926, 0.1079545, 
    0.1013173, 0.06048173, 0.001214606, 0.0001109738, -2.814335e-09, 
    -4.699114e-09, 8.537145e-09, 1.027088e-08, 6.182452e-07, 0.009273938, 
    0.04193022, -0.0004391281, 1.811142e-08, 2.596306e-08,
  1.192501e-07, 0.0001102299, 2.265121e-06, -4.483883e-09, 0.0001137155, 
    0.002024712, 0.07394102, 0.07436448, 0.04486448, 0.00449447, 0.0063156, 
    0.003867676, 0.02271436, 0.0821979, 0.008720819, 0.03282437, 
    0.0007402104, 2.566766e-05, 3.48558e-09, 2.396052e-08, 5.555785e-09, 
    9.903503e-08, 1.274948e-06, 0.002131574, 0.007279629, 0.0002499377, 
    5.148746e-08, 5.364268e-09, 6.464028e-09,
  0.0225779, 0.04125771, 0.02344686, 0.002160335, 0.0002592293, 0.05552921, 
    0.007939728, 0.01638241, 0.07004687, 0.2215734, 0.03041135, 0.1157363, 
    0.2664486, 0.04932443, 0.0253718, 0.01129541, 0.005592544, 0.01552194, 
    0.01069459, 0.0002359795, 0.01212436, 0.003290463, 0.06766852, 
    0.02336396, 0.01756674, 0.01226823, 0.01706595, 0.001869443, 0.00558988,
  0.1993213, 0.1356051, 0.09051392, 0.1088846, 0.02811904, 0.02775593, 
    0.03076852, 0.007429131, 0.01050447, 0.004121846, 0.002575216, 
    0.007162859, 0.04881537, 0.03793453, 0.05365534, 0.04678784, 0.07854223, 
    0.1569092, 0.2521367, 0.2592848, 0.1182316, 0.07687962, 0.2018695, 
    0.06680444, 0.01227003, 0.04084848, 0.0735564, 0.164501, 0.2758689,
  0.002239454, 3.25607e-05, -1.328556e-05, 0.002204745, 0.01150718, 
    0.09027348, 0.2044076, 0.03657098, 0.1774973, 0.07313138, 0.152161, 
    0.1029807, 0.05424627, 0.08088055, 0.0301155, 0.0359362, 1.407987e-05, 
    2.747426e-06, 0.0035779, 0.0103283, 0.03697167, 0.07717077, 0.01395301, 
    0.01512799, 0.006106806, 0.0008082257, 0.002534497, 0.001036137, 
    0.004112058,
  -0.0004266017, 0.01119082, 0, -1.332062e-11, 0.00573378, 0.0003793002, 
    0.06455317, 0.1848076, 0.225514, 0.03186192, 0.08696292, 0.07239054, 
    0.1867122, 0.08662678, 0.1406523, 0.03451791, 0.0128438, 0.0002550861, 
    1.51563e-05, 0.01919628, 0.02512703, 0.01270712, 0.07190578, 0.01227123, 
    0.004651154, 0.003169832, 0.0007871779, 4.194794e-08, 0.04475814,
  0.0134096, 0.005941547, 0.001942881, 0.01953242, 0.02007136, 0.001474832, 
    0.1023602, 0.09978273, 0.1036263, 0.102036, 0.1089995, 0.0827749, 
    0.05346826, 0.1095153, 0.1345729, 0.08806422, 0.071558, 0.03795286, 
    0.008228343, -6.770476e-05, 0.1199546, 0.01646766, 0.03798514, 
    0.03320251, 0.09184647, 0.03321362, 0.06431331, 0.02433188, 0.004028275,
  0.1008783, 0.1784484, 0.1887423, 0.07333343, 0.03425134, 0.04531281, 
    0.01322211, 0.05252404, 0.1546327, 0.1438557, 0.05127169, 0.07647124, 
    0.09607302, 0.1604148, 0.09776656, 0.07808381, 0.1142307, 0.1054864, 
    0.183827, 0.02123361, 0.04685071, 0.07837029, 0.06147223, 0.06548888, 
    0.09959923, 0.1389034, 0.1134852, 0.1083301, 0.1002825,
  0.122901, 0.1149465, 0.1013807, 0.08619386, 0.03444915, 0.1224464, 
    0.1647511, 0.08971696, 0.07168194, 0.109888, 0.1353974, 0.1546288, 
    0.06377257, 0.08936106, 0.125874, 0.1422978, 0.1851797, 0.2850612, 
    0.3601667, 0.09690278, 0.1390927, 0.1111049, 0.1641465, 0.1721874, 
    0.1580092, 0.2671201, 0.1390707, 0.2545918, 0.159638,
  0.1149071, 0.2151822, 0.1355181, 0.1872034, 0.2259028, 0.1526843, 0.210703, 
    0.2036107, 0.1728325, 0.1814529, 0.1838448, 0.2297032, 0.2034767, 
    0.2098072, 0.2756321, 0.1521771, 0.2157078, 0.200083, 0.2003235, 
    0.177327, 0.1512628, 0.1314928, 0.1390285, 0.1874608, 0.122978, 0.215628, 
    0.1161963, 0.1393342, 0.07653743,
  0.1080503, 0.1593662, 0.1398835, 0.1926668, 0.2234242, 0.2362394, 
    0.1476749, 0.1284079, 0.1878278, 0.2076762, 0.2604854, 0.2098755, 
    0.2283393, 0.3154088, 0.3406235, 0.3110034, 0.2734166, 0.2832541, 
    0.3034379, 0.2825605, 0.3045405, 0.3995381, 0.1988769, 0.1285304, 
    0.1433531, 0.1189709, 0.1201948, 0.08974492, 0.1289875,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0002184165, -0.0002184165, 
    -0.0002184165, -0.0002184165, -0.0002184165, -0.0002184165, 
    -0.0002184165, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.000329046, 0.2129536, 0.1923478, 
    0.09337036, 0.08720624, 0.09404679, 0.06784976, 0.08880296, 0.03416189, 
    0.01296637, 0.05308892, 0.2048258, 0.2265832, 0.1677098, 0.2370286, 
    0.1022976, 0,
  0.1772096, 0.2725687, 0.1962801, 0.1812821, 0.02393849, 0.006294556, 
    0.1153177, 0.006358207, 0.007573265, -0.002357541, 0.02591716, 
    0.02095005, 0.1725722, 0.3174548, 0.3458972, 0.2410218, 0.2302627, 
    0.1994517, 0.2230504, 0.2648659, 0.3108827, 0.3278148, 0.3074995, 
    0.3703009, 0.2411116, 0.2198112, 0.2610749, 0.2604663, 0.2067319,
  0.2566402, 0.2532483, 0.2654736, 0.2956732, 0.2701927, 0.2566589, 
    0.2900196, 0.271694, 0.2445098, 0.3101892, 0.2657489, 0.3137599, 
    0.3056298, 0.2608719, 0.2104309, 0.2216998, 0.2736428, 0.2767826, 
    0.2326957, 0.2842404, 0.2554828, 0.2725568, 0.2491923, 0.2325344, 
    0.3139546, 0.2082316, 0.1843011, 0.2430882, 0.3205389,
  0.1862206, 0.1664178, 0.2104921, 0.1655962, 0.1807467, 0.1535147, 
    0.1572067, 0.1955332, 0.2102273, 0.220963, 0.2599374, 0.2398503, 
    0.1598797, 0.1310438, 0.1347215, 0.2038045, 0.126049, 0.1535946, 
    0.1392977, 0.1161109, 0.1517104, 0.1546362, 0.2218275, 0.1792725, 
    0.1718506, 0.1795, 0.20161, 0.2296646, 0.2060321,
  0.1421602, 0.08505967, 0.07018039, 0.1236594, 0.05165741, 0.07673968, 
    0.100628, 0.0944709, 0.05562678, 0.05296902, 0.06184258, 0.08453323, 
    0.06427191, 0.07989507, 0.1618239, 0.1303, 0.07252102, 0.07428823, 
    0.1069442, 0.1216091, 0.1713412, 0.1490042, 0.1654428, 0.1348737, 
    0.09435288, 0.08408833, 0.06973612, 0.1050884, 0.1458558,
  0.0046522, 0.0003971857, 0.04832483, 0.01646738, 0.06518964, 0.0826491, 
    0.01488283, 0.005122272, -4.588209e-06, 0.005083308, 0.01214343, 
    0.04691598, 0.02865241, 0.04840695, 0.05697918, 0.0828338, 0.1759575, 
    0.2631985, 0.1498513, 0.02206196, 0.05673191, 0.02687227, 0.001173616, 
    -1.700273e-06, 0.08215422, 0.06536276, 0.05994945, 0.03815705, 0.03091518,
  1.936595e-07, 5.763031e-07, 6.90442e-05, 0.002441898, 0.03498096, 
    0.02476786, -6.300078e-06, 0.002250423, 2.380577e-07, 0.02335301, 
    0.006202775, 1.551349e-05, 0.0009360298, 0.0175969, 0.1017973, 0.1279226, 
    0.05949312, 0.002187604, 0.0002596076, 1.489093e-08, -2.897138e-09, 
    1.007608e-08, 1.163423e-08, 8.580383e-07, 0.01769544, 0.04440985, 
    0.001023586, 2.019039e-07, 3.274704e-07,
  3.313655e-07, 0.0003470655, 1.493802e-05, 1.856824e-07, 0.000353559, 
    0.005207425, 0.07412995, 0.07536116, 0.05111014, 0.00454722, 0.01677149, 
    0.01015002, 0.03160698, 0.08479371, 0.01219627, 0.03655833, 0.003344264, 
    0.0001062291, 1.557799e-07, 9.549886e-08, 4.172429e-08, 4.816717e-07, 
    7.80351e-06, 0.003513414, 0.004206622, 0.0006270029, 3.098592e-07, 
    1.411893e-08, 3.170489e-08,
  0.01594242, 0.05046386, 0.0355876, 0.0003476429, 0.001108292, 0.06360543, 
    0.0110988, 0.02060058, 0.08527476, 0.2604413, 0.04830448, 0.1423126, 
    0.2763498, 0.06598231, 0.0264664, 0.01362218, 0.01177674, 0.01419849, 
    0.01009755, 0.002664812, 0.004365679, 0.005426765, 0.07342478, 
    0.03262766, 0.01886319, 0.01281763, 0.03719407, 0.001448029, 0.002454942,
  0.220657, 0.1681486, 0.1211062, 0.1344786, 0.01742675, 0.02113422, 
    0.03302165, 0.01555095, 0.05680561, 0.00607933, 0.005344774, 0.01187362, 
    0.04913627, 0.04912741, 0.07618664, 0.06885974, 0.09614886, 0.2209015, 
    0.2771264, 0.2890266, 0.1165573, 0.1030231, 0.1951872, 0.09343497, 
    0.01775526, 0.05558961, 0.08523013, 0.2057765, 0.3216655,
  0.05614682, -0.0001302982, 1.250034e-05, 0.0001587928, 0.00245584, 
    0.05616578, 0.2338826, 0.07796928, 0.1995174, 0.08770504, 0.1880615, 
    0.1210585, 0.0653962, 0.09708407, 0.04135475, 0.03892607, 1.941244e-05, 
    3.524099e-06, 0.002033825, 0.02885109, 0.0414198, 0.08729257, 0.0193154, 
    0.0231895, 0.007922133, 0.006483898, 0.001306687, 0.0008616832, 
    0.004845237,
  -0.0001824685, 0.04995241, 0, -3.617539e-09, 0.005573206, -5.694925e-05, 
    0.07807709, 0.1915452, 0.2598146, 0.03351199, 0.09798802, 0.09136872, 
    0.2082858, 0.108398, 0.1497718, 0.02993887, 0.001961404, 0.0009050499, 
    9.918665e-07, 0.01054638, 0.04463582, 0.01824106, 0.07316072, 
    0.009767302, 0.004847555, 0.003135684, 0.0008898673, 5.352195e-08, 
    0.03388645,
  0.009963163, 0.005229265, 0.001755383, 0.02968028, 0.01770554, 0.001189907, 
    0.1235575, 0.09477618, 0.08694284, 0.1027018, 0.1172586, 0.0786114, 
    0.06384235, 0.106974, 0.1368401, 0.08048648, 0.08455185, 0.04510382, 
    0.01182851, -7.2635e-05, 0.09411594, 0.01904566, 0.0422951, 0.04127898, 
    0.09777245, 0.03563714, 0.06393952, 0.02465036, 0.001862329,
  0.1021129, 0.1748753, 0.1786429, 0.07726902, 0.03567365, 0.03944108, 
    0.01394057, 0.0565459, 0.1502364, 0.1570275, 0.05535926, 0.07122451, 
    0.09906018, 0.1658857, 0.08544809, 0.08245979, 0.1120788, 0.09707317, 
    0.1903017, 0.0219964, 0.04589775, 0.06639305, 0.06408403, 0.07243361, 
    0.1032017, 0.1309505, 0.1105141, 0.09920812, 0.1050836,
  0.1587307, 0.1137068, 0.09370786, 0.06102275, 0.02880508, 0.1124847, 
    0.1527149, 0.07466891, 0.08492455, 0.1276306, 0.1260496, 0.1684951, 
    0.07523159, 0.1084293, 0.1113658, 0.1467687, 0.1625641, 0.2713028, 
    0.3834881, 0.09848092, 0.1354718, 0.1241507, 0.1788931, 0.2138523, 
    0.1408227, 0.2648535, 0.129474, 0.2027082, 0.1651887,
  0.08096766, 0.1821791, 0.1384882, 0.1375991, 0.2476511, 0.2459314, 
    0.2557574, 0.2824835, 0.1722981, 0.2135429, 0.2202012, 0.2446899, 
    0.1890876, 0.2155417, 0.2583182, 0.1367757, 0.2469265, 0.2046727, 
    0.2245157, 0.2277844, 0.1756578, 0.1261362, 0.09775919, 0.2044684, 
    0.08229116, 0.2198328, 0.1030865, 0.1130312, 0.06967379,
  0.09705459, 0.1043163, 0.1296965, 0.1726283, 0.1848672, 0.2288369, 
    0.1748897, 0.1360137, 0.1750373, 0.2509806, 0.2884136, 0.2421738, 
    0.3051139, 0.401428, 0.4315405, 0.34074, 0.3213944, 0.2896287, 0.3264412, 
    0.2520624, 0.2360172, 0.3842484, 0.2136743, 0.1570953, 0.1645259, 
    0.1328462, 0.1589917, 0.07490317, 0.1080063,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0001670188, -0.0001670188, 
    -0.0001670188, -0.0001670188, -0.0001670188, -0.0001670188, 
    -0.0001670188, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.148176e-05, 0.002504447, 0.2343522, 
    0.1838798, 0.1255063, 0.1170021, 0.1369257, 0.08608368, 0.1288853, 
    0.08379475, 0.04867915, 0.09972566, 0.2095856, 0.2410965, 0.2382757, 
    0.2630099, 0.2449595, 0.002407756,
  0.1959556, 0.2814604, 0.2361202, 0.2341946, 0.03313804, 0.02033828, 
    0.1218871, 0.03509638, 0.02692407, 0.001678401, 0.03936908, 0.03971129, 
    0.2407241, 0.3291289, 0.3468599, 0.2710558, 0.231278, 0.2177932, 
    0.2669403, 0.2679822, 0.2962787, 0.2898545, 0.2802764, 0.3468411, 
    0.2347263, 0.2207033, 0.2438442, 0.2658792, 0.2065719,
  0.2456109, 0.2322178, 0.2427163, 0.3063661, 0.2766862, 0.2588653, 
    0.2583431, 0.2654684, 0.2468661, 0.3246558, 0.2543921, 0.2879704, 
    0.2901698, 0.2591426, 0.204387, 0.2117072, 0.2582948, 0.274621, 
    0.2298606, 0.3103043, 0.2669111, 0.2632999, 0.2464765, 0.2259177, 
    0.3059664, 0.1905009, 0.1813665, 0.2389175, 0.2942219,
  0.1756718, 0.1678003, 0.1915028, 0.1668388, 0.1920383, 0.1736648, 
    0.1667949, 0.212017, 0.1991179, 0.216426, 0.2692955, 0.2437715, 
    0.1631598, 0.1512443, 0.1088323, 0.201808, 0.1257313, 0.1519099, 
    0.1363005, 0.1219786, 0.1396808, 0.1617906, 0.2129155, 0.1720813, 
    0.1501444, 0.1682762, 0.1873401, 0.2215711, 0.1910979,
  0.1216529, 0.09276605, 0.07791242, 0.1189493, 0.05352139, 0.09099266, 
    0.1058259, 0.09178753, 0.05164352, 0.06060576, 0.07395516, 0.1018175, 
    0.0661223, 0.07917428, 0.1677365, 0.1047783, 0.07023484, 0.08808498, 
    0.1128188, 0.112099, 0.1683655, 0.1375997, 0.1512572, 0.1404993, 
    0.09563268, 0.0780274, 0.06886619, 0.1171216, 0.1646253,
  0.004675225, 0.0007059926, 0.0976492, 0.02125506, 0.06630783, 0.09891132, 
    0.01469331, 0.006449348, 0.0002139229, 0.01915477, 0.04076758, 
    0.04303004, 0.03946501, 0.04551617, 0.07402845, 0.09377173, 0.1717429, 
    0.2510169, 0.1370598, 0.03262161, 0.07190171, 0.04300968, 0.0005963101, 
    3.1582e-05, 0.1236417, 0.06797385, 0.06300046, 0.04734609, 0.03309517,
  1.33277e-07, 0.0001161136, 0.01089834, 0.002099839, 0.06713707, 0.02887057, 
    0.006353778, -3.632794e-05, 8.400121e-07, 0.02056067, 0.02561714, 
    0.0003700716, 0.0002913242, 0.01796524, 0.09807409, 0.1538672, 
    0.06088091, 0.002281342, 0.0002823873, -7.745928e-07, 1.238181e-07, 
    1.340044e-08, 6.438679e-09, 6.387759e-07, 0.03383163, 0.05019935, 
    0.003919306, 9.574309e-07, 2.741106e-07,
  9.531869e-07, 0.000704067, 0.0003378065, 4.810327e-06, 0.0002698327, 
    0.006911333, 0.0827068, 0.08614575, 0.07242405, 0.007108492, 0.01908377, 
    0.01207874, 0.05108699, 0.1065795, 0.01828383, 0.03774212, 0.002885346, 
    0.0001979884, 5.176737e-05, 1.023853e-07, 8.497705e-08, 5.256434e-07, 
    1.168329e-05, 0.00494309, 0.01345062, 0.005320703, 6.210896e-07, 
    1.411499e-08, 4.594831e-08,
  0.02134822, 0.08167255, 0.08738215, 0.003742858, 0.00690283, 0.06621223, 
    0.01605383, 0.03668861, 0.1228134, 0.3040658, 0.05724259, 0.1729073, 
    0.2894128, 0.07642758, 0.02897691, 0.01404558, 0.01302119, 0.006267443, 
    0.001848478, 0.0003151107, 0.002829668, 0.0009334999, 0.0553826, 
    0.06164963, 0.02569892, 0.01226053, 0.02144322, 0.009813128, 0.009938656,
  0.2647916, 0.2161408, 0.1537642, 0.1709045, 0.01170532, 0.006962708, 
    0.03917708, 0.02613463, 0.0957368, 0.008175506, 0.008983514, 0.01763143, 
    0.05872708, 0.06501268, 0.1028531, 0.08287607, 0.1165, 0.2607126, 
    0.2936789, 0.3238685, 0.1153533, 0.1085002, 0.207891, 0.1202844, 
    0.02277901, 0.06714176, 0.1055506, 0.2263035, 0.3577533,
  0.0217597, 0.0047308, 4.634447e-06, -5.613597e-06, 0.0002671, 0.01666293, 
    0.2712616, 0.08303659, 0.2250051, 0.08190636, 0.1611021, 0.1059978, 
    0.06876073, 0.1184014, 0.05947861, 0.04194029, 1.977695e-05, 
    7.610231e-05, 0.002083501, 0.02093498, 0.0643972, 0.1007309, 0.01920754, 
    0.02392983, 0.007081036, 0.001717165, 6.472149e-05, 0.0001357844, 
    0.001471903,
  -2.895272e-05, 0.02261201, -1.53828e-10, -3.003627e-11, 0.001801495, 
    -5.01033e-06, 0.06908689, 0.2251243, 0.2682154, 0.02303511, 0.1034731, 
    0.08905857, 0.234331, 0.1251431, 0.1662497, 0.02442136, 0.0006233018, 
    0.01399175, 1.020384e-06, 0.0006100895, 0.0604896, 0.02941585, 
    0.08025146, 0.01346823, 0.005791132, 0.00512385, 0.002301139, 
    5.295858e-08, 0.01177699,
  0.002340052, 0.005169933, 0.002024582, 0.03067187, 0.0147644, 0.002408395, 
    0.1210119, 0.09286348, 0.07016061, 0.1237273, 0.1316101, 0.08699906, 
    0.07394959, 0.1145194, 0.143636, 0.07175412, 0.07678182, 0.04622241, 
    0.00849981, -1.813143e-05, 0.04640864, 0.01995973, 0.05054097, 
    0.05802848, 0.1188425, 0.03960051, 0.07404557, 0.02438748, 0.001509276,
  0.100348, 0.1647398, 0.172778, 0.07505704, 0.05057833, 0.04125058, 
    0.0201224, 0.06407105, 0.154298, 0.1644613, 0.07566036, 0.07840728, 
    0.1097985, 0.1904761, 0.07713969, 0.07784033, 0.1281548, 0.111064, 
    0.1871206, 0.01902357, 0.02817464, 0.04160703, 0.06926506, 0.07064765, 
    0.1294326, 0.1316092, 0.09982682, 0.107371, 0.1056817,
  0.1356555, 0.1174416, 0.07796751, 0.05431288, 0.03600658, 0.121217, 
    0.1715493, 0.09489044, 0.0821399, 0.1423656, 0.1289969, 0.1918793, 
    0.08150642, 0.12525, 0.1135549, 0.1360149, 0.1465434, 0.2962814, 
    0.3971812, 0.08754697, 0.1292831, 0.1239002, 0.1849556, 0.1886857, 
    0.1395286, 0.2746847, 0.1204483, 0.1965774, 0.146376,
  0.07758893, 0.1674169, 0.1307278, 0.1901844, 0.2479842, 0.2219758, 
    0.2576509, 0.2358023, 0.2401969, 0.2368497, 0.2362338, 0.2174655, 
    0.1840633, 0.2570826, 0.2911806, 0.1597922, 0.2390047, 0.1660844, 
    0.2187709, 0.2262632, 0.1738712, 0.1196521, 0.08705808, 0.1976111, 
    0.06355403, 0.2603256, 0.1016704, 0.1200937, 0.0604194,
  0.1087244, 0.1294631, 0.1451127, 0.1674932, 0.1989048, 0.2148539, 0.212803, 
    0.1976785, 0.2448592, 0.2754918, 0.3584361, 0.3963245, 0.3593581, 
    0.4691282, 0.4784584, 0.3768457, 0.4057131, 0.3230228, 0.4025375, 
    0.3437754, 0.2497068, 0.3658606, 0.2240963, 0.1614741, 0.1600989, 
    0.1605865, 0.1653033, 0.06630258, 0.1341195,
  0.0001481954, 9.430615e-05, 4.041692e-05, -1.347231e-05, -6.736154e-05, 
    -0.0001212508, -0.00017514, -0.0001166826, -8.405105e-05, -5.141949e-05, 
    -1.878793e-05, 1.384363e-05, 4.647519e-05, 7.910676e-05, -0.002677071, 
    -0.002143893, -0.001610715, -0.001077537, -0.0005443587, -1.118071e-05, 
    0.0005219973, 0.0002520553, -0.000259865, -0.0007717854, -0.001283706, 
    -0.001795626, -0.002307547, -0.002819467, 0.0001913068,
  -0.003089417, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0001792608, 0.01183662, 
    0.2248425, 0.16538, 0.1162691, 0.1344704, 0.1723982, 0.1551976, 
    0.1948744, 0.1309487, 0.08787776, 0.1454271, 0.2381978, 0.2148647, 
    0.2304648, 0.250213, 0.3014946, 0.04920447,
  0.2064344, 0.297418, 0.2427551, 0.2730003, 0.06503031, 0.04559088, 
    0.1334064, 0.07353593, 0.03700501, 0.04190014, 0.07745418, 0.07149008, 
    0.249857, 0.3393807, 0.3688274, 0.2900759, 0.2674015, 0.26098, 0.266156, 
    0.2699402, 0.2871666, 0.2986041, 0.2924348, 0.3825919, 0.2567449, 
    0.213374, 0.2484211, 0.2784143, 0.2077834,
  0.2232786, 0.2165785, 0.237638, 0.2966751, 0.2689331, 0.2483527, 0.2645259, 
    0.2751789, 0.254752, 0.3218017, 0.2494708, 0.2729007, 0.2961382, 
    0.2641538, 0.2372132, 0.228001, 0.2524228, 0.2647915, 0.2608022, 
    0.3146457, 0.2641091, 0.2882946, 0.2365681, 0.220946, 0.3215731, 
    0.1858401, 0.1789914, 0.2198733, 0.2934299,
  0.1825939, 0.1678706, 0.1801444, 0.1591626, 0.1742828, 0.1785682, 
    0.1692953, 0.2156847, 0.2091709, 0.2372607, 0.2841749, 0.244877, 
    0.1757619, 0.156679, 0.1309315, 0.1974766, 0.1309726, 0.1505752, 
    0.1202474, 0.1317302, 0.1349607, 0.1555713, 0.2021672, 0.1634465, 
    0.1419759, 0.1629848, 0.1866782, 0.2202821, 0.1783671,
  0.1129636, 0.1007411, 0.0829639, 0.1222516, 0.0626384, 0.08813762, 
    0.1017029, 0.08441031, 0.04743067, 0.07127733, 0.08785231, 0.11327, 
    0.07396055, 0.08686908, 0.1628536, 0.1044475, 0.06783247, 0.094438, 
    0.1102975, 0.1050748, 0.1522174, 0.1389049, 0.1493718, 0.1416084, 
    0.09813033, 0.06590605, 0.06294136, 0.127766, 0.1851619,
  0.007001288, 0.0004757864, 0.1194311, 0.02653174, 0.07243592, 0.1160794, 
    0.01747244, 0.00712283, 0.0007273075, 0.01383421, 0.06385473, 0.0179517, 
    0.052201, 0.05116264, 0.07529523, 0.111224, 0.1742257, 0.2374422, 
    0.1345771, 0.04849359, 0.08132993, 0.0546636, 0.001158706, 2.936478e-05, 
    0.1686715, 0.08183621, 0.06924062, 0.04996916, 0.03403005,
  7.435116e-08, 8.245873e-07, 0.00274327, 0.002653682, 0.07569665, 
    0.02819296, 0.01683499, 1.06647e-06, 1.711038e-06, 0.009333105, 
    0.0491425, 0.008559504, 0.01293153, 0.01741203, 0.08272031, 0.1548764, 
    0.07944312, 0.004254733, 0.001170826, 2.337309e-05, 1.367859e-06, 
    1.045361e-08, 2.319408e-09, 3.351648e-07, 0.02585406, 0.05641126, 
    0.006566081, 7.051314e-07, 2.324463e-07,
  1.041039e-06, -0.0005326149, 0.001984445, 0.001235006, 0.0001405347, 
    0.01107448, 0.08901377, 0.08234976, 0.07619111, 0.01272988, 0.01782849, 
    0.009858967, 0.06156725, 0.09450504, 0.0206498, 0.04265875, 0.002684022, 
    0.001331733, 8.162761e-05, 5.177841e-08, 1.69826e-07, 5.73369e-07, 
    1.156957e-05, 0.005641128, 0.06828885, 0.0237799, 1.629474e-05, 
    3.386327e-08, 7.645097e-08,
  0.02337515, 0.1060373, 0.1262329, 0.00950312, 0.0003085119, 0.06377791, 
    0.01812364, 0.03119071, 0.1312058, 0.3405593, 0.04172318, 0.1375129, 
    0.2657026, 0.06123183, 0.02875295, 0.01075443, 0.01868913, 0.01093663, 
    0.0130403, 0.0009210171, 0.0001822606, 0.002429501, 0.033172, 0.0928821, 
    0.03513609, 0.01441291, 0.01242156, 0.002491161, 0.02263244,
  0.2428165, 0.2371627, 0.1414709, 0.2226823, 0.007655095, 0.003804051, 
    0.03390775, 0.02654903, 0.05827156, 0.007889352, 0.007660507, 0.01370642, 
    0.04334294, 0.0495893, 0.08985928, 0.07476365, 0.1226222, 0.2865471, 
    0.2851428, 0.3187235, 0.09339352, 0.08576334, 0.2149674, 0.1205572, 
    0.02121167, 0.06443643, 0.0972164, 0.184268, 0.3917011,
  0.002272601, 0.0004260011, 3.287333e-06, 2.595935e-06, 1.853465e-05, 
    0.002490138, 0.1732959, 0.07635338, 0.2378861, 0.07047746, 0.110158, 
    0.08121711, 0.04198916, 0.07907154, 0.03994776, 0.03558296, 1.131151e-05, 
    2.114931e-05, 0.0001548851, 0.01214585, 0.05069278, 0.100297, 0.01431288, 
    0.0185606, 0.005809331, 0.001083698, 0.0001292573, 0.0001193923, 
    0.001071542,
  -1.324629e-06, 0.002617309, 6.869132e-10, 1.655784e-09, 0.0002255071, 
    -1.44582e-06, 0.06139971, 0.2828247, 0.3025555, 0.01340385, 0.09402367, 
    0.08035074, 0.198414, 0.09535521, 0.1424927, 0.02200292, 0.001765561, 
    0.007960333, 9.181459e-07, 1.659374e-05, 0.05548236, 0.0300127, 
    0.07681681, 0.01088497, 0.006975812, 0.005680757, 0.001818251, 
    2.807953e-08, 0.0008368955,
  0.00183674, 0.004136232, 0.003288372, 0.02735456, 0.007315458, 0.005988449, 
    0.1005322, 0.06829865, 0.04723522, 0.1240216, 0.1509161, 0.07808359, 
    0.09032926, 0.1195572, 0.1405361, 0.07023964, 0.0971239, 0.05482316, 
    0.009171288, 3.287091e-05, 0.02361405, 0.02272809, 0.04690982, 
    0.06384855, 0.1249479, 0.04309769, 0.0791624, 0.03075816, 0.002119775,
  0.09483496, 0.1628763, 0.1798518, 0.0995864, 0.04625594, 0.05484313, 
    0.02930503, 0.07603786, 0.1588068, 0.1650834, 0.1027356, 0.08569244, 
    0.1179387, 0.2006938, 0.07173929, 0.08478816, 0.1683991, 0.1004519, 
    0.1860881, 0.02349794, 0.02751452, 0.03201364, 0.07207131, 0.1028906, 
    0.1371668, 0.156147, 0.1025811, 0.1214185, 0.1190981,
  0.1333746, 0.1426809, 0.08115525, 0.06301635, 0.02884289, 0.1149744, 
    0.1650754, 0.08565607, 0.0827507, 0.1464258, 0.1391642, 0.2119066, 
    0.08857797, 0.1504737, 0.1222653, 0.1561459, 0.1565994, 0.3817404, 
    0.425219, 0.07306305, 0.1199364, 0.1450743, 0.2195509, 0.1882441, 
    0.1587639, 0.3001258, 0.1258523, 0.1801241, 0.1504738,
  0.05833662, 0.1885631, 0.1443089, 0.1349714, 0.1939696, 0.1924355, 
    0.2438123, 0.261927, 0.2243103, 0.227077, 0.2503727, 0.230175, 0.2450492, 
    0.2697158, 0.3099339, 0.1961373, 0.2540197, 0.1435876, 0.2124397, 
    0.2156897, 0.204659, 0.1518958, 0.108642, 0.2390765, 0.04883362, 
    0.2910702, 0.13255, 0.0806701, 0.04899772,
  0.09949026, 0.08563891, 0.1408879, 0.1294186, 0.1640427, 0.257847, 
    0.2073369, 0.1972503, 0.2410679, 0.3609818, 0.4332996, 0.4055107, 
    0.3799514, 0.5207968, 0.4936283, 0.428174, 0.3828822, 0.3177107, 
    0.354352, 0.3038397, 0.2309316, 0.3837533, 0.2458048, 0.1966971, 
    0.1817713, 0.1485374, 0.1571338, 0.05932069, 0.1099356,
  0.01355244, 0.01171181, 0.009871185, 0.008030555, 0.006189925, 0.004349295, 
    0.002508665, 0.0001598558, 0.000647026, 0.001134196, 0.001621366, 
    0.002108537, 0.002595707, 0.003082877, 0.01047933, 0.01269164, 
    0.01490394, 0.01711625, 0.01932855, 0.02154086, 0.02375316, 0.02445713, 
    0.02359828, 0.02273944, 0.02188059, 0.02102175, 0.0201629, 0.01930406, 
    0.01502495,
  0.02348906, -4.27804e-05, -1.005468e-07, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0001123916, 0.0405795, 0.1914037, 0.1263936, 0.139865, 0.125223, 
    0.1942758, 0.1991169, 0.2635525, 0.1858352, 0.1931442, 0.1864914, 
    0.2340904, 0.20567, 0.2123979, 0.2571411, 0.2950574, 0.1717867,
  0.2110143, 0.2945851, 0.2306467, 0.2837086, 0.1244305, 0.1053081, 
    0.1611947, 0.1286332, 0.03451061, 0.1428862, 0.1335112, 0.1476884, 
    0.2568811, 0.3599697, 0.382914, 0.3425016, 0.3103036, 0.3232343, 
    0.3589277, 0.3003049, 0.2832297, 0.2991326, 0.3490941, 0.415338, 
    0.2812381, 0.2347126, 0.2594987, 0.2700872, 0.2285155,
  0.2434804, 0.2149837, 0.2489024, 0.2978282, 0.2809098, 0.249164, 0.26807, 
    0.2895563, 0.2911472, 0.3048075, 0.2932665, 0.2791843, 0.2976764, 
    0.2833138, 0.2457105, 0.2560886, 0.2781797, 0.3081516, 0.3173601, 
    0.3194369, 0.2849986, 0.3166272, 0.2400074, 0.2238864, 0.3143887, 
    0.1784874, 0.1905843, 0.2365227, 0.2894319,
  0.2061282, 0.1678381, 0.1583256, 0.1571877, 0.1630103, 0.1750509, 
    0.1798747, 0.2298701, 0.2254599, 0.2502444, 0.3037881, 0.2802364, 
    0.1965711, 0.1963005, 0.1352724, 0.2017746, 0.1383859, 0.1786683, 
    0.1723895, 0.1702711, 0.1768401, 0.1606801, 0.2132074, 0.1542348, 
    0.128352, 0.1516506, 0.184265, 0.2450367, 0.1703648,
  0.1224836, 0.131107, 0.09247179, 0.117514, 0.08372001, 0.09390853, 
    0.1018238, 0.07941727, 0.0569937, 0.09080424, 0.09905753, 0.1148218, 
    0.07985128, 0.08901305, 0.1510343, 0.1214257, 0.07837845, 0.1055237, 
    0.1104284, 0.100746, 0.1420805, 0.1446175, 0.1403266, 0.1391976, 
    0.07996187, 0.05987071, 0.07677215, 0.1390417, 0.1965768,
  0.01082194, 0.0005714351, 0.1034954, 0.02771651, 0.08542287, 0.1124648, 
    0.01669072, 0.01333263, 0.004225403, 0.01635395, 0.05139248, 0.01338166, 
    0.06494132, 0.05950978, 0.08281584, 0.1269079, 0.1806274, 0.2116584, 
    0.1228548, 0.06232162, 0.1130646, 0.05948861, 0.002797588, 4.603714e-05, 
    0.1760626, 0.08437536, 0.0748426, 0.05155602, 0.03788394,
  7.532876e-08, -6.107793e-05, 0.008727116, 0.009258009, 0.0778574, 
    0.03985759, 0.01302356, 0.00428057, 0.001081123, 0.002668317, 0.03891781, 
    0.03802452, 0.03737861, 0.03748745, 0.1387505, 0.1419402, 0.1159085, 
    0.01566045, 0.006039233, 0.0004519472, 0.0001959272, 5.313151e-08, 
    7.712142e-09, 1.095596e-07, 0.03209461, 0.05638814, 0.01603173, 
    8.402807e-07, 1.072733e-05,
  -6.33746e-07, -0.000384843, 0.003305548, 0.008923102, 0.001268111, 
    0.01433686, 0.07095892, 0.0800663, 0.06507006, 0.003858504, 0.01770691, 
    0.007014161, 0.06545546, 0.09647041, 0.0186407, 0.0461637, 0.003367248, 
    0.0009178007, 0.00118291, 3.667698e-08, 2.751256e-07, 4.946369e-07, 
    5.499243e-06, 0.006504325, 0.08321638, 0.04420412, 0.001568182, 
    4.273381e-08, 1.017165e-07,
  0.007346584, 0.09940286, 0.1019632, 0.003406726, 6.428894e-05, 0.05962969, 
    0.01842272, 0.02977109, 0.0971601, 0.2745737, 0.0397134, 0.1068947, 
    0.2330504, 0.05151648, 0.03024448, 0.008665587, 0.008369087, 0.005842087, 
    0.02014481, 9.682676e-05, 1.723239e-05, 0.004476409, 0.01812499, 
    0.08407981, 0.03714309, 0.0124468, 0.00661153, 0.0007744792, 0.006543088,
  0.1127275, 0.1274205, 0.05150417, 0.3249712, 0.003556205, 0.001787422, 
    0.0275262, 0.02448084, 0.0406967, 0.008980097, 0.005936112, 0.0107111, 
    0.03602939, 0.03854871, 0.07919573, 0.06484982, 0.1306869, 0.2584789, 
    0.2682495, 0.320253, 0.07340942, 0.0776195, 0.1951651, 0.1110416, 
    0.02296303, 0.05579657, 0.09516503, 0.144115, 0.3158249,
  0.0002947271, -6.11659e-06, 2.468035e-06, 1.778265e-06, 5.206493e-06, 
    0.0004793074, 0.1326885, 0.08585516, 0.1930553, 0.07216672, 0.09001283, 
    0.06858077, 0.03268505, 0.0529907, 0.02662943, 0.01280173, 4.185823e-06, 
    2.589356e-07, 3.33458e-05, 0.008802428, 0.0394886, 0.1076896, 0.01196328, 
    0.0121424, 0.005686826, 0.00122547, 6.226645e-05, 7.240712e-06, 
    0.0005846909,
  -1.063467e-07, 0.0002812295, 7.245848e-09, 2.206555e-09, 3.215421e-05, 
    -5.921422e-07, 0.05286885, 0.3140232, 0.3233378, 0.01128868, 0.09000755, 
    0.08466446, 0.1420132, 0.07465731, 0.1014686, 0.01261205, 0.006060412, 
    0.0003266352, 4.254723e-07, 9.086939e-06, 0.06400028, 0.03137369, 
    0.06086854, 0.009722704, 0.005689136, 0.004779934, 0.0005615122, 
    3.281516e-08, 7.068392e-05,
  0.001430854, 0.00128351, 0.004975803, 0.03434565, 0.002491038, 0.009305126, 
    0.08987633, 0.0468188, 0.03846429, 0.1267418, 0.1459126, 0.06682056, 
    0.08468558, 0.1251778, 0.1311644, 0.05623948, 0.0983355, 0.06373042, 
    0.009013508, 0.0001339924, 0.009170693, 0.008319763, 0.05312462, 
    0.05293896, 0.09170187, 0.04024554, 0.0615695, 0.02900655, 0.001578558,
  0.1061357, 0.1901442, 0.170329, 0.1187161, 0.06976032, 0.05543461, 
    0.04793918, 0.08586851, 0.178493, 0.1807935, 0.1115786, 0.08647782, 
    0.08823946, 0.204724, 0.0804392, 0.0779127, 0.1622169, 0.09842248, 
    0.1762336, 0.02120951, 0.01451867, 0.02278738, 0.07528692, 0.1013387, 
    0.150702, 0.1572211, 0.1084955, 0.122721, 0.1240668,
  0.1967101, 0.1432314, 0.1265694, 0.09375021, 0.02689563, 0.1247529, 
    0.2006863, 0.1467948, 0.116163, 0.1694518, 0.1407454, 0.2341712, 
    0.1062892, 0.1836989, 0.140257, 0.1633368, 0.1565618, 0.4257598, 
    0.4181305, 0.08188533, 0.1243347, 0.1615423, 0.233232, 0.197074, 
    0.166019, 0.2912292, 0.1310353, 0.1868173, 0.1458382,
  0.06390698, 0.205185, 0.1595173, 0.132136, 0.2431125, 0.1852069, 0.2490359, 
    0.2845456, 0.2102491, 0.2160903, 0.2641248, 0.2310539, 0.2320782, 
    0.2413973, 0.2793851, 0.2264073, 0.2504308, 0.170797, 0.1893051, 
    0.2150524, 0.1902347, 0.1585253, 0.1318821, 0.2125181, 0.1068078, 
    0.286332, 0.2135209, 0.07328235, 0.0666829,
  0.1182169, 0.08719014, 0.1091958, 0.1782036, 0.2094914, 0.2375672, 
    0.2089781, 0.2095122, 0.2872884, 0.3296124, 0.3128692, 0.4069448, 
    0.4101523, 0.5050184, 0.5082127, 0.4040009, 0.3903646, 0.3276598, 
    0.3439931, 0.2630859, 0.2360148, 0.37756, 0.2791695, 0.2668436, 
    0.1516447, 0.1582625, 0.1522226, 0.05299747, 0.1073738,
  0.02967546, 0.02777132, 0.02586718, 0.02396303, 0.02205889, 0.02015474, 
    0.0182506, 0.02348379, 0.02446851, 0.02545322, 0.02643793, 0.02742264, 
    0.02840735, 0.02939206, 0.0261152, 0.02797682, 0.02983844, 0.03170007, 
    0.03356169, 0.03542331, 0.03728493, 0.03571803, 0.03477585, 0.03383366, 
    0.03289147, 0.03194928, 0.03100709, 0.0300649, 0.03119878,
  0.122583, -0.005069637, -1.96162e-06, 0, 0, 0, 0, 0, 0, 0, -2.013761e-05, 
    0.001079691, 0.0727468, 0.1366198, 0.07756297, 0.09842167, 0.1373173, 
    0.2561666, 0.2505167, 0.2663694, 0.2673229, 0.2793983, 0.1894829, 
    0.2584883, 0.2075321, 0.2088875, 0.2636204, 0.2936607, 0.2604911,
  0.2141372, 0.2930604, 0.2377211, 0.299708, 0.1916684, 0.1686564, 0.1771623, 
    0.1729567, 0.09298785, 0.2620941, 0.227424, 0.2279993, 0.2634324, 
    0.368218, 0.4433187, 0.3404076, 0.2776427, 0.30302, 0.3843096, 0.3412306, 
    0.3212548, 0.3333393, 0.3167639, 0.452206, 0.3255328, 0.2270514, 
    0.2352333, 0.3017837, 0.2353613,
  0.2406098, 0.2121321, 0.2514492, 0.3003139, 0.3084102, 0.2592029, 
    0.2755757, 0.2814443, 0.3284027, 0.3272841, 0.3014349, 0.2933254, 
    0.3127144, 0.3316799, 0.2955381, 0.2767063, 0.2741977, 0.3259606, 
    0.3518786, 0.3518486, 0.3189372, 0.326755, 0.2489349, 0.2142518, 
    0.3141118, 0.1976883, 0.2157388, 0.2503116, 0.2944225,
  0.2246473, 0.1895878, 0.1779921, 0.1807536, 0.1872988, 0.1909557, 
    0.2172427, 0.2697738, 0.2416369, 0.268052, 0.3010901, 0.3309698, 
    0.2148636, 0.1850816, 0.1155349, 0.2150188, 0.1402134, 0.1963107, 
    0.17915, 0.1849129, 0.2164006, 0.2173261, 0.2453172, 0.1540728, 
    0.1132208, 0.1487063, 0.2095496, 0.2736024, 0.2148726,
  0.1319139, 0.1479142, 0.09991205, 0.1243138, 0.1111239, 0.1087191, 
    0.1178005, 0.08498924, 0.08151025, 0.1162388, 0.1095173, 0.1376471, 
    0.08127997, 0.09340169, 0.155771, 0.1542264, 0.1133885, 0.1178162, 
    0.1138957, 0.1113893, 0.1563509, 0.1573707, 0.1406484, 0.1428584, 
    0.07752424, 0.06034019, 0.1145355, 0.1644811, 0.2076075,
  0.0134271, 0.001829745, 0.09069698, 0.02353546, 0.08770407, 0.1150043, 
    0.02655948, 0.02762239, 0.0105184, 0.01709585, 0.03656037, 0.01579184, 
    0.1059205, 0.0656926, 0.09819376, 0.1310572, 0.1858359, 0.2098839, 
    0.1246066, 0.08123837, 0.12851, 0.07780939, 0.009713712, 5.230865e-05, 
    0.1669131, 0.07737383, 0.07975169, 0.05133675, 0.04129704,
  1.627241e-07, -3.432157e-06, 0.03220335, 0.01498337, 0.07096469, 
    0.03634625, 0.02695397, 0.04816091, 0.0216114, 0.001536617, 0.01053187, 
    0.03612064, 0.07323552, 0.02819016, 0.156331, 0.1217876, 0.1282125, 
    0.05959034, 0.01207989, 0.006687113, 0.004823009, -2.478726e-06, 
    5.2398e-08, 9.485959e-08, 0.04408332, 0.0676481, 0.0283788, 0.0005610058, 
    0.002331716,
  -4.730756e-08, -2.922691e-05, 0.01214316, 0.03914328, 0.005985311, 
    0.02072296, 0.05297814, 0.08559957, 0.05494613, 0.002720732, 0.02369397, 
    0.006820019, 0.08270016, 0.09132566, 0.02119202, 0.05092688, 0.009936011, 
    0.002019964, 0.001381339, -3.166888e-07, 2.799459e-07, 3.741064e-07, 
    1.418513e-06, 0.00684878, 0.02727243, 0.01814765, 0.01545535, 
    3.022337e-06, 1.278746e-07,
  0.0003218762, 0.1050964, 0.06300356, 0.001728288, 0.0002635085, 0.05984004, 
    0.01617294, 0.02808927, 0.08972269, 0.2494007, 0.04549111, 0.07103651, 
    0.196257, 0.04639173, 0.03353011, 0.01554577, 0.00506017, 0.002340221, 
    0.008205481, 0.000188714, 0.000389106, 0.00692769, 0.01241293, 
    0.07828794, 0.02776874, 0.008307473, 0.007144135, 8.208364e-05, 
    0.0004713311,
  0.09084214, 0.08805598, 0.03348516, 0.3500549, 0.0007973908, 0.001462949, 
    0.02489353, 0.02721828, 0.02849841, 0.009592212, 0.006536821, 0.01103123, 
    0.03733496, 0.03206139, 0.07468377, 0.06402776, 0.142566, 0.2264274, 
    0.248793, 0.307563, 0.05444501, 0.06856108, 0.1868607, 0.1042028, 
    0.02350927, 0.05406083, 0.1003966, 0.1402247, 0.275268,
  9.397417e-05, 3.538549e-09, 6.649473e-07, 7.404848e-07, 1.334875e-06, 
    1.72661e-05, 0.09651081, 0.1024373, 0.2033045, 0.0800607, 0.07707869, 
    0.06381037, 0.03219073, 0.04865577, 0.02404952, 0.01430203, 3.835987e-05, 
    4.935326e-07, 3.368454e-05, 0.008064251, 0.03746126, 0.1166437, 
    0.01150505, 0.01163658, 0.006624992, 0.002197772, 4.059509e-06, 
    2.16241e-06, 0.0002968674,
  -3.327555e-08, 4.919454e-05, 1.888067e-08, 1.429826e-09, 7.345196e-06, 
    -4.162372e-08, 0.04982478, 0.333808, 0.3715321, 0.01483283, 0.09220841, 
    0.09532727, 0.1090365, 0.0655895, 0.06412981, 0.0151737, 0.01033953, 
    0.0002340791, 2.500381e-07, 3.500415e-06, 0.0413577, 0.03709393, 
    0.05542913, 0.009553367, 0.00455344, 0.007674293, 0.001040606, 
    2.705637e-08, 1.677592e-05,
  0.0009127474, 0.0007855695, 0.009086125, 0.02418459, 0.0001352657, 
    0.007782831, 0.064026, 0.02599197, 0.02498941, 0.1354565, 0.1332049, 
    0.06625219, 0.09719314, 0.1133133, 0.1259591, 0.04612624, 0.1021914, 
    0.07508412, 0.009762176, 5.808065e-05, 0.005073048, 0.007894418, 
    0.0541316, 0.04667052, 0.07485393, 0.03891721, 0.06271749, 0.03010455, 
    0.001670783,
  0.1333266, 0.2148437, 0.1617786, 0.1452472, 0.05835773, 0.06053475, 
    0.05759034, 0.1141073, 0.2114104, 0.1946428, 0.1099101, 0.07943885, 
    0.07408659, 0.1815478, 0.06191534, 0.06227881, 0.1739577, 0.1075167, 
    0.1986188, 0.02286671, 0.00828461, 0.01140819, 0.06703813, 0.1254437, 
    0.1703093, 0.1711394, 0.1121125, 0.1200197, 0.1250222,
  0.2047297, 0.1843756, 0.1351449, 0.1123136, 0.06079983, 0.138788, 
    0.2164337, 0.1477633, 0.1496114, 0.2076258, 0.1495588, 0.2500593, 
    0.1348952, 0.1911195, 0.1657094, 0.1730158, 0.2237001, 0.4795788, 
    0.4569709, 0.1312258, 0.1384955, 0.1800867, 0.2247554, 0.1889831, 
    0.1519058, 0.3002764, 0.1700169, 0.2068225, 0.1648814,
  0.1214437, 0.1761562, 0.1619456, 0.1491429, 0.2615604, 0.1884804, 
    0.2586106, 0.3305647, 0.2069157, 0.2160516, 0.2605249, 0.2373797, 
    0.2418959, 0.2651762, 0.3005305, 0.2548356, 0.2507076, 0.2000172, 
    0.2112645, 0.2253487, 0.2291588, 0.2016188, 0.147143, 0.1794974, 
    0.1161098, 0.2897629, 0.1479412, 0.07136548, 0.07956061,
  0.1622527, 0.1792465, 0.1953784, 0.2099295, 0.2490075, 0.2951775, 
    0.2949684, 0.272567, 0.2838658, 0.3387093, 0.410391, 0.5113818, 
    0.5313352, 0.5633385, 0.5644696, 0.4703459, 0.4138452, 0.3114395, 
    0.3227285, 0.2794025, 0.2382168, 0.4030639, 0.2761595, 0.2349788, 
    0.1603965, 0.1719984, 0.1606846, 0.08319212, 0.1715015,
  0.05576523, 0.051435, 0.04710477, 0.04277454, 0.03844431, 0.03411408, 
    0.02978385, 0.03542552, 0.03728193, 0.03913834, 0.04099475, 0.04285116, 
    0.04470757, 0.04656398, 0.04175255, 0.04496554, 0.04817853, 0.05139152, 
    0.0546045, 0.05781749, 0.06103048, 0.07497329, 0.07423413, 0.07349496, 
    0.07275579, 0.07201663, 0.07127746, 0.0705383, 0.05922941,
  0.1631925, 0.01606301, -7.133435e-05, 0, 0, -0.0004520692, 0.0001231653, 0, 
    0, 0, 0.0005825327, 0.02249188, 0.08804929, 0.1114691, 0.05751512, 
    0.07515104, 0.122616, 0.2404257, 0.2692552, 0.2837373, 0.3083985, 
    0.3544021, 0.1847469, 0.243065, 0.2129292, 0.2113634, 0.2535324, 
    0.2949123, 0.2898274,
  0.2356709, 0.2744496, 0.2349201, 0.2944775, 0.2592428, 0.2066784, 
    0.1814548, 0.2508464, 0.1864792, 0.3568704, 0.2886183, 0.2513781, 
    0.246193, 0.381291, 0.3892101, 0.2944962, 0.2371062, 0.2744953, 
    0.2683393, 0.3001439, 0.3333761, 0.3303948, 0.2574695, 0.481858, 
    0.3049393, 0.2156217, 0.2283427, 0.2606821, 0.2414996,
  0.2434934, 0.2529395, 0.2662612, 0.3014288, 0.3442549, 0.3036676, 
    0.2886968, 0.2945692, 0.3514616, 0.3328497, 0.3226083, 0.2844242, 
    0.3164999, 0.3243922, 0.2801481, 0.2534202, 0.3041216, 0.348187, 
    0.3731453, 0.3483886, 0.3392227, 0.3153887, 0.2481561, 0.2408613, 
    0.3026075, 0.1948044, 0.2372546, 0.2612312, 0.2859504,
  0.2538092, 0.2143637, 0.1922782, 0.2097996, 0.1912415, 0.1931125, 
    0.2228968, 0.2852876, 0.2436064, 0.2846676, 0.3053057, 0.3100384, 
    0.2311975, 0.2067419, 0.1196515, 0.234947, 0.1565032, 0.1987607, 
    0.1565326, 0.1949181, 0.200598, 0.2041589, 0.2550209, 0.1582103, 
    0.1056585, 0.1590122, 0.2138156, 0.2862396, 0.2127967,
  0.1430303, 0.1792236, 0.1149534, 0.1495914, 0.1246269, 0.1413352, 
    0.1274335, 0.1084086, 0.1216406, 0.1494229, 0.1183908, 0.1498348, 
    0.1003839, 0.09777173, 0.1720859, 0.1911268, 0.1229499, 0.1502252, 
    0.121117, 0.123854, 0.1884673, 0.163784, 0.1596446, 0.1534926, 
    0.08198556, 0.07232256, 0.139935, 0.1717879, 0.2324576,
  0.0229066, 0.00781458, 0.07006341, 0.02491222, 0.08982112, 0.121558, 
    0.03151833, 0.03633132, 0.02088557, 0.02581656, 0.01508397, 0.01261044, 
    0.1433844, 0.07383527, 0.1112334, 0.1492488, 0.189558, 0.1873305, 
    0.1291987, 0.1030534, 0.1346613, 0.1133078, 0.009702871, 2.449199e-05, 
    0.1182477, 0.06269392, 0.07051922, 0.06451587, 0.04836458,
  2.015682e-07, -1.756955e-07, 0.02451951, 0.02446559, 0.0668892, 0.03551492, 
    0.04964824, 0.04516318, 0.03526857, 0.0004284738, 0.00076974, 0.08198639, 
    0.09042278, 0.03389865, 0.1278539, 0.1056689, 0.1345554, 0.06436483, 
    0.01738591, 0.02861225, 0.01457482, 0.0001650348, 3.34668e-07, 
    8.421165e-08, 0.01259416, 0.07383432, 0.06199149, 0.008291531, 0.007187949,
  2.330145e-08, -2.50768e-06, 0.002908018, 0.1147126, 0.01213495, 0.02753566, 
    0.05020811, 0.1015925, 0.04693643, 0.004004442, 0.03327519, 0.008835425, 
    0.1102209, 0.0875989, 0.02459323, 0.05890819, 0.01611208, 0.007042665, 
    0.005947908, 1.416467e-06, 3.489678e-07, 1.660114e-07, 7.407212e-07, 
    0.006904302, 0.004118179, 0.006390123, 0.02934981, 0.0004224102, 
    3.901602e-07,
  0.0001459897, 0.1144829, 0.03829153, 0.006911012, 0.002281752, 0.05908855, 
    0.01503787, 0.0265771, 0.0900815, 0.2482389, 0.0498182, 0.05133619, 
    0.1759692, 0.04123331, 0.03284086, 0.02343585, 0.01205009, 0.001968838, 
    0.001573685, 0.001717805, 0.004075201, 0.007491476, 0.01107758, 
    0.07513439, 0.02233965, 0.006270466, 0.01026167, 2.618662e-05, 0.001522318,
  0.06786784, 0.06526776, 0.0290904, 0.2611176, 0.0008749234, 0.001673832, 
    0.02748707, 0.02844405, 0.02491597, 0.01024725, 0.008294746, 0.01353052, 
    0.04165555, 0.02709242, 0.06500105, 0.06253636, 0.1423604, 0.2047398, 
    0.2417862, 0.2865825, 0.04420356, 0.06823314, 0.1931914, 0.1013617, 
    0.02399653, 0.05357953, 0.09744657, 0.1376686, 0.2342309,
  4.094822e-05, 3.767248e-07, 1.393068e-07, -7.874556e-08, 4.564474e-07, 
    4.254176e-06, 0.09870897, 0.1029565, 0.2106296, 0.07750171, 0.06327181, 
    0.06097452, 0.03201439, 0.04663772, 0.02338787, 0.02243985, 0.001097793, 
    8.863551e-05, 0.0002634597, 0.008979258, 0.03597732, 0.1256462, 
    0.01334689, 0.01192785, 0.01343913, 0.009131646, 9.973917e-05, 
    4.310668e-07, 8.950382e-05,
  -3.093424e-09, 2.129716e-05, -2.302116e-08, 1.858342e-10, 2.369248e-06, 
    -1.564965e-08, 0.03768658, 0.413149, 0.3652776, 0.02066706, 0.09558436, 
    0.1058071, 0.0950375, 0.06087358, 0.04305432, 0.01580941, 0.02946071, 
    0.001164196, 1.488337e-07, 1.44533e-06, 0.01666741, 0.04412863, 
    0.05103114, 0.01123825, 0.004772622, 0.008370202, 0.00822672, 
    1.565686e-05, 7.687017e-06,
  0.0006553612, 0.001333436, 0.009321552, 0.02894089, -7.791309e-05, 
    0.002864462, 0.04381867, 0.01708041, 0.01417455, 0.07960071, 0.1359847, 
    0.07147882, 0.09612408, 0.1176968, 0.1239398, 0.05165659, 0.09307504, 
    0.07953345, 0.02200996, 2.362991e-05, 0.002375186, 0.003889524, 
    0.05327983, 0.04548674, 0.06742894, 0.04106521, 0.06616416, 0.03255159, 
    0.002453834,
  0.1170677, 0.2209192, 0.1736714, 0.1437213, 0.02101429, 0.05403779, 
    0.06544983, 0.1441493, 0.2344441, 0.1861078, 0.1119647, 0.08744403, 
    0.06378906, 0.1699068, 0.06521513, 0.04974203, 0.1766592, 0.1263253, 
    0.1744965, 0.03419438, 0.007891783, 0.005280337, 0.06340671, 0.1700916, 
    0.1678235, 0.1878203, 0.1345526, 0.112922, 0.1206154,
  0.2575987, 0.1976705, 0.1365547, 0.1090227, 0.09706423, 0.1476563, 
    0.2052841, 0.1488741, 0.2036645, 0.2159432, 0.1759684, 0.2662331, 
    0.1200591, 0.2177819, 0.1746141, 0.1842265, 0.2889329, 0.4931833, 
    0.4509642, 0.1066127, 0.132167, 0.1427652, 0.2190645, 0.2093107, 
    0.1362315, 0.3307635, 0.2083625, 0.2833217, 0.198451,
  0.1259088, 0.2517197, 0.2016958, 0.1733458, 0.3195566, 0.2650176, 
    0.2645114, 0.3317988, 0.2509557, 0.2314634, 0.3044683, 0.2927328, 
    0.2708986, 0.2617123, 0.3170965, 0.2400682, 0.2801789, 0.2448371, 
    0.2135484, 0.2425319, 0.2166569, 0.2502958, 0.1603687, 0.1766039, 
    0.08096711, 0.2898813, 0.1283753, 0.07730496, 0.1042245,
  0.2292139, 0.2849824, 0.2334974, 0.2379365, 0.2666642, 0.3237133, 
    0.2608443, 0.3094022, 0.3489231, 0.3617654, 0.3808584, 0.4620696, 
    0.4605144, 0.545851, 0.5811075, 0.4648212, 0.4162416, 0.3149541, 
    0.3481198, 0.3107409, 0.2425502, 0.4553847, 0.3255346, 0.2037404, 
    0.1392581, 0.154681, 0.141622, 0.08766792, 0.1748795,
  0.1170336, 0.1128706, 0.1087075, 0.1045445, 0.1003815, 0.09621852, 
    0.09205551, 0.1154888, 0.1181907, 0.1208926, 0.1235944, 0.1262963, 
    0.1289982, 0.1317001, 0.1152283, 0.1189116, 0.1225948, 0.126278, 
    0.1299612, 0.1336444, 0.1373276, 0.1266653, 0.1244432, 0.1222211, 
    0.1199991, 0.117777, 0.1155549, 0.1133328, 0.120364,
  0.2129585, 0.05194824, 0.007872252, -0.0001444329, 0, -0.001948192, 
    -0.0008910495, 0, 0, 5.511761e-05, 0.02087785, 0.0488483, 0.121643, 
    0.1009165, 0.05706367, 0.1007129, 0.1373389, 0.2095933, 0.2642531, 
    0.2705658, 0.3365416, 0.3944078, 0.2118172, 0.2408417, 0.2042862, 
    0.2428589, 0.2393144, 0.2898466, 0.2851023,
  0.2709178, 0.2452294, 0.2490335, 0.3055143, 0.2927099, 0.2199252, 
    0.1863167, 0.3180059, 0.2431424, 0.3955542, 0.3069772, 0.2556472, 
    0.2275292, 0.3781529, 0.3675247, 0.254269, 0.1986342, 0.2411071, 
    0.2431409, 0.3028496, 0.3929959, 0.2954886, 0.2987944, 0.4697596, 
    0.3089778, 0.1655474, 0.2202577, 0.2696427, 0.2495049,
  0.2843794, 0.2408646, 0.2651601, 0.3446832, 0.390646, 0.3094402, 0.3129891, 
    0.3085684, 0.3431764, 0.3350372, 0.3398396, 0.2875393, 0.2684049, 
    0.2917222, 0.235434, 0.2384652, 0.2851693, 0.2807908, 0.348672, 
    0.3530409, 0.3505113, 0.2998783, 0.2589365, 0.2435084, 0.2839364, 
    0.1723902, 0.1921581, 0.2601765, 0.308343,
  0.2846932, 0.2380799, 0.2123069, 0.2162827, 0.2094457, 0.2155903, 
    0.2397979, 0.3120877, 0.270977, 0.2895288, 0.3132254, 0.2999795, 
    0.2443034, 0.262151, 0.152173, 0.2615669, 0.1785222, 0.2350567, 
    0.2009539, 0.2006819, 0.2289567, 0.2017801, 0.243728, 0.1636436, 
    0.09841489, 0.1879757, 0.2299007, 0.2747476, 0.2320672,
  0.1805546, 0.2098275, 0.1362676, 0.1756558, 0.1257482, 0.1463933, 
    0.1265646, 0.1400772, 0.1593308, 0.1985934, 0.1538375, 0.160531, 
    0.1217917, 0.1065149, 0.1890521, 0.2018666, 0.1451637, 0.144379, 
    0.1316276, 0.1393586, 0.2067806, 0.1731542, 0.1684997, 0.1716503, 
    0.07845976, 0.1050998, 0.1494353, 0.1819486, 0.2642477,
  0.05910584, 0.02712383, 0.05520044, 0.03713553, 0.09679367, 0.1148366, 
    0.05359442, 0.03312086, 0.03855102, 0.04299061, 0.0100081, 0.01047918, 
    0.1280388, 0.08706658, 0.1080767, 0.1659229, 0.1981125, 0.1728899, 
    0.1451325, 0.1083441, 0.146671, 0.1285415, 0.01341194, 1.139422e-05, 
    0.08286151, 0.05179856, 0.05268314, 0.07280339, 0.08246344,
  -1.486719e-05, 3.217511e-08, 0.002493095, 0.03883042, 0.07525562, 
    0.02635961, 0.04026507, 0.05090513, 0.05163512, 0.0001104503, 
    3.721446e-05, 0.0162513, 0.09706505, 0.04372215, 0.1225975, 0.08827923, 
    0.1287636, 0.07009445, 0.02720961, 0.04490248, 0.0484732, 0.001885469, 
    7.51236e-06, 8.589487e-08, 0.0005302952, 0.1297519, 0.07390185, 
    0.03655355, 0.01820784,
  3.882719e-08, -2.962678e-07, -8.274927e-06, 0.104253, 0.01849645, 
    0.02330294, 0.04711832, 0.1052769, 0.06575982, 0.01335402, 0.04356093, 
    0.02618928, 0.1277431, 0.08396427, 0.02570658, 0.05449909, 0.01370954, 
    0.008700841, 0.01111145, 0.0001205781, 1.521898e-06, 4.054022e-07, 
    5.858587e-07, 0.009902867, 0.002045445, 0.001074346, 0.04042974, 
    0.002963763, 6.16634e-06,
  0.0004520049, 0.1459642, 0.02285241, 0.02017201, 0.01305052, 0.05448942, 
    0.01338323, 0.02558265, 0.08648368, 0.2598307, 0.05008968, 0.03975255, 
    0.1367057, 0.03386301, 0.02935442, 0.02653171, 0.02586296, 0.005942434, 
    0.002648988, 0.004463342, 0.005182327, 0.01200818, 0.01342096, 
    0.07902799, 0.02121353, 0.006399905, 0.014438, 0.001469074, 0.000164607,
  0.0527496, 0.05660306, 0.03149837, 0.1840534, 2.787344e-05, 0.002289508, 
    0.02961965, 0.0254259, 0.02272038, 0.01142547, 0.01658759, 0.01657145, 
    0.04028659, 0.02561159, 0.05168819, 0.05897193, 0.124999, 0.2005174, 
    0.2377581, 0.2807897, 0.05731671, 0.06761842, 0.208867, 0.09888976, 
    0.02169042, 0.04621686, 0.08952597, 0.1350229, 0.1898528,
  9.483235e-06, 1.423251e-07, 4.055562e-08, -5.213919e-07, 1.414016e-07, 
    1.495231e-06, 0.1131864, 0.1002109, 0.2219591, 0.07090553, 0.05069871, 
    0.05641837, 0.03094567, 0.04176657, 0.02402597, 0.02392493, 0.01180232, 
    0.001006501, 0.0001152763, 0.01067554, 0.03381876, 0.1221299, 0.012666, 
    0.01164043, 0.023071, 0.01842603, 0.005203291, 7.185739e-08, 2.666465e-05,
  -4.227823e-09, 1.260455e-05, -1.593485e-07, 9.818275e-12, 1.086057e-06, 
    -9.817078e-09, 0.02146959, 0.3941826, 0.363603, 0.03787839, 0.09653991, 
    0.1077004, 0.09210936, 0.05901097, 0.03574133, 0.02308434, 0.04612613, 
    0.003594591, -1.17773e-07, 6.09015e-07, 0.008270445, 0.05327972, 
    0.04668521, 0.0116232, 0.007006137, 0.01245176, 0.03361139, 0.002670741, 
    3.759638e-06,
  0.002855788, 0.003773205, 0.009895099, 0.03869173, -2.221647e-05, 
    0.003393854, 0.02580049, 0.008709302, 0.006916753, 0.062304, 0.1461281, 
    0.08602463, 0.1135907, 0.1135964, 0.1316555, 0.07204986, 0.09322675, 
    0.09655579, 0.01868363, 1.746518e-05, 0.001087057, 0.002562291, 
    0.04252104, 0.0400776, 0.07870957, 0.04882309, 0.07852865, 0.05206471, 
    0.007941033,
  0.1168432, 0.2158249, 0.1871205, 0.09145676, 0.006970086, 0.06706608, 
    0.04130579, 0.1133988, 0.2293911, 0.1616518, 0.1220219, 0.09770373, 
    0.05284452, 0.1762825, 0.06862946, 0.0504869, 0.1626763, 0.1731814, 
    0.2022045, 0.03837357, 0.005437417, 0.006952811, 0.06767475, 0.1740466, 
    0.171398, 0.1658492, 0.1294835, 0.1345353, 0.1325861,
  0.2430753, 0.2007276, 0.1467497, 0.1112648, 0.09737647, 0.1529365, 
    0.210032, 0.1670494, 0.1961711, 0.2055007, 0.1470503, 0.2612342, 
    0.09951203, 0.2325218, 0.1797306, 0.2167931, 0.3622993, 0.4893211, 
    0.462917, 0.1079229, 0.1084701, 0.1407681, 0.20324, 0.2356558, 0.1357031, 
    0.3256274, 0.2381325, 0.2574839, 0.2136986,
  0.1789817, 0.2312616, 0.2689605, 0.1677473, 0.2847129, 0.2298902, 
    0.2342607, 0.3517101, 0.2797345, 0.2700745, 0.3531011, 0.2622384, 
    0.2483169, 0.2435033, 0.2900545, 0.1953504, 0.2577909, 0.2121744, 
    0.2429682, 0.2464348, 0.2381957, 0.2573197, 0.1847325, 0.1823184, 
    0.08142107, 0.3167822, 0.1324978, 0.07105293, 0.1138094,
  0.1781633, 0.2684598, 0.2755611, 0.2082019, 0.2225589, 0.330579, 0.2986231, 
    0.2737, 0.2592086, 0.2926746, 0.3197879, 0.4210386, 0.3973686, 0.4776438, 
    0.5191882, 0.4538382, 0.4258171, 0.3092201, 0.3394333, 0.3260985, 
    0.2551705, 0.492007, 0.352112, 0.2397326, 0.127933, 0.1476714, 0.1321894, 
    0.1111613, 0.1609576,
  0.1466008, 0.1404632, 0.1343256, 0.1281881, 0.1220505, 0.1159129, 
    0.1097754, 0.1360871, 0.139215, 0.142343, 0.145471, 0.1485989, 0.1517269, 
    0.1548549, 0.1514076, 0.1568441, 0.1622806, 0.1677171, 0.1731537, 
    0.1785902, 0.1840267, 0.1654709, 0.163044, 0.1606171, 0.1581902, 
    0.1557633, 0.1533364, 0.1509095, 0.1515108,
  0.2292565, 0.1133222, 0.01344637, 0.002720024, -0.0004937006, -0.002477397, 
    0.005675649, -0.0005507059, 0.0002225076, -0.0001845549, 0.05066545, 
    0.0508181, 0.1156403, 0.09448563, 0.07048365, 0.1089253, 0.1068954, 
    0.1843485, 0.2551883, 0.2493173, 0.3880188, 0.4209013, 0.2567407, 
    0.2241816, 0.2076723, 0.2508806, 0.2416681, 0.2708912, 0.2904742,
  0.2880358, 0.2311431, 0.2587294, 0.303864, 0.3089938, 0.2337098, 0.1853247, 
    0.3504332, 0.291153, 0.3879098, 0.2993031, 0.2475727, 0.2156461, 
    0.3627015, 0.375572, 0.2405493, 0.2067044, 0.218724, 0.2923835, 
    0.3157037, 0.3983714, 0.3193969, 0.3164916, 0.4637212, 0.2892188, 
    0.2071736, 0.2226882, 0.3294084, 0.2820491,
  0.2884189, 0.2234979, 0.3229594, 0.436334, 0.4227915, 0.3262362, 0.2998239, 
    0.3123532, 0.3980292, 0.344146, 0.324707, 0.3186541, 0.263852, 0.3188291, 
    0.2543144, 0.2694651, 0.2969691, 0.3011393, 0.4072299, 0.3961651, 
    0.3746172, 0.3512428, 0.2524674, 0.245316, 0.276455, 0.170663, 0.232622, 
    0.2303293, 0.3372453,
  0.3186027, 0.2758538, 0.2520935, 0.2416614, 0.2609694, 0.251932, 0.2820219, 
    0.3473004, 0.250643, 0.2845089, 0.324445, 0.3031722, 0.2690668, 
    0.2593399, 0.1711421, 0.2747479, 0.2235042, 0.3109013, 0.2452066, 
    0.2205781, 0.2388185, 0.1863722, 0.2408094, 0.176995, 0.1050698, 
    0.2203057, 0.2415219, 0.3192893, 0.2570701,
  0.2164146, 0.2381034, 0.1771602, 0.2260361, 0.1807436, 0.2502024, 
    0.1750132, 0.1676585, 0.2201207, 0.2295076, 0.1794545, 0.1898335, 
    0.1336136, 0.1276626, 0.2077982, 0.2167819, 0.1708279, 0.1582619, 
    0.1599553, 0.1658424, 0.2266796, 0.192925, 0.1928588, 0.1970333, 
    0.06913357, 0.1776885, 0.2200199, 0.2456031, 0.2865375,
  0.1663655, 0.04063114, 0.04125974, 0.0615115, 0.1015403, 0.1090632, 
    0.09123898, 0.06172118, 0.07987906, 0.07258166, 0.01060551, 0.000571867, 
    0.08198556, 0.1182593, 0.1190891, 0.1733381, 0.1974983, 0.1894031, 
    0.1612451, 0.1161632, 0.1864414, 0.1732204, 0.03686891, 0.0005038265, 
    0.08313618, 0.06667814, 0.07831848, 0.1123144, 0.09945166,
  0.06544739, -3.36555e-07, 0.0001030094, 0.03641533, 0.08738535, 0.02984349, 
    0.04305824, 0.07933455, 0.1427567, 0.01980312, -1.243327e-05, 
    0.001952445, 0.09830494, 0.08742084, 0.1182517, 0.07157255, 0.1219033, 
    0.07437322, 0.02802911, 0.05279026, 0.0856601, 0.1154854, 0.006400954, 
    4.717759e-08, 0.0006058309, 0.02028158, 0.05351755, 0.09738272, 0.06733226,
  7.218752e-07, 2.218676e-06, -2.001628e-05, 0.05914885, 0.01519452, 
    0.03055911, 0.05127324, 0.0950302, 0.08136017, 0.0229148, 0.04422544, 
    0.03797873, 0.1624929, 0.08048096, 0.02487909, 0.04825579, 0.01700245, 
    0.01021133, 0.0169924, 0.01569464, 0.0008436851, 6.563185e-06, 
    4.071543e-07, 0.01234934, 0.00155371, 0.0001822791, 0.03597571, 
    0.03638712, 0.0001661586,
  0.0006067194, 0.1776024, 0.01732338, 0.02429125, 0.02731961, 0.05046235, 
    0.01222972, 0.02358207, 0.07670403, 0.2424693, 0.04829684, 0.02695819, 
    0.1057383, 0.02903824, 0.0256801, 0.02300209, 0.03630599, 0.0152679, 
    0.01610184, 0.01596729, 0.003061804, 0.01023771, 0.01718517, 0.07892808, 
    0.02396271, 0.007634995, 0.01647858, 0.01530928, 0.0004371174,
  0.0634798, 0.05012301, 0.02869866, 0.1456734, -0.0001245334, 0.006223965, 
    0.03119154, 0.02451837, 0.01804919, 0.01298911, 0.08048712, 0.02068112, 
    0.03426002, 0.02182663, 0.04041872, 0.05083639, 0.1049516, 0.191609, 
    0.2052822, 0.2610657, 0.06672136, 0.06211503, 0.2151311, 0.09772665, 
    0.01988059, 0.0399222, 0.08163484, 0.1248363, 0.1613956,
  2.887382e-07, 5.289617e-08, 2.011543e-08, -6.025433e-07, 8.809745e-08, 
    -7.884306e-05, 0.1358334, 0.08147421, 0.2205036, 0.06206966, 0.03829433, 
    0.04655395, 0.02794345, 0.03774058, 0.02785725, 0.03615845, 0.02655797, 
    0.005991986, 3.998318e-05, 0.0129611, 0.03264317, 0.1166032, 0.01289905, 
    0.01329308, 0.02870971, 0.02420493, 0.01313145, 2.303159e-07, 6.114592e-06,
  -3.896837e-09, 6.561976e-06, 5.792101e-06, 2.583185e-12, 6.06792e-07, 
    -7.355487e-09, 0.0147103, 0.3458354, 0.351641, 0.05147048, 0.09318392, 
    0.09845743, 0.09001437, 0.05269976, 0.03714945, 0.02951275, 0.06074892, 
    0.02583653, 0.0007757021, 2.87151e-07, 0.003106236, 0.05589961, 
    0.04309997, 0.01450714, 0.009226136, 0.01833908, 0.0406166, 0.01023461, 
    2.353135e-06,
  0.006120597, 0.009763212, 0.00479961, 0.0533394, -3.62424e-05, 
    0.0009741858, 0.01658533, 0.003315392, 0.003769763, 0.0603218, 0.1760233, 
    0.1092708, 0.1417398, 0.1220573, 0.1640941, 0.1066116, 0.1509496, 
    0.1425697, 0.03502851, -6.832843e-05, 0.0005423889, 0.001264862, 
    0.02939961, 0.03531763, 0.08952943, 0.05332576, 0.1033935, 0.1030542, 
    0.01004972,
  0.1377123, 0.2371785, 0.1830219, 0.06177298, 0.01091171, 0.04605597, 
    0.04164841, 0.1164725, 0.2301731, 0.1496353, 0.1336849, 0.1051119, 
    0.05100131, 0.1874506, 0.0765609, 0.04218063, 0.1861508, 0.2199857, 
    0.2652757, 0.05218922, 0.003370752, 0.00798439, 0.08736333, 0.1782288, 
    0.1702741, 0.1690058, 0.1725321, 0.1828001, 0.1397676,
  0.2337405, 0.2212103, 0.1608916, 0.1499666, 0.1277443, 0.1485225, 
    0.1938086, 0.1962147, 0.1930026, 0.2421252, 0.1701218, 0.284131, 
    0.102171, 0.2626984, 0.1824706, 0.3000889, 0.4066747, 0.518755, 
    0.4438373, 0.08408436, 0.08384244, 0.1411292, 0.1767177, 0.2251109, 
    0.1414722, 0.3080682, 0.2445583, 0.2812478, 0.2231806,
  0.2369823, 0.2688667, 0.2836136, 0.1728792, 0.2857179, 0.2237802, 
    0.2387802, 0.4076325, 0.3220907, 0.2692749, 0.3403895, 0.2719954, 
    0.2851337, 0.3058704, 0.351329, 0.1829266, 0.2914021, 0.1928569, 
    0.2202704, 0.2123037, 0.2132761, 0.2381396, 0.1719164, 0.1747881, 
    0.09029482, 0.3159407, 0.1461213, 0.07620668, 0.1446326,
  0.1962149, 0.2110795, 0.2531707, 0.2595035, 0.2744653, 0.3716711, 
    0.3105909, 0.269782, 0.2374054, 0.2838637, 0.3092856, 0.4817515, 
    0.4401572, 0.5402843, 0.5711415, 0.4346447, 0.4102283, 0.3052295, 
    0.3327746, 0.3363708, 0.278165, 0.5106578, 0.4011302, 0.2994513, 
    0.1352606, 0.184929, 0.1573327, 0.1131261, 0.1820894,
  0.2039614, 0.1972816, 0.1906018, 0.1839219, 0.1772421, 0.1705622, 
    0.1638824, 0.1761573, 0.1780302, 0.1799031, 0.1817759, 0.1836488, 
    0.1855217, 0.1873946, 0.1765869, 0.1832751, 0.1899633, 0.1966515, 
    0.2033396, 0.2100278, 0.216716, 0.2174007, 0.2155194, 0.2136382, 
    0.211757, 0.2098758, 0.2079946, 0.2061134, 0.2093053,
  0.2318809, 0.1477728, 0.02311045, 0.01724694, 4.272915e-05, 0.005612806, 
    0.02632305, 0.001194485, 0.0003043015, 0.03387197, 0.06331589, 
    0.06413606, 0.1409233, 0.09150515, 0.08104878, 0.1186943, 0.0999831, 
    0.1680094, 0.2601346, 0.2185666, 0.3825891, 0.4257429, 0.3040628, 
    0.2313771, 0.2356643, 0.2276514, 0.2469568, 0.244777, 0.2922482,
  0.304369, 0.2082943, 0.2852816, 0.2852374, 0.3128636, 0.2277738, 0.1765913, 
    0.3650738, 0.3093239, 0.3792585, 0.2924865, 0.2095508, 0.2244163, 
    0.351989, 0.3776976, 0.2554299, 0.2615214, 0.2163722, 0.3994622, 
    0.3158876, 0.3485199, 0.3280665, 0.3283358, 0.4513352, 0.2547335, 
    0.1966562, 0.2337262, 0.3784251, 0.319589,
  0.318678, 0.2907575, 0.4353006, 0.4587951, 0.4660494, 0.3911639, 0.2992977, 
    0.3683546, 0.5390061, 0.3618183, 0.340422, 0.3179289, 0.3399724, 
    0.3423811, 0.2678944, 0.3179853, 0.3425413, 0.3626739, 0.4473357, 
    0.3846121, 0.2592911, 0.2752655, 0.2436526, 0.2434438, 0.2704827, 
    0.1976757, 0.2437233, 0.3102323, 0.3664277,
  0.2726339, 0.2881332, 0.2687002, 0.2941478, 0.2886544, 0.2875988, 
    0.3088377, 0.3369588, 0.2590045, 0.2566081, 0.3114072, 0.3173644, 
    0.2626107, 0.2837943, 0.197045, 0.3254916, 0.2921102, 0.3400505, 
    0.2785714, 0.233351, 0.2218269, 0.1825484, 0.2628452, 0.2031492, 
    0.1220745, 0.2369647, 0.3038001, 0.3794714, 0.2689985,
  0.3025406, 0.2578746, 0.1915172, 0.2377308, 0.2615562, 0.3131321, 0.269966, 
    0.2708818, 0.259156, 0.1885011, 0.1670795, 0.1642048, 0.114303, 
    0.1982827, 0.218457, 0.1888582, 0.1972609, 0.1958684, 0.2019653, 
    0.2368026, 0.2584699, 0.2577851, 0.2069913, 0.2207482, 0.06046465, 
    0.2398834, 0.2219633, 0.2526382, 0.2951416,
  0.1911768, 0.08833166, 0.02962384, 0.09784523, 0.09982512, 0.1330479, 
    0.09977185, 0.1877315, 0.1358076, 0.1627905, 0.005649095, -3.069118e-05, 
    0.06003477, 0.1009086, 0.1421849, 0.1736151, 0.2179488, 0.2133487, 
    0.1700184, 0.1409962, 0.2213977, 0.2239187, 0.1493684, 0.001495673, 
    0.08535248, 0.1139402, 0.1784254, 0.1581714, 0.1319295,
  0.1478903, -9.002762e-05, 5.842059e-06, 0.04221128, 0.07895967, 0.03105053, 
    0.05869704, 0.1587264, 0.1467485, 0.0213717, -1.504213e-06, 0.0003941484, 
    0.1179972, 0.1300836, 0.1150687, 0.07404568, 0.1089988, 0.07711684, 
    0.03772684, 0.1318983, 0.1867765, 0.2158933, 0.0395707, 6.438325e-09, 
    4.829014e-05, 0.008086604, 0.05029776, 0.1654624, 0.3705601,
  6.752742e-05, 2.716965e-05, -0.0001567823, 0.02388858, 0.01823458, 
    0.03663019, 0.05802623, 0.07861313, 0.08243843, 0.02988307, 0.0403147, 
    0.03666848, 0.1930159, 0.07405822, 0.02643961, 0.04968857, 0.02492082, 
    0.01655334, 0.02399622, 0.03728926, 0.05010514, 0.002731411, 
    1.231097e-06, 0.01635216, 0.0007531762, 2.64029e-05, 0.05925507, 
    0.09492056, 0.009291681,
  0.01742628, 0.2009881, 0.01447157, 0.01821554, 0.03510544, 0.04862059, 
    0.01317665, 0.02351134, 0.06051271, 0.2241482, 0.04745111, 0.0256767, 
    0.0839546, 0.0258714, 0.02521322, 0.02221608, 0.02695997, 0.01366348, 
    0.01797176, 0.03059277, 0.003441748, 0.005919863, 0.01308835, 0.07418443, 
    0.02902451, 0.01380904, 0.02282184, 0.04641251, 0.005076258,
  0.0664176, 0.04742184, 0.02417996, 0.1191709, -8.015755e-05, 0.01431664, 
    0.02986146, 0.02602516, 0.01617425, 0.01666444, 0.0412744, 0.03154239, 
    0.02828294, 0.02023369, 0.03376102, 0.04364179, 0.08734541, 0.1692933, 
    0.1657862, 0.2191817, 0.06792111, 0.05251677, 0.2150456, 0.09934194, 
    0.02052012, 0.03722684, 0.07067759, 0.1142135, 0.1523652,
  1.942377e-07, 3.360459e-08, 1.554836e-08, -3.835821e-07, 6.405693e-08, 
    0.001143949, 0.1370556, 0.0688367, 0.2027473, 0.05508692, 0.02822849, 
    0.0393791, 0.02714648, 0.03958472, 0.03129152, 0.03997955, 0.083313, 
    0.04913042, 0.001242328, 0.02123628, 0.03260849, 0.1142363, 0.0159703, 
    0.01713955, 0.04451536, 0.03605332, 0.02957276, -9.045843e-06, 
    -1.886247e-06,
  -3.32313e-09, 1.73737e-06, 3.96715e-05, -1.457882e-10, 3.624435e-07, 
    -5.383745e-09, 0.008244977, 0.3256603, 0.3763051, 0.05047343, 0.09996053, 
    0.1000386, 0.08007468, 0.05720495, 0.04652388, 0.03373865, 0.08738792, 
    0.1020867, 0.01901331, 1.410429e-07, 0.00159962, 0.05328646, 0.04205328, 
    0.02285228, 0.025365, 0.03511102, 0.08052023, 0.02227779, 1.624951e-06,
  0.01805302, 0.004183786, 0.0008741936, 0.08947396, -1.856102e-05, 
    -4.042034e-05, 0.01337346, 0.0006561439, 0.001909143, 0.05052963, 
    0.1879836, 0.1084654, 0.1390231, 0.1344528, 0.2015656, 0.1625411, 
    0.2427867, 0.1872134, 0.0585688, -6.059175e-05, 0.0001604946, 
    0.0006985833, 0.0295552, 0.03140472, 0.1098391, 0.06146196, 0.104243, 
    0.1351888, 0.009911896,
  0.1484313, 0.2351802, 0.1504031, 0.06699857, 0.009919852, 0.03668221, 
    0.0396418, 0.1313398, 0.2458562, 0.1635319, 0.1385831, 0.1290786, 
    0.05355635, 0.2033221, 0.1028294, 0.06490649, 0.2063201, 0.2250841, 
    0.2784441, 0.04657647, 0.003161598, 0.003019089, 0.08739441, 0.2098483, 
    0.1670142, 0.2187184, 0.2271534, 0.2098966, 0.1693446,
  0.2742886, 0.2084701, 0.1660569, 0.1510207, 0.1235852, 0.1378039, 
    0.1493825, 0.1921882, 0.1696027, 0.2304935, 0.1822232, 0.3006926, 
    0.1402665, 0.2807521, 0.1873754, 0.3497812, 0.4127817, 0.5160901, 
    0.4454987, 0.08122839, 0.07108597, 0.1402906, 0.1708629, 0.2960465, 
    0.156087, 0.2813435, 0.3232573, 0.3454612, 0.2828215,
  0.3176924, 0.3308655, 0.3695665, 0.2162597, 0.2880859, 0.2271412, 
    0.3242964, 0.4062441, 0.3358578, 0.3454719, 0.3983073, 0.350794, 
    0.3557646, 0.3424458, 0.3589486, 0.2498749, 0.3478266, 0.2097135, 
    0.1891038, 0.2288731, 0.2037822, 0.2754504, 0.1844285, 0.1764602, 
    0.08007265, 0.320311, 0.1383458, 0.08359072, 0.1784174,
  0.2061406, 0.2991627, 0.2797614, 0.2454748, 0.3656213, 0.3751143, 0.310784, 
    0.319162, 0.331676, 0.3499606, 0.4366322, 0.5684802, 0.5425791, 
    0.6013916, 0.6384416, 0.4950944, 0.4148983, 0.3474496, 0.3896428, 
    0.3700874, 0.345486, 0.5075006, 0.432138, 0.3540598, 0.1628243, 
    0.2057407, 0.154589, 0.1467507, 0.1831356,
  0.2218536, 0.2178232, 0.2137928, 0.2097625, 0.2057321, 0.2017018, 
    0.1976714, 0.2232282, 0.2247619, 0.2262957, 0.2278294, 0.2293632, 
    0.2308969, 0.2324307, 0.2088432, 0.2135221, 0.2182011, 0.22288, 
    0.2275589, 0.2322378, 0.2369167, 0.2353394, 0.2331571, 0.2309748, 
    0.2287925, 0.2266102, 0.2244279, 0.2222456, 0.2250779,
  0.2319861, 0.1528771, 0.04487194, 0.03329983, 0.01099475, 0.0132857, 
    0.02670721, 0.0133094, 0.0004268664, 0.04191322, 0.07902863, 0.1003884, 
    0.1534792, 0.05605228, 0.07306233, 0.1139036, 0.1431372, 0.1571161, 
    0.2460111, 0.1720861, 0.3915298, 0.4242586, 0.3456203, 0.2385569, 
    0.2344858, 0.2148751, 0.2084989, 0.2201854, 0.2881954,
  0.2779225, 0.1974079, 0.2833397, 0.2525463, 0.3270012, 0.2212463, 
    0.1498815, 0.3489636, 0.314713, 0.3735997, 0.2860096, 0.1785485, 
    0.2372783, 0.3167688, 0.383996, 0.3555703, 0.2915743, 0.2320359, 
    0.5075208, 0.3246142, 0.3395763, 0.3919087, 0.373751, 0.4709439, 
    0.2354174, 0.2276386, 0.2581049, 0.3709224, 0.3438578,
  0.3997156, 0.4047867, 0.5796245, 0.4061339, 0.4346255, 0.4477029, 
    0.3347157, 0.4923192, 0.5408539, 0.2923409, 0.3222903, 0.3209074, 
    0.372612, 0.3659954, 0.2974879, 0.3173402, 0.4044757, 0.4436831, 
    0.4084992, 0.2703344, 0.2145408, 0.2288005, 0.2351509, 0.2626615, 
    0.2825634, 0.2258014, 0.311623, 0.3431002, 0.3522178,
  0.2618821, 0.2822523, 0.2889687, 0.3000815, 0.3134886, 0.3094531, 
    0.3250637, 0.3157555, 0.2451927, 0.2224077, 0.2854726, 0.3241076, 
    0.2328352, 0.2477829, 0.2643244, 0.2821929, 0.2858784, 0.3071727, 
    0.268178, 0.1802102, 0.217316, 0.2345539, 0.2767084, 0.2398758, 
    0.1236944, 0.2093365, 0.3333929, 0.3759376, 0.2958718,
  0.2636073, 0.2238273, 0.183752, 0.2449739, 0.2860025, 0.2876247, 0.3093684, 
    0.312274, 0.225313, 0.127912, 0.125, 0.1186037, 0.06988221, 0.2310765, 
    0.2595417, 0.1653874, 0.1881863, 0.2692636, 0.2043927, 0.2338516, 
    0.2120145, 0.2356213, 0.2073906, 0.2652436, 0.05371544, 0.2550209, 
    0.2191512, 0.2376131, 0.3166759,
  0.1720194, 0.07953159, 0.02776061, 0.07861541, 0.1442768, 0.1469343, 
    0.1988545, 0.3232725, 0.2540422, 0.09841222, 0.00107456, 0.0001444629, 
    0.04267589, 0.05181749, 0.1038213, 0.172724, 0.2056481, 0.2116976, 
    0.149214, 0.1239381, 0.1964054, 0.227777, 0.2061568, 0.007315591, 
    0.08514624, 0.1173813, 0.2133455, 0.1772578, 0.1076469,
  0.4084406, 0.0002471985, -1.650721e-05, 0.03587165, 0.08774106, 0.04541327, 
    0.07571287, 0.1344016, 0.1878604, 0.007675699, 1.3471e-07, 0.0001699819, 
    0.1263075, 0.1309206, 0.1975347, 0.08556699, 0.1108711, 0.08412619, 
    0.06078681, 0.222694, 0.1780369, 0.3768843, 0.2425046, 1.258899e-06, 
    -3.920425e-06, 0.006207218, 0.1406018, 0.1229965, 0.3700871,
  0.007594304, 0.0007597505, -7.565336e-05, 0.01066007, 0.03725466, 
    0.05096457, 0.07611136, 0.08744982, 0.08965314, 0.1324676, 0.04231384, 
    0.0647557, 0.2015965, 0.1014049, 0.04857178, 0.06910628, 0.0514388, 
    0.03563621, 0.04859322, 0.08734111, 0.1373569, 0.1230799, 6.206321e-05, 
    0.01335946, 0.0003261107, 4.429006e-06, 0.1009931, 0.09601559, 0.1359982,
  0.1053604, 0.2204237, 0.008618276, 0.02794293, 0.04283315, 0.05322414, 
    0.03329106, 0.02623959, 0.04965732, 0.2026378, 0.05178709, 0.0259821, 
    0.06964164, 0.02944807, 0.0277706, 0.02655594, 0.01877853, 0.01184006, 
    0.0152818, 0.04346776, 0.01915701, 0.0005925692, 0.01190452, 0.06722153, 
    0.01983791, 0.03048654, 0.04540748, 0.06083268, 0.03852948,
  0.06247296, 0.04346981, 0.01705027, 0.08732686, -2.359157e-05, 0.02032008, 
    0.02523003, 0.03479511, 0.01228392, 0.02272386, 0.01026138, 0.04264459, 
    0.03069927, 0.02423126, 0.03387312, 0.04240884, 0.07633666, 0.1502178, 
    0.1432242, 0.1756769, 0.06816897, 0.04720543, 0.22833, 0.09653641, 
    0.02517561, 0.03892518, 0.07060855, 0.1034634, 0.1287305,
  1.383196e-07, 2.98561e-08, 1.416041e-08, -4.948484e-09, 5.574837e-08, 
    0.02587039, 0.1006358, 0.06329712, 0.1824058, 0.03493738, 0.02492537, 
    0.04875072, 0.0326786, 0.04392087, 0.03668583, 0.04859802, 0.1576237, 
    0.1593884, 0.03797501, 0.03268973, 0.03636548, 0.1171254, 0.02638789, 
    0.0215165, 0.05445318, 0.06650557, 0.05057072, 0.0009497099, -7.010817e-07,
  -2.895886e-09, 3.465311e-07, 3.697634e-05, -4.476182e-10, 2.53746e-07, 
    -3.959703e-09, 0.003071258, 0.3415721, 0.3545658, 0.03903515, 0.131787, 
    0.1051945, 0.09135094, 0.05901154, 0.05434732, 0.04095528, 0.09717974, 
    0.1690339, 0.07669085, 6.235265e-07, 0.0005337929, 0.04884215, 
    0.04144914, 0.03428482, 0.04551912, 0.05434605, 0.09527759, 0.1017082, 
    9.898929e-07,
  0.02159568, 0.001180801, 0.0002970624, 0.1272159, -1.608167e-05, 
    -9.929929e-05, 0.01566284, 7.635226e-05, 0.0008192057, 0.04275525, 
    0.1670169, 0.1256929, 0.1807027, 0.1836037, 0.2395744, 0.1824869, 
    0.2823375, 0.2123879, 0.1153934, -7.279421e-05, 5.90566e-05, 
    0.0003786108, 0.03645785, 0.02328869, 0.1210037, 0.09033387, 0.1374741, 
    0.2654873, 0.04130443,
  0.1265581, 0.2102225, 0.1476431, 0.08728351, 0.008019388, 0.02841993, 
    0.01939928, 0.1294415, 0.2419176, 0.1817414, 0.1429732, 0.133441, 
    0.06051118, 0.2186435, 0.1448745, 0.1704777, 0.3104347, 0.2757827, 
    0.302967, 0.034741, 0.0029221, 0.0006526727, 0.08745437, 0.2023807, 
    0.1539251, 0.2505358, 0.2867682, 0.3339725, 0.2035347,
  0.3218615, 0.2034493, 0.1387257, 0.108031, 0.09808405, 0.1761879, 
    0.1528113, 0.1600256, 0.1363681, 0.2207311, 0.1774434, 0.296029, 
    0.154672, 0.2967215, 0.1866122, 0.3846293, 0.4007287, 0.4848422, 
    0.4549374, 0.05401909, 0.07303327, 0.170102, 0.2274781, 0.3279859, 
    0.2415419, 0.2387552, 0.4011776, 0.4473186, 0.2657445,
  0.4305277, 0.3122184, 0.3611661, 0.2428012, 0.3828928, 0.2900369, 
    0.3761185, 0.4215242, 0.2923328, 0.3313416, 0.3988425, 0.3514484, 
    0.3688932, 0.3638365, 0.3585359, 0.385557, 0.3619663, 0.24921, 0.244509, 
    0.237569, 0.2413876, 0.3297684, 0.2422395, 0.2031659, 0.088432, 0.305052, 
    0.108521, 0.08485487, 0.2698285,
  0.1986485, 0.3852159, 0.34642, 0.3425465, 0.4664841, 0.4693528, 0.4282862, 
    0.4667355, 0.5135611, 0.4724419, 0.5815826, 0.7188178, 0.7422069, 
    0.6746334, 0.6747417, 0.5992269, 0.4699979, 0.3585998, 0.497089, 
    0.4346443, 0.4454572, 0.5400915, 0.4489889, 0.3538875, 0.1784087, 
    0.1747873, 0.1543422, 0.1744916, 0.1553986,
  0.2261455, 0.2239303, 0.2217151, 0.2194999, 0.2172848, 0.2150696, 
    0.2128544, 0.2250108, 0.2267782, 0.2285457, 0.2303131, 0.2320805, 
    0.233848, 0.2356154, 0.2293059, 0.2314829, 0.2336598, 0.2358368, 
    0.2380138, 0.2401908, 0.2423677, 0.2379922, 0.236263, 0.2345338, 
    0.2328046, 0.2310754, 0.2293462, 0.2276169, 0.2279177,
  0.2264886, 0.1551652, 0.05184202, 0.04212821, 0.01895225, 0.018736, 
    0.02815455, 0.02191204, 0.0006386611, 0.0445007, 0.1013989, 0.1257714, 
    0.1539601, 0.02119054, 0.07709923, 0.1120756, 0.1634833, 0.1570061, 
    0.2101469, 0.1436848, 0.4488805, 0.4753069, 0.3635942, 0.2473581, 
    0.2204074, 0.2114036, 0.1706979, 0.2107434, 0.2861766,
  0.2325248, 0.1784082, 0.2611617, 0.1895905, 0.3030664, 0.216521, 
    0.09840874, 0.3206955, 0.3183063, 0.3744052, 0.2744224, 0.157959, 
    0.2144448, 0.2575015, 0.3925294, 0.4044546, 0.3229658, 0.2472436, 
    0.5749659, 0.3030736, 0.3463019, 0.3996734, 0.3902397, 0.4693846, 
    0.2171622, 0.2716204, 0.3199291, 0.3636511, 0.3605498,
  0.4667745, 0.4292441, 0.5661909, 0.322833, 0.3825285, 0.4831391, 0.3591862, 
    0.5770278, 0.4345677, 0.2190526, 0.2708177, 0.3191091, 0.4070643, 
    0.3925882, 0.3516241, 0.3490512, 0.4421273, 0.4503665, 0.3838557, 
    0.206192, 0.181871, 0.2037639, 0.2467386, 0.2590295, 0.2792338, 
    0.2494623, 0.3841562, 0.4071825, 0.4164895,
  0.3186041, 0.2806599, 0.249934, 0.3010924, 0.3212213, 0.3272196, 0.3305153, 
    0.281294, 0.2437993, 0.2257343, 0.2637866, 0.3378323, 0.2047634, 
    0.2012339, 0.2799575, 0.2748904, 0.2582926, 0.2854693, 0.2280056, 
    0.1676293, 0.1920289, 0.2602081, 0.2566198, 0.2529733, 0.123912, 
    0.2362573, 0.333391, 0.3674057, 0.3447431,
  0.1912299, 0.1640067, 0.1103073, 0.2355233, 0.2317363, 0.2271021, 
    0.2696467, 0.2096686, 0.1489192, 0.0775038, 0.1046657, 0.07220285, 
    0.03484988, 0.149967, 0.3142928, 0.1285275, 0.1234085, 0.2355404, 
    0.15909, 0.2058766, 0.1725218, 0.2030191, 0.2007953, 0.3181887, 
    0.0515084, 0.1713131, 0.171862, 0.2094432, 0.3191474,
  0.1493206, 0.1104473, 0.02360699, 0.05424031, 0.1453398, 0.1475153, 
    0.2147989, 0.2617012, 0.1978822, 0.02437361, 0.000299287, 4.387819e-05, 
    0.03619315, 0.03118498, 0.07666666, 0.178764, 0.16326, 0.2098265, 
    0.1199481, 0.09835198, 0.1683051, 0.2358965, 0.1961679, 0.0075522, 
    0.09712332, 0.125822, 0.1825786, 0.1494088, 0.1378266,
  0.502903, 0.003547288, -7.647688e-06, 0.04175977, 0.1226234, 0.04306547, 
    0.04153589, 0.06885428, 0.09751534, 0.002475125, 8.707789e-08, 
    4.693288e-05, 0.08955397, 0.0685703, 0.1881854, 0.1181142, 0.1244691, 
    0.129955, 0.1084891, 0.1197688, 0.07759992, 0.2741966, 0.5920517, 
    3.564481e-05, 0.0006261817, 0.007831793, 0.0691414, 0.0364592, 0.1730913,
  0.2858463, 0.01604691, -7.863058e-05, 0.007880521, 0.04750251, 0.06345949, 
    0.09828867, 0.08032104, 0.07393824, 0.07106802, 0.0391692, 0.05635639, 
    0.2061445, 0.1463386, 0.05685388, 0.04259961, 0.03924567, 0.02253992, 
    0.02412991, 0.03555922, 0.1322557, 0.4445216, 0.008147715, 0.005258351, 
    0.0001341858, 1.170276e-06, 0.07936912, 0.07405879, 0.3875839,
  0.1956388, 0.2001827, 0.003567952, 0.04124505, 0.04590249, 0.07639474, 
    0.1408424, 0.1002317, 0.03109356, 0.1659736, 0.08978578, 0.03330667, 
    0.06860279, 0.03320352, 0.02814057, 0.0279334, 0.02037934, 0.01640945, 
    0.01872958, 0.0251347, 0.08750406, 0.01489754, 0.01219144, 0.04359166, 
    0.007675121, 0.1067461, 0.08946295, 0.1203638, 0.08479298,
  0.05808715, 0.03989905, 0.01019254, 0.06890451, -8.133416e-06, 0.0166511, 
    0.0222315, 0.0641212, 0.01064037, 0.07745648, 0.002157137, 0.2086778, 
    0.03230683, 0.04896482, 0.04432501, 0.04828442, 0.08143718, 0.1344953, 
    0.12136, 0.1520009, 0.09050426, 0.05469641, 0.2189133, 0.09538728, 
    0.03981758, 0.05768454, 0.09148914, 0.1042487, 0.1071231,
  1.094068e-07, 2.735301e-08, 1.366895e-08, 5.313271e-09, 5.262294e-08, 
    0.06584411, 0.05409563, 0.05149533, 0.1606314, 0.02346419, 0.04163203, 
    0.04720666, 0.03654788, 0.09379604, 0.03581036, 0.06211292, 0.09140042, 
    0.2058357, 0.3032133, 0.06900523, 0.0347568, 0.1313778, 0.02576938, 
    0.02142127, 0.0681039, 0.1220936, 0.1500228, 0.02957046, -1.554909e-07,
  -2.503417e-09, -2.906327e-06, 0.0004420496, -3.645966e-09, 1.942401e-07, 
    -3.290271e-09, -0.0008057333, 0.375196, 0.3243988, 0.02873435, 0.1489487, 
    0.08974079, 0.1219361, 0.08320622, 0.05682812, 0.04500622, 0.07201132, 
    0.1931802, 0.2572089, 1.111721e-05, 0.0002155421, 0.04214358, 0.03685426, 
    0.1860771, 0.078839, 0.1199251, 0.1150847, 0.2113678, -6.232862e-05,
  0.02517345, 0.0001690171, 0.0001474356, 0.1591587, -3.266776e-05, 
    -4.886214e-05, 0.01119221, -4.248667e-06, -0.000107365, 0.03743853, 
    0.1373463, 0.1472415, 0.246457, 0.2372934, 0.2244001, 0.201843, 
    0.3140702, 0.1864435, 0.3506366, -0.0001231858, 2.251433e-05, 
    0.0002014724, 0.02597618, 0.05441, 0.1393992, 0.1449393, 0.2087551, 
    0.3352485, 0.08507932,
  0.130106, 0.1905105, 0.1272056, 0.08610677, 0.005568602, 0.03396323, 
    0.01336799, 0.1250095, 0.2268588, 0.1780258, 0.1198981, 0.1324854, 
    0.08140103, 0.2387696, 0.2966865, 0.3417298, 0.4763844, 0.3682488, 
    0.314372, 0.03026226, 0.002359066, 0.0009442521, 0.1003804, 0.191213, 
    0.1486705, 0.2916766, 0.3828365, 0.3457423, 0.1863387,
  0.3216123, 0.1943932, 0.1083678, 0.06678352, 0.08199108, 0.1428196, 
    0.1491053, 0.1045169, 0.1278826, 0.2016691, 0.1572887, 0.3006344, 
    0.158666, 0.3444476, 0.1652894, 0.4308704, 0.40804, 0.4522898, 0.4204584, 
    0.03392782, 0.05997763, 0.2043026, 0.2617832, 0.2958265, 0.3585684, 
    0.1945943, 0.4829279, 0.3678757, 0.2983642,
  0.5941242, 0.3572102, 0.3806266, 0.3561356, 0.4879822, 0.3983821, 
    0.4210292, 0.4682654, 0.2636334, 0.2464828, 0.4323105, 0.3705193, 
    0.3217295, 0.4201807, 0.4298477, 0.5757479, 0.4193172, 0.3361684, 
    0.256897, 0.2606342, 0.3366805, 0.4359217, 0.2915915, 0.244602, 
    0.1433733, 0.2661253, 0.102292, 0.1078935, 0.4917275,
  0.249034, 0.4453655, 0.4811785, 0.480479, 0.5501366, 0.5661417, 0.5547153, 
    0.6435935, 0.6604302, 0.6629851, 0.6327991, 0.7513901, 0.7513276, 
    0.6989174, 0.7070175, 0.6773685, 0.6804416, 0.5033669, 0.6207212, 
    0.5782614, 0.553632, 0.5972927, 0.4569865, 0.3513396, 0.199925, 
    0.1992901, 0.1586754, 0.2043173, 0.1835229,
  0.2194332, 0.218079, 0.2167247, 0.2153705, 0.2140163, 0.212662, 0.2113078, 
    0.2031297, 0.2059465, 0.2087633, 0.2115801, 0.2143969, 0.2172137, 
    0.2200305, 0.2175337, 0.2177089, 0.2178842, 0.2180594, 0.2182346, 
    0.2184098, 0.218585, 0.2085639, 0.2069261, 0.2052883, 0.2036505, 
    0.2020127, 0.200375, 0.1987372, 0.2205166,
  0.2210793, 0.1512545, 0.05277501, 0.05024358, 0.02364637, 0.02270303, 
    0.03658057, 0.02631328, 0.001555658, 0.04033508, 0.1216631, 0.1414724, 
    0.1457819, 0.003736347, 0.08614498, 0.1035421, 0.1536361, 0.1891899, 
    0.1944449, 0.1202002, 0.4528278, 0.4899669, 0.3579538, 0.2470862, 
    0.1914469, 0.2130374, 0.1897391, 0.2040055, 0.2895569,
  0.209057, 0.1538882, 0.2396119, 0.1384886, 0.2619072, 0.2026637, 
    0.05957842, 0.2994541, 0.3173063, 0.3784987, 0.2529213, 0.1554414, 
    0.1778371, 0.2146878, 0.4096633, 0.4147924, 0.3708692, 0.2840363, 
    0.5678635, 0.2921261, 0.35222, 0.3844711, 0.4336299, 0.4407883, 
    0.2131723, 0.3515756, 0.3771076, 0.382266, 0.3740441,
  0.4802067, 0.4131792, 0.4963623, 0.2656823, 0.3236355, 0.4523106, 
    0.3424361, 0.5918447, 0.2899893, 0.163309, 0.2274767, 0.2691454, 0.40091, 
    0.4576824, 0.3902637, 0.4035027, 0.4380378, 0.4593822, 0.3756752, 
    0.1691257, 0.1452045, 0.1916676, 0.2180084, 0.2383331, 0.2749691, 
    0.2627835, 0.4479056, 0.5252639, 0.4966257,
  0.2866364, 0.2858626, 0.2525252, 0.2851585, 0.3486048, 0.3336792, 
    0.3466417, 0.2520044, 0.237066, 0.2208497, 0.2455406, 0.3269748, 
    0.2287979, 0.199398, 0.1884325, 0.2207878, 0.195764, 0.2506085, 
    0.1838044, 0.1796004, 0.1611163, 0.2348609, 0.22727, 0.2269748, 0.133453, 
    0.250706, 0.2991565, 0.3354831, 0.3269089,
  0.1608624, 0.1199026, 0.08255218, 0.208351, 0.2067229, 0.1790595, 
    0.2055853, 0.1520045, 0.118939, 0.04215863, 0.07135533, 0.04438613, 
    0.01532035, 0.08598094, 0.317755, 0.1053959, 0.09192462, 0.1811688, 
    0.1417175, 0.1369909, 0.1463273, 0.207238, 0.1564276, 0.334667, 
    0.05987622, 0.1400688, 0.1483739, 0.1382481, 0.2979954,
  0.1132784, 0.03891709, 0.01852203, 0.02134018, 0.1723108, 0.1258564, 
    0.1056768, 0.1257684, 0.06499785, 0.008574555, 0.0001388684, 
    -5.479524e-05, 0.03445471, 0.01240452, 0.04600728, 0.1504543, 0.1202234, 
    0.1695542, 0.1192244, 0.0744475, 0.1707563, 0.1411252, 0.109162, 
    0.009174887, 0.1030423, 0.2130949, 0.1153765, 0.1123718, 0.1428335,
  0.2215774, 0.007526964, -3.138832e-05, 0.02021773, 0.1134313, 0.01590071, 
    0.01440837, 0.02007731, 0.02607895, 0.001573598, 5.889859e-08, 
    3.768522e-06, 0.05370314, 0.01698911, 0.1273314, 0.1429058, 0.1812705, 
    0.1176524, 0.03374379, 0.03780826, 0.02870327, 0.09878255, 0.3292091, 
    -0.0002202799, 2.805335e-05, 0.01100379, 0.0351988, 0.006127619, 
    0.05469352,
  0.5420231, 0.1413065, -2.067109e-05, 0.009135623, 0.03693789, 0.03382221, 
    0.04722093, 0.04566623, 0.02927469, 0.02859472, 0.04320617, 0.02343999, 
    0.1648693, 0.07694515, 0.01834064, 0.01337707, 0.009602583, 0.004575104, 
    0.006977547, 0.00671248, 0.03836609, 0.2289616, 0.2083042, 0.001473637, 
    7.408046e-05, 4.619978e-07, 0.01024901, 0.01768011, 0.1567731,
  0.2898913, 0.1721035, 0.001154258, 0.03921162, 0.04007157, 0.05969397, 
    0.03662624, 0.0327015, 0.02549149, 0.132774, 0.06498039, 0.04903829, 
    0.07014048, 0.02778537, 0.01234835, 0.007892037, 0.01610864, 0.01253156, 
    0.01678237, 0.02152119, 0.1406831, 0.2739292, 0.04698044, 0.01573529, 
    0.00216166, 0.03013242, 0.0237894, 0.0673569, 0.293103,
  0.04309926, 0.03474266, 0.006386847, 0.06584607, -9.638878e-07, 0.01142599, 
    0.02991557, 0.0245665, 0.0010971, 0.02935822, 0.0005446978, 0.09539152, 
    0.03269748, 0.1390661, 0.0427524, 0.03871326, 0.07379764, 0.1229886, 
    0.1145943, 0.1453699, 0.08183203, 0.1048454, 0.2440663, 0.07704174, 
    0.01673584, 0.0335136, 0.1047996, 0.1048342, 0.09044527,
  9.256978e-08, 2.598422e-08, 1.347872e-08, 2.681408e-09, 5.132123e-08, 
    0.08332757, 0.04998663, 0.0304745, 0.1383556, 0.02012572, 0.03480352, 
    0.02250316, 0.0164747, 0.04656127, 0.01732994, 0.01515751, 0.02142422, 
    0.08305494, 0.3187718, 0.2071459, 0.05481322, 0.1690299, 0.005707919, 
    0.001974582, 0.02034335, 0.06942112, 0.3123648, 0.04979131, -3.635254e-08,
  -2.23258e-09, -9.494724e-07, 0.0001710663, -8.474333e-08, 1.585238e-07, 
    -2.862766e-09, -0.004077656, 0.3895454, 0.3118362, 0.02495384, 0.1284584, 
    0.07411127, 0.08271868, 0.04689227, 0.068367, 0.1096909, 0.03129024, 
    0.1058712, 0.4926576, 0.001148691, 8.316948e-05, 0.04434218, 0.0287709, 
    0.07856277, 0.1164677, 0.1511488, 0.09444241, 0.2238463, -0.0004002665,
  0.01293192, -5.538453e-05, 0.0002199835, 0.210709, -4.79096e-05, 
    -7.811336e-06, 0.008915305, -2.300243e-05, -0.0002230705, 0.03262321, 
    0.09781422, 0.184615, 0.3086885, 0.2757984, 0.2613673, 0.2673817, 
    0.247404, 0.1674681, 0.3654712, -0.0001327793, 1.061053e-05, 8.78061e-05, 
    0.007854498, 0.02786263, 0.1412308, 0.1312279, 0.2206363, 0.2349931, 
    0.1241644,
  0.1239248, 0.156582, 0.1074441, 0.06867833, 0.00561319, 0.02990986, 
    0.005226764, 0.1269065, 0.2273491, 0.1635498, 0.1074458, 0.1021483, 
    0.1506856, 0.3548484, 0.4330391, 0.4292172, 0.4944791, 0.3829071, 
    0.3371648, 0.0356289, 0.0005646982, 0.00118954, 0.07096532, 0.1522288, 
    0.1516319, 0.3834878, 0.4021366, 0.3296777, 0.1712232,
  0.2899665, 0.1723235, 0.07418856, 0.05400492, 0.03884132, 0.1126103, 
    0.1496468, 0.07228979, 0.1094028, 0.1846564, 0.1458112, 0.3220617, 
    0.196133, 0.397867, 0.1789823, 0.4235289, 0.3630095, 0.4180436, 0.405913, 
    0.03040119, 0.05638308, 0.2241234, 0.2974966, 0.3216889, 0.5272945, 
    0.1611971, 0.4941421, 0.3377911, 0.327599,
  0.5930858, 0.3302039, 0.3576838, 0.2912976, 0.4785442, 0.399347, 0.4382308, 
    0.4866345, 0.1932101, 0.2302479, 0.4004664, 0.3464123, 0.2605751, 
    0.4145591, 0.4819983, 0.5003706, 0.4103732, 0.2793363, 0.3624401, 
    0.2783274, 0.4010621, 0.5514652, 0.2243009, 0.300599, 0.2408344, 
    0.2863501, 0.08464622, 0.197191, 0.6832088,
  0.3911152, 0.6021878, 0.556755, 0.6111425, 0.7079491, 0.725885, 0.6996928, 
    0.6624553, 0.6750206, 0.710443, 0.6604694, 0.7308382, 0.6815687, 
    0.721442, 0.7079294, 0.6812204, 0.7043176, 0.6662724, 0.6864986, 
    0.7309631, 0.7170885, 0.645188, 0.4636536, 0.3896973, 0.2176185, 
    0.1570067, 0.13687, 0.1873395, 0.2688971,
  0.1769586, 0.1744665, 0.1719744, 0.1694822, 0.1669901, 0.164498, 0.1620059, 
    0.1441463, 0.1498348, 0.1555233, 0.1612117, 0.1669002, 0.1725886, 
    0.1782771, 0.1667029, 0.1649702, 0.1632375, 0.1615047, 0.159772, 
    0.1580393, 0.1563066, 0.180759, 0.1792954, 0.1778318, 0.1763681, 
    0.1749045, 0.1734408, 0.1719772, 0.1789523,
  0.2225234, 0.1258079, 0.04366329, 0.04938712, 0.02300602, 0.02366212, 
    0.03263562, 0.02621369, 0.0011385, 0.00834681, 0.07935815, 0.1319846, 
    0.1640232, -0.002386998, 0.10537, 0.1276823, 0.1878855, 0.2356975, 
    0.1938485, 0.1447783, 0.4634927, 0.4983656, 0.3156655, 0.2206676, 
    0.2145985, 0.2217141, 0.2298651, 0.1909505, 0.2842912,
  0.179964, 0.1257677, 0.2175043, 0.09102583, 0.209201, 0.1788194, 
    0.02537654, 0.2873979, 0.3131845, 0.3645, 0.2242358, 0.1608121, 
    0.1458766, 0.1860468, 0.4309639, 0.4411516, 0.4126325, 0.3282302, 
    0.5499821, 0.3455589, 0.3924672, 0.3960823, 0.443276, 0.4120362, 
    0.2372831, 0.4258753, 0.4195642, 0.4318696, 0.381159,
  0.4881479, 0.4052791, 0.3938821, 0.2227838, 0.263503, 0.385134, 0.3294426, 
    0.4797338, 0.1854257, 0.1178112, 0.1838133, 0.2265126, 0.3860097, 
    0.4507671, 0.3929003, 0.4114313, 0.4463061, 0.4620653, 0.3317788, 
    0.1408612, 0.1147686, 0.1622341, 0.193858, 0.2232383, 0.2737554, 
    0.2963606, 0.4817503, 0.6156617, 0.5711349,
  0.2431296, 0.2422796, 0.2616653, 0.2984576, 0.3373204, 0.3635394, 
    0.3205916, 0.2282517, 0.2059389, 0.1940389, 0.1916642, 0.2368142, 
    0.1650555, 0.2160746, 0.1616221, 0.1731261, 0.1348886, 0.190076, 
    0.153289, 0.1630685, 0.1334759, 0.2034263, 0.1870544, 0.1874928, 
    0.1260278, 0.2127871, 0.2439662, 0.2828439, 0.2719786,
  0.1551923, 0.08237422, 0.06555662, 0.1713302, 0.1828679, 0.1647468, 
    0.1700252, 0.09865238, 0.09033587, 0.01896494, 0.04544576, 0.02566851, 
    0.007359643, 0.05240079, 0.2625669, 0.08288787, 0.08463715, 0.133356, 
    0.08987422, 0.1023685, 0.1289987, 0.1835525, 0.1292325, 0.332249, 
    0.04430975, 0.1149569, 0.1272642, 0.09814522, 0.2680317,
  0.04644864, 0.01231764, 0.01266238, 0.009364198, 0.1595524, 0.09667318, 
    0.06773283, 0.04152406, 0.02660954, 0.004120635, 4.298098e-05, 
    -0.000213881, 0.03057268, 0.006167401, 0.03333502, 0.1164113, 0.0893449, 
    0.1563676, 0.1093514, 0.06642365, 0.1227845, 0.09343622, 0.03474513, 
    0.008695932, 0.09507672, 0.177766, 0.073857, 0.06178974, 0.06122776,
  0.08393507, 0.01205376, -4.049546e-05, 0.004989647, 0.03941343, 
    0.001869653, 0.005927878, 0.004394839, 0.007938578, 0.0005569739, 
    4.386392e-08, 7.194552e-07, 0.03747188, 0.003657117, 0.09888265, 
    0.1250939, 0.09980065, 0.02810273, 0.007485882, 0.009478038, 0.005016294, 
    0.03799345, 0.1425924, 0.01760594, 1.285634e-06, 0.01951462, 0.02314033, 
    0.00141466, 0.01742521,
  0.2584836, 0.3198299, 9.809799e-05, 0.01431595, 0.007868021, 0.01312916, 
    0.02049034, 0.02108297, 0.007106571, 0.00598965, 0.02201444, 0.003986406, 
    0.1053898, 0.03981064, 0.002167665, 0.008583827, 0.001049307, 
    0.0003871942, 0.0006552655, 0.000703107, 0.007225624, 0.08045878, 
    0.1790533, 0.0001678545, 2.599903e-05, 1.92849e-07, -0.0007388562, 
    0.004238017, 0.05302827,
  0.1598037, 0.146513, 0.0005019414, 0.02095776, 0.01334897, 0.02260717, 
    0.007114804, 0.01472461, 0.02946471, 0.1003515, 0.02204509, 0.02359382, 
    0.06305849, 0.00930583, 0.002390269, 0.0004687927, 0.004477446, 
    0.004945697, 0.0128573, 0.0198597, 0.08166628, 0.5066212, 0.1764762, 
    0.006562217, 0.0006308304, 0.004589578, 0.003667941, 0.009100824, 
    0.1524545,
  0.02049919, 0.03540662, 0.004280149, 0.06702043, -2.572667e-07, 0.0043893, 
    0.04018657, 0.004747821, -0.00356898, 0.005254934, 0.0001860938, 
    0.02021594, 0.01675518, 0.02170674, 0.01361488, 0.01750622, 0.04627686, 
    0.09242909, 0.0834605, 0.1309459, 0.02400197, 0.02510732, 0.2780567, 
    0.05222006, 0.002458188, 0.01056281, 0.04736896, 0.08824484, 0.07557668,
  8.148976e-08, 2.462968e-08, 1.334509e-08, 9.621928e-10, 5.026634e-08, 
    0.06153939, 0.03320451, 0.01722413, 0.1393596, 0.01497124, 0.01660663, 
    0.005993909, 0.003906539, 0.01587449, 0.002162896, 0.002053646, 
    0.00348833, 0.02697297, 0.192716, 0.4541268, 0.1350682, 0.1441416, 
    0.0003719425, -0.002829109, 0.003835418, 0.01733548, 0.1407654, 
    0.1329713, 3.392971e-09,
  -2.032311e-09, -8.609003e-07, 0.0006996202, -8.186267e-08, 1.354092e-07, 
    -2.567198e-09, -0.005942712, 0.3820289, 0.302201, 0.01795082, 0.138886, 
    0.03337513, 0.04977347, 0.02027529, 0.04386699, 0.02198013, 0.007466774, 
    0.05265877, 0.2627046, 0.1830832, 2.458343e-05, 0.03433178, 0.01774929, 
    0.02807954, 0.02637897, 0.03247288, 0.04328547, 0.09785764, -0.0005202723,
  0.006400552, 4.302779e-05, 0.0002971105, 0.2534246, -4.464046e-05, 
    -2.052113e-06, 0.007884861, -2.857469e-06, -0.0001909771, 0.02677514, 
    0.07605463, 0.1649504, 0.4490281, 0.3726432, 0.3217667, 0.3699764, 
    0.2150168, 0.1474079, 0.2475041, -0.0002088623, 1.1701e-05, 2.620978e-05, 
    0.003203988, 0.04306032, 0.1323595, 0.1358704, 0.1386135, 0.1905136, 
    0.1144439,
  0.09497923, 0.1329404, 0.09336012, 0.05454857, 0.002581341, 0.02034489, 
    0.001793424, 0.1387012, 0.2087109, 0.1493022, 0.09897043, 0.09376621, 
    0.2857061, 0.5052311, 0.5685627, 0.579573, 0.4755039, 0.3151774, 
    0.3458633, 0.04372916, 0.0001368751, 0.0001247205, 0.05295581, 0.118493, 
    0.1516096, 0.4017203, 0.3563994, 0.2773823, 0.1410371,
  0.2360108, 0.1519531, 0.04814681, 0.04495944, 0.02278918, 0.1028557, 
    0.1425205, 0.05327145, 0.0935978, 0.17564, 0.1450715, 0.365542, 
    0.2857406, 0.4376176, 0.1939485, 0.4169627, 0.3238889, 0.3951668, 
    0.431945, 0.02603995, 0.04606145, 0.2453681, 0.3353638, 0.3582186, 
    0.600078, 0.1283842, 0.4681817, 0.2909803, 0.2854538,
  0.4250672, 0.2297654, 0.3008842, 0.2002779, 0.4035875, 0.3188328, 
    0.4249202, 0.4305864, 0.1652001, 0.1799978, 0.3421756, 0.2993615, 
    0.2204162, 0.3396415, 0.431752, 0.4356177, 0.3507829, 0.2388891, 
    0.3704189, 0.2897797, 0.4196864, 0.5518346, 0.1891166, 0.3152097, 
    0.549227, 0.2832068, 0.06786768, 0.2680752, 0.6048401,
  0.5100804, 0.7020515, 0.4656218, 0.6054718, 0.7123379, 0.7190766, 
    0.7068973, 0.6559977, 0.576192, 0.6207303, 0.5980371, 0.6712949, 
    0.6251838, 0.6822287, 0.702995, 0.6803842, 0.6706604, 0.6965725, 
    0.6867449, 0.8424646, 0.7951532, 0.6151071, 0.4795403, 0.4203099, 
    0.2746988, 0.1424941, 0.108597, 0.1564364, 0.3022997,
  0.09321445, 0.09017443, 0.08713441, 0.08409438, 0.08105436, 0.07801434, 
    0.07497431, 0.0712798, 0.07708111, 0.08288242, 0.08868372, 0.09448504, 
    0.1002863, 0.1060876, 0.1016139, 0.1017404, 0.1018668, 0.1019933, 
    0.1021198, 0.1022462, 0.1023727, 0.1392143, 0.1363266, 0.1334388, 
    0.1305511, 0.1276633, 0.1247755, 0.1218878, 0.09564647,
  0.2157615, 0.1073802, 0.03268296, 0.04393383, 0.01716501, 0.01545439, 
    0.02222181, 0.02231413, 0.00064896, 0.0008062187, 0.04364469, 0.07749972, 
    0.1822377, -0.002041949, 0.135399, 0.209927, 0.2746392, 0.2720376, 
    0.2017617, 0.1959104, 0.4864536, 0.5122522, 0.2754667, 0.2059021, 
    0.2394598, 0.2837904, 0.2857885, 0.1519183, 0.2437097,
  0.1706351, 0.1035688, 0.2044765, 0.05843979, 0.1475384, 0.1617802, 
    0.01391966, 0.2633772, 0.2801388, 0.3261128, 0.2149888, 0.1683217, 
    0.1252413, 0.1493256, 0.4545659, 0.4758011, 0.4619617, 0.3859374, 
    0.5723547, 0.3980808, 0.4269266, 0.3986459, 0.4525716, 0.4077904, 
    0.2662159, 0.4813324, 0.4640801, 0.4786383, 0.4010173,
  0.5129005, 0.4390399, 0.3109707, 0.1686679, 0.2104091, 0.3146917, 
    0.3412347, 0.3831826, 0.1275954, 0.08474235, 0.1317228, 0.1883277, 
    0.3453754, 0.4010362, 0.3513747, 0.3789299, 0.409965, 0.4039115, 
    0.2748652, 0.107239, 0.09016301, 0.1330874, 0.1667118, 0.173734, 
    0.2621376, 0.3089549, 0.4696128, 0.6186343, 0.5984827,
  0.1996825, 0.1981326, 0.236181, 0.2774985, 0.2909231, 0.3309613, 0.2838294, 
    0.1964858, 0.1717531, 0.1589824, 0.1335635, 0.1692168, 0.1035827, 
    0.1900312, 0.1329916, 0.1296301, 0.07556769, 0.1441426, 0.1228068, 
    0.1207417, 0.1031856, 0.1515141, 0.1399999, 0.1525759, 0.09559571, 
    0.1583763, 0.2114928, 0.23509, 0.2281357,
  0.1398241, 0.05229494, 0.05807288, 0.1238439, 0.1701607, 0.1463015, 
    0.1273321, 0.06862254, 0.06103724, 0.007514812, 0.02286141, 0.01471949, 
    0.003673784, 0.03549886, 0.2100614, 0.06239392, 0.06342713, 0.1055606, 
    0.07210886, 0.08462131, 0.112696, 0.1601283, 0.1005072, 0.3173601, 
    0.0282973, 0.08251704, 0.1002392, 0.06511192, 0.2298095,
  0.01522521, 0.00593036, 0.008235137, 0.003029926, 0.09857711, 0.07410528, 
    0.03935007, 0.02234051, 0.01471196, 0.002562555, 5.882302e-06, 
    -0.0005862793, 0.02230796, 0.003181303, 0.02920422, 0.08195654, 
    0.06631248, 0.1377021, 0.07629646, 0.03589802, 0.07875063, 0.0495591, 
    0.01289317, 0.003517148, 0.09823788, 0.07490186, 0.03805903, 0.03565872, 
    0.0242268,
  0.03798886, 0.0209251, -3.894925e-05, 0.001465166, 0.009719239, 
    0.0002470635, 0.00232181, 0.001229244, 0.003305069, 0.0002636242, 
    3.69737e-08, 3.912746e-07, 0.02987363, 0.001567077, 0.06255889, 
    0.0842467, 0.04414487, 0.008142623, 0.002483537, 0.003888917, 
    0.001276904, 0.01548337, 0.06576424, 0.01062156, -5.82805e-07, 
    0.03020135, 0.01301773, 0.0007086693, 0.007183707,
  0.1193478, 0.211126, 0.0002206204, 0.03334019, 0.001826259, 0.004328323, 
    0.006916525, 0.009535177, 0.001454291, 0.0002850064, 0.01405528, 
    0.0006391095, 0.06129192, 0.0127718, 0.0002633709, 0.0122323, 
    0.0002688942, 3.438425e-05, 0.0002702157, 0.0002916207, 0.002581901, 
    0.03019799, 0.07074293, 2.352848e-05, 9.771203e-06, 1.100376e-07, 
    -0.0005120937, 0.00161929, 0.01942893,
  0.04972155, 0.1249659, 0.0003583705, 0.008489945, 0.002370173, 0.009786384, 
    0.002002696, 0.003107974, 0.04285963, 0.08896288, 0.00252678, 
    0.006191934, 0.03661286, 0.001802035, 0.0003890148, 2.118606e-05, 
    0.0001823402, 8.218395e-05, 0.0008866282, 0.006259728, 0.01542237, 
    0.2161631, 0.1090672, 0.002442115, 0.000215512, 0.001645066, 
    0.0009999354, 0.003053184, 0.04136696,
  0.01004269, 0.03332308, 0.002239177, 0.06962706, -1.075392e-07, 
    0.0006695931, 0.05118126, 0.0008204428, -0.004540467, 0.001606148, 
    1.65561e-05, 0.006625955, 0.004508275, 0.005150355, 0.003107368, 
    0.002222956, 0.02338792, 0.07549981, 0.03974187, 0.07055479, 0.006068093, 
    0.003539357, 0.3097384, 0.04141546, 0.000249719, 0.003377534, 0.01299303, 
    0.03604157, 0.07004012,
  7.505343e-08, 2.309511e-08, 1.325657e-08, 2.50417e-10, 4.88121e-08, 
    0.01744941, 0.01608348, 0.001629605, 0.1332213, 0.00760442, 0.002455364, 
    0.001116846, 0.0003155459, 0.007864338, 0.0001151144, 0.0006122802, 
    0.00128926, 0.008804858, 0.07543562, 0.2469499, 0.03682791, 0.1068408, 
    3.523232e-05, -0.002277616, 0.0007302302, 0.004794205, 0.04679691, 
    0.09693832, -2.389049e-09,
  -1.903762e-09, 1.536862e-07, 0.000936618, -6.718481e-07, 1.205207e-07, 
    -2.368029e-09, -0.006499924, 0.352153, 0.2819744, 0.0125168, 0.1005939, 
    0.01036934, 0.02056386, 0.01146056, 0.02281871, 0.007547477, 
    0.0009620583, 0.03736104, 0.1070693, 0.2746966, 1.088433e-05, 0.02351535, 
    0.01302504, 0.008501871, 0.007162706, 0.00981926, 0.01166158, 0.03802432, 
    -0.0004852653,
  0.003593649, -2.023093e-05, 0.0001049531, 0.2638905, -5.436263e-05, 
    -1.070601e-06, 0.008368054, 1.893398e-07, -0.0001675612, 0.01946666, 
    0.07123785, 0.1487914, 0.4338206, 0.3948629, 0.3661378, 0.38237, 
    0.1361191, 0.1018033, 0.1640161, -0.0007439697, 9.098007e-06, 
    -1.515114e-05, 0.005697222, 0.057366, 0.1346132, 0.1048561, 0.09341135, 
    0.1325857, 0.0895128,
  0.06765085, 0.1095615, 0.0826694, 0.04607796, 0.002373209, 0.01292048, 
    0.0006064108, 0.1276888, 0.1877452, 0.1427203, 0.08536198, 0.09535513, 
    0.4087495, 0.6565937, 0.7147828, 0.6430963, 0.4259178, 0.2562534, 
    0.3253357, 0.04165479, 4.940854e-05, -8.652531e-06, 0.04202942, 
    0.09859849, 0.1614248, 0.4056754, 0.2883541, 0.2295482, 0.1433803,
  0.181822, 0.1285878, 0.03284876, 0.03221713, 0.01546241, 0.09443845, 
    0.1314124, 0.04457521, 0.0809787, 0.1678739, 0.1316092, 0.3737388, 
    0.3067161, 0.43865, 0.2114421, 0.3674018, 0.3037301, 0.3663627, 
    0.4014817, 0.02366446, 0.03965693, 0.2306048, 0.3021201, 0.3679486, 
    0.5068977, 0.1160551, 0.4146235, 0.2313281, 0.2180479,
  0.3039865, 0.1689863, 0.2844602, 0.1824895, 0.3288232, 0.3746251, 
    0.3498567, 0.3741567, 0.1578103, 0.1421586, 0.3080526, 0.2675615, 
    0.1993694, 0.274324, 0.3430479, 0.3615046, 0.2903653, 0.2235668, 
    0.3386626, 0.277408, 0.4437075, 0.5098943, 0.1962668, 0.2683085, 
    0.7087664, 0.2477659, 0.06512231, 0.2341339, 0.4308046,
  0.5871084, 0.6274559, 0.3563057, 0.5319147, 0.6198515, 0.6289653, 0.620536, 
    0.5281453, 0.4558566, 0.5096145, 0.5346089, 0.6291518, 0.5902197, 
    0.6283798, 0.685581, 0.6694548, 0.6499802, 0.6422168, 0.6672978, 
    0.8162898, 0.7457654, 0.5399797, 0.5112402, 0.4133072, 0.2526478, 
    0.1273604, 0.07121637, 0.1284977, 0.346772,
  0.02515564, 0.02247247, 0.0197893, 0.01710612, 0.01442295, 0.01173978, 
    0.009056605, 0.02104703, 0.0259025, 0.03075798, 0.03561345, 0.04046892, 
    0.0453244, 0.05017987, 0.05924453, 0.06041449, 0.06158445, 0.06275441, 
    0.06392436, 0.06509433, 0.06626429, 0.07915778, 0.07581552, 0.07247327, 
    0.069131, 0.06578874, 0.06244648, 0.05910422, 0.02730218,
  0.1819369, 0.09167586, 0.007878589, 0.00639797, 0.0003699312, 0.007201408, 
    0.0038371, 0.0051479, 0.0006867303, 0.0006980027, 0.01308207, 0.04790327, 
    0.1912086, -0.001561808, 0.1652866, 0.3795421, 0.3416577, 0.2682271, 
    0.1832055, 0.238589, 0.5381192, 0.5591047, 0.225848, 0.1811682, 
    0.2658515, 0.369457, 0.2918483, 0.1109469, 0.1893347,
  0.1693224, 0.08955872, 0.2014332, 0.04007291, 0.1033487, 0.1389208, 
    0.006351597, 0.2059734, 0.2160109, 0.2723083, 0.1881202, 0.1657093, 
    0.1036712, 0.1083223, 0.4783421, 0.4694469, 0.4239219, 0.365342, 
    0.4892024, 0.3960948, 0.4119941, 0.3787076, 0.4631843, 0.3584358, 
    0.227603, 0.4742145, 0.4997609, 0.490186, 0.4120464,
  0.4658175, 0.3953427, 0.2336133, 0.1149981, 0.1421818, 0.2347403, 
    0.3080807, 0.3121637, 0.08926174, 0.05564203, 0.09158901, 0.1461615, 
    0.2917698, 0.3327039, 0.2762367, 0.28588, 0.3238715, 0.309396, 0.2092615, 
    0.07776739, 0.06738151, 0.1073337, 0.1241789, 0.13206, 0.2429547, 
    0.2735773, 0.404303, 0.5441833, 0.5349618,
  0.157125, 0.1542612, 0.1857922, 0.236894, 0.2408983, 0.2642897, 0.2397338, 
    0.144549, 0.1334293, 0.1189672, 0.08816694, 0.108399, 0.0608954, 
    0.1377897, 0.1166978, 0.08909708, 0.04115235, 0.1039068, 0.09651613, 
    0.08611918, 0.07401151, 0.104906, 0.09657041, 0.1261696, 0.07108539, 
    0.1177331, 0.1724367, 0.1839802, 0.1755201,
  0.1059823, 0.03164252, 0.04969173, 0.0880857, 0.1261353, 0.1014331, 
    0.08247622, 0.04358784, 0.03685419, 0.00318716, 0.01011001, 0.007384835, 
    0.001553834, 0.02301043, 0.1528459, 0.04921655, 0.04709719, 0.08551884, 
    0.06167149, 0.06706288, 0.09186076, 0.1335447, 0.06466538, 0.2900077, 
    0.0193275, 0.06226789, 0.06742375, 0.0400414, 0.1806589,
  0.00838776, 0.003854583, 0.005000647, 0.001267791, 0.06041776, 0.04467537, 
    0.02036976, 0.01318123, 0.009937176, 0.001831748, 4.555846e-06, 
    -0.0007780634, 0.01390661, 0.001076852, 0.02158601, 0.05128593, 
    0.04834314, 0.09668162, 0.04381564, 0.01688441, 0.04422235, 0.03079856, 
    0.006769518, 0.001474545, 0.09420034, 0.039078, 0.02144799, 0.02064464, 
    0.01338824,
  0.02178903, 0.02096215, -2.799744e-05, 0.0007512706, 0.002009387, 
    0.0001019744, 0.0005609472, 0.0005252208, 0.001787149, 0.0001797177, 
    3.246063e-08, -1.453809e-08, 0.01799082, 0.0009092276, 0.02830725, 
    0.0381097, 0.01658745, 0.003228507, 0.001257169, 0.001951642, 
    0.0006112464, 0.007808404, 0.03734058, 0.004193428, -5.954694e-07, 
    0.03950939, 0.0070932, 0.0004471896, 0.003861562,
  0.06558208, 0.09600563, 9.071498e-05, 0.04870217, 0.0009061974, 
    0.001789809, 0.00219938, 0.003784586, 0.000314872, -0.0004576493, 
    0.01502118, 0.0003081248, 0.03124456, 0.004084218, 9.713606e-05, 
    0.0093037, 0.0001553249, 1.775479e-05, 0.0001470756, 0.0001598826, 
    0.001334217, 0.0148959, 0.03747357, 6.118642e-05, 2.686572e-06, 
    1.811182e-07, -0.0005173807, 0.0008332666, 0.009908102,
  0.02400096, 0.1135885, 0.0003294748, 0.003164024, 0.000131931, 0.003688388, 
    0.001107067, 0.001197935, 0.03835987, 0.079793, 0.0004825453, 
    0.004719061, 0.01660788, 0.0004416171, 7.313539e-05, 5.739312e-06, 
    4.067894e-05, 1.766624e-05, 7.146146e-05, 0.0005632505, 0.004896871, 
    0.09198236, 0.05393021, 0.0009936769, 0.0001316866, 0.0008807606, 
    0.0005605645, 0.001615116, 0.01859768,
  0.006006565, 0.03809988, 0.001006331, 0.06172979, -5.23505e-08, 
    4.181532e-05, 0.04230513, 0.0002908205, -0.002604995, 0.0008336286, 
    5.200671e-08, 0.003470897, 0.001915971, 0.002629153, 0.0006884777, 
    0.0003184381, 0.009111304, 0.05790262, 0.01528348, 0.03128687, 
    0.00174417, 0.0007200642, 0.261048, 0.0390384, 0.0001184315, 0.002065259, 
    0.003818451, 0.01408949, 0.05298483,
  6.948392e-08, 2.219832e-08, 1.320094e-08, 6.730656e-11, 4.778123e-08, 
    0.003048142, 0.003330054, -1.724959e-05, 0.1233404, 0.002108525, 
    0.000455822, 0.0004750936, 7.249894e-05, 0.003589987, 4.477959e-05, 
    0.0002936553, 0.0007048161, 0.004553109, 0.03204649, 0.1285404, 
    0.01262564, 0.08723667, 1.560634e-05, -0.001723547, 0.0003423356, 
    0.002191245, 0.02047382, 0.03988089, 4.700414e-09,
  -1.810302e-09, 2.47399e-07, 0.001207925, -7.017129e-07, 1.100943e-07, 
    -2.224599e-09, -0.006232414, 0.3265839, 0.2545747, 0.0067346, 0.05484083, 
    0.003136473, 0.006855939, 0.005405731, 0.01221428, 0.004150875, 
    0.0003737084, 0.01913103, 0.05155957, 0.1997521, 1.290681e-06, 
    0.01756447, 0.009356701, 0.004352866, 0.003372211, 0.004832909, 
    0.005708992, 0.01891807, -0.0003272619,
  0.002610822, -8.09143e-05, 2.191207e-05, 0.2513993, -4.192513e-05, 
    -1.506522e-07, 0.007626079, 5.074553e-07, -0.0001332843, 0.01414945, 
    0.05898472, 0.1475821, 0.3775699, 0.3202767, 0.2993493, 0.2571067, 
    0.06424253, 0.05110678, 0.09840461, -0.001410263, 6.152749e-06, 
    -1.60089e-05, 0.004411853, 0.04906235, 0.09616178, 0.06965167, 
    0.05498121, 0.09022639, 0.08598813,
  0.04229379, 0.09014335, 0.05995191, 0.03459802, 0.001044618, 0.006502996, 
    0.0002419924, 0.1127952, 0.1619128, 0.1332707, 0.07371625, 0.09616854, 
    0.487723, 0.7026047, 0.7025685, 0.6282674, 0.3603213, 0.2073745, 
    0.2789319, 0.0358132, 2.662112e-05, -1.494039e-05, 0.03846183, 
    0.08227956, 0.1350568, 0.4221778, 0.2199123, 0.1867962, 0.1293313,
  0.1440057, 0.1102736, 0.02247199, 0.02658996, 0.01101385, 0.08438477, 
    0.1088623, 0.0381262, 0.07379024, 0.161671, 0.1152469, 0.3538028, 
    0.3003027, 0.4030818, 0.2403403, 0.3171403, 0.2815582, 0.3236719, 
    0.3400937, 0.01947526, 0.03265565, 0.211275, 0.264317, 0.3697405, 
    0.4007651, 0.1278269, 0.3593596, 0.1812257, 0.1656812,
  0.2337383, 0.1310126, 0.246926, 0.1510971, 0.2868474, 0.3623608, 0.2758364, 
    0.3160507, 0.1440039, 0.1154626, 0.2766135, 0.2321791, 0.180052, 
    0.238098, 0.2839297, 0.3007158, 0.2635186, 0.2285383, 0.2986235, 0.25483, 
    0.4372549, 0.4905431, 0.1922877, 0.2510428, 0.6668595, 0.2177759, 
    0.05800059, 0.21788, 0.3206188,
  0.5508924, 0.5318123, 0.2784961, 0.4371156, 0.5068032, 0.5121281, 
    0.5396092, 0.4294172, 0.3679709, 0.4198015, 0.4134665, 0.500256, 
    0.4980842, 0.5400562, 0.6091133, 0.6003119, 0.5928191, 0.5671698, 
    0.6113928, 0.715028, 0.6900213, 0.4193621, 0.4753344, 0.410316, 
    0.2122017, 0.0927941, 0.04133598, 0.1048799, 0.3769285,
  0.01440501, 0.01380268, 0.01320036, 0.01259803, 0.01199571, 0.01139338, 
    0.01079106, 0.02012765, 0.0234531, 0.02677855, 0.03010399, 0.03342944, 
    0.03675489, 0.04008034, 0.04353616, 0.04380924, 0.04408232, 0.0443554, 
    0.04462848, 0.04490156, 0.04517464, 0.04467896, 0.04168276, 0.03868655, 
    0.03569035, 0.03269415, 0.02969794, 0.02670174, 0.01488687,
  0.1586076, 0.06623261, 0.001942633, 0.001561152, 0.0005651913, 0.001652003, 
    0.001445772, 0.00131015, 2.537547e-05, 0.0008195419, 0.006973812, 
    0.03011072, 0.09720844, -0.001414366, 0.2421139, 0.3867514, 0.2754426, 
    0.3346552, 0.1686206, 0.3203866, 0.5626186, 0.5877253, 0.2031748, 
    0.1623367, 0.2548318, 0.4689552, 0.2628969, 0.08585817, 0.1564041,
  0.1829372, 0.06835436, 0.1766426, 0.03069893, 0.0767692, 0.1230552, 
    0.004885595, 0.1456578, 0.1456581, 0.2154946, 0.1597793, 0.1267643, 
    0.09017797, 0.0914905, 0.4628915, 0.4428509, 0.3800761, 0.3283251, 
    0.4335019, 0.3676099, 0.3700953, 0.3633264, 0.4703068, 0.3000465, 
    0.1989613, 0.4549689, 0.4843868, 0.4389616, 0.3770683,
  0.3711624, 0.3363437, 0.1858609, 0.08027911, 0.1028975, 0.1819497, 
    0.2769186, 0.2553832, 0.06371297, 0.03880606, 0.06682949, 0.1110914, 
    0.2346191, 0.2631828, 0.2049866, 0.2053101, 0.2382414, 0.2417964, 
    0.1632382, 0.05814687, 0.05170463, 0.08297245, 0.0969792, 0.09800987, 
    0.2118187, 0.2320603, 0.3438004, 0.4505256, 0.4415579,
  0.1216957, 0.117756, 0.1343143, 0.1896809, 0.2078783, 0.2085376, 0.1973003, 
    0.107925, 0.1036372, 0.08725625, 0.05708724, 0.06647343, 0.03684441, 
    0.08560582, 0.09803695, 0.06224297, 0.02493505, 0.06894784, 0.07637084, 
    0.05986666, 0.04854858, 0.06816535, 0.0604731, 0.1031751, 0.04969602, 
    0.07306448, 0.1318908, 0.140061, 0.1303945,
  0.07541437, 0.01789716, 0.03671475, 0.05637767, 0.07060104, 0.05354299, 
    0.04987656, 0.02825693, 0.02030112, 0.00181407, 0.005717854, 0.004472079, 
    0.0008605976, 0.01212021, 0.1118479, 0.03505262, 0.0291261, 0.06341096, 
    0.05018377, 0.0457385, 0.06570921, 0.09724689, 0.03974745, 0.2564924, 
    0.01316977, 0.04556668, 0.04261258, 0.02231928, 0.1312753,
  0.00572994, 0.002865077, 0.002902774, 0.0007555357, 0.03390429, 0.02160916, 
    0.01132016, 0.008601642, 0.007484035, 0.001422231, 9.315355e-07, 
    -0.0004818169, 0.007762699, 0.0003961996, 0.01181813, 0.02987077, 
    0.0282493, 0.05334235, 0.02396982, 0.007634686, 0.02066724, 0.01730134, 
    0.004626014, 0.0007626608, 0.08160982, 0.01791216, 0.01205981, 
    0.009537647, 0.009315408,
  0.01464631, 0.01812429, -1.749994e-05, 0.0004832023, 4.848198e-05, 
    5.79964e-05, 0.0001971485, 0.0003042383, 0.001142323, 0.0001353745, 
    2.937672e-08, -5.214154e-06, 0.007795785, 0.000631407, 0.01147565, 
    0.01240676, 0.007287207, 0.002052073, 0.0007788575, 0.00115426, 
    0.0003701274, 0.004818222, 0.02521549, 0.002363232, -4.404551e-07, 
    0.0296794, 0.003713242, 0.0003212069, 0.002462186,
  0.04270234, 0.04746733, 2.897364e-05, 0.04878031, 0.0005965917, 
    0.0004909221, 0.001004595, 0.001298148, 0.0001357379, 7.844888e-05, 
    0.01063722, 0.0001948451, 0.01269152, 0.001673406, 6.449244e-05, 
    0.005161725, 0.0001047812, 1.151578e-05, 9.584668e-05, 0.0001041292, 
    0.0008320631, 0.00909153, 0.02406587, 4.237632e-05, 1.042907e-06, 
    6.092446e-08, -0.0001537486, 0.0005148558, 0.006244367,
  0.01502807, 0.09514298, 0.0001914136, 0.001425192, 5.838121e-05, 
    0.001504808, 0.0007249287, 0.0006620468, 0.02765153, 0.0737143, 
    0.0002602394, 0.002988665, 0.006698226, 0.000141805, 3.352007e-05, 
    3.063062e-06, 2.078803e-05, 7.669657e-06, 3.267061e-05, 0.0001939661, 
    0.002709399, 0.05070264, 0.0353687, 0.0009605263, 7.17716e-05, 
    0.0005727654, 0.0003693592, 0.001036672, 0.01121806,
  0.004904113, 0.02978032, 0.0005481953, 0.0495911, -1.461058e-08, 
    1.567327e-05, 0.02382563, 0.0001813623, -0.001015338, 0.0005182374, 
    9.837833e-07, 0.002195156, 0.0006739269, 0.001437106, 0.0001962563, 
    6.250538e-05, 0.003381324, 0.02923357, 0.005455681, 0.0129715, 
    0.0008957706, 0.0003072738, 0.2124562, 0.04152987, 7.289094e-05, 
    0.001034835, 0.001137458, 0.00562332, 0.03715186,
  6.622857e-08, 2.162718e-08, 1.316963e-08, -5.575919e-11, 4.711288e-08, 
    0.001381126, -0.0008834354, -2.99433e-05, 0.1035149, 0.0003137537, 
    0.0002460644, 0.0002428423, 3.315879e-05, 0.001634481, 2.410063e-05, 
    0.0001734731, 0.000461527, 0.00240209, 0.0180626, 0.07274783, 
    0.006029329, 0.07077621, 9.141832e-06, -0.001255872, 0.0002127273, 
    0.001351033, 0.01185017, 0.02079315, 4.338599e-09,
  -1.747448e-09, 2.674449e-07, 0.0004324049, -1.310553e-06, 1.026337e-07, 
    -2.123266e-09, -0.00574256, 0.300305, 0.2212254, 0.00336423, 0.0214162, 
    0.001133327, 0.00266526, 0.001730756, 0.005498083, 0.002775982, 
    0.0002176108, 0.0074319, 0.03107546, 0.1652217, -1.725305e-06, 
    0.01148644, 0.004557579, 0.002803778, 0.002171465, 0.00303314, 
    0.003592173, 0.01153606, -0.0002571957,
  0.001679943, -0.0001152555, -2.819577e-05, 0.2315067, -4.022582e-05, 
    -2.51007e-07, 0.006738297, 5.941016e-07, -0.0001010139, 0.01143902, 
    0.04827124, 0.1303083, 0.3021037, 0.2476224, 0.1893459, 0.1605811, 
    0.02645722, 0.02428697, 0.06364504, -0.002293649, 4.382616e-06, 
    -4.567641e-06, 0.006885787, 0.04963331, 0.0516651, 0.03931852, 
    0.02778333, 0.04899093, 0.08746844,
  0.02154119, 0.06663384, 0.03956797, 0.02035962, 0.0005075421, 0.003066243, 
    0.0001234638, 0.1068602, 0.1388594, 0.1242258, 0.06380412, 0.08202519, 
    0.4580899, 0.6673773, 0.6475275, 0.5567111, 0.2763746, 0.1435465, 
    0.2039916, 0.03396699, 1.510499e-05, -4.622071e-06, 0.03256899, 
    0.06548431, 0.1081776, 0.397166, 0.1606733, 0.1351527, 0.0938818,
  0.09986918, 0.09046515, 0.01722242, 0.01905316, 0.007867479, 0.07301765, 
    0.09037045, 0.03162999, 0.06376079, 0.1414136, 0.09720715, 0.3141266, 
    0.2869544, 0.3435406, 0.2261669, 0.2570834, 0.243449, 0.2668701, 
    0.2643265, 0.01301328, 0.02570168, 0.19787, 0.223464, 0.3395252, 
    0.3228303, 0.1131981, 0.2488891, 0.1201414, 0.1014319,
  0.1615719, 0.09896921, 0.2100056, 0.1254092, 0.2284777, 0.3081576, 
    0.2122329, 0.2644456, 0.1219383, 0.08760925, 0.2385202, 0.1907123, 
    0.1555246, 0.2211164, 0.2374446, 0.2527848, 0.21913, 0.2177045, 
    0.2744621, 0.2540354, 0.377947, 0.4622189, 0.1728325, 0.2279034, 
    0.5915294, 0.1838086, 0.0603452, 0.1887635, 0.2454639,
  0.4958204, 0.4632038, 0.2125311, 0.3513593, 0.4112421, 0.4112504, 
    0.4325193, 0.3425487, 0.2786122, 0.3075175, 0.2689007, 0.3336248, 
    0.3097084, 0.3403885, 0.4194879, 0.4273908, 0.4558899, 0.441808, 
    0.5236931, 0.5976725, 0.6121768, 0.3367011, 0.4273322, 0.4000974, 
    0.179661, 0.06700943, 0.02994668, 0.08493348, 0.3721734,
  0.003076577, 0.003191179, 0.003305781, 0.003420383, 0.003534985, 
    0.003649588, 0.00376419, 0.01048744, 0.01328853, 0.01608963, 0.01889073, 
    0.02169183, 0.02449292, 0.02729402, 0.03491892, 0.03480327, 0.03468761, 
    0.03457196, 0.0344563, 0.03434064, 0.03422499, 0.02177066, 0.01897062, 
    0.01617057, 0.01337053, 0.01057049, 0.007770444, 0.004970401, 0.002984896,
  0.06755415, 0.03215805, 0.00207996, 0.001998526, 6.610027e-05, 0.001805818, 
    0.001556749, 0.001303023, -2.814307e-06, 8.467206e-05, 0.003408546, 
    0.02286398, 0.06924308, -0.000749802, 0.2897987, 0.2845693, 0.2428338, 
    0.3457178, 0.1356919, 0.3725578, 0.5846575, 0.6087115, 0.1845135, 
    0.1538688, 0.2225132, 0.4266412, 0.2653883, 0.05312473, 0.08418812,
  0.1689648, 0.05499205, 0.154594, 0.02277465, 0.0620441, 0.1114696, 
    0.004249717, 0.1106027, 0.06808143, 0.163751, 0.1411598, 0.08803605, 
    0.0849181, 0.08495806, 0.4359057, 0.4041598, 0.3426897, 0.3039074, 
    0.4025588, 0.3345257, 0.3382658, 0.3501832, 0.4479232, 0.2668644, 
    0.1874077, 0.4265053, 0.4410213, 0.3573096, 0.3166667,
  0.3179598, 0.2905777, 0.1559855, 0.06353942, 0.07808559, 0.1511251, 
    0.24373, 0.2212799, 0.05115723, 0.02965332, 0.0525162, 0.09054253, 
    0.1909881, 0.2145409, 0.1604296, 0.1600537, 0.1907824, 0.203528, 
    0.133623, 0.0458985, 0.04271424, 0.07187849, 0.08226428, 0.07794511, 
    0.183997, 0.210213, 0.3064044, 0.3788051, 0.3779491,
  0.09715022, 0.09751786, 0.1006402, 0.1610187, 0.1860104, 0.1757295, 
    0.1674243, 0.08619077, 0.08566803, 0.06743556, 0.04091861, 0.04601769, 
    0.02249362, 0.05918997, 0.06925217, 0.04330488, 0.01696619, 0.05085066, 
    0.06353623, 0.04244428, 0.03540905, 0.04980003, 0.04129143, 0.0943592, 
    0.03655891, 0.05134371, 0.1023246, 0.1139036, 0.1039003,
  0.05117298, 0.01213053, 0.02529527, 0.03722747, 0.04207625, 0.03148473, 
    0.02990089, 0.01724364, 0.01282613, 0.001290302, 0.003814202, 
    0.003157205, 0.0006409381, 0.00719641, 0.08469774, 0.02239478, 
    0.01793529, 0.04481261, 0.03852283, 0.03043022, 0.04648271, 0.07331707, 
    0.02514912, 0.2317163, 0.01076112, 0.03435588, 0.02914637, 0.01250316, 
    0.0943383,
  0.004425881, 0.002323758, 0.001816214, 0.0005516507, 0.02072161, 0.0115135, 
    0.007397854, 0.006337684, 0.006104141, 0.001179554, 6.794622e-07, 
    -0.0001571667, 0.005369527, 0.0002881527, 0.006931884, 0.01485224, 
    0.01431484, 0.02570096, 0.01321824, 0.004117906, 0.0107627, 0.009930765, 
    0.003584434, 0.0005643782, 0.06634276, 0.01052661, 0.006357643, 
    0.005675247, 0.007320189,
  0.01108273, 0.01518509, -1.205825e-05, 0.0003356455, -0.0002068915, 
    4.003181e-05, 0.0001015517, 0.0002108276, 0.0008352475, 0.000110467, 
    2.739249e-08, -8.215216e-06, 0.003564067, 0.0004861497, 0.005578043, 
    0.005644064, 0.004133772, 0.001535667, 0.0005583517, 0.0007915557, 
    0.000260254, 0.003445494, 0.01913354, 0.001622554, -3.156472e-07, 
    0.02195339, 0.001879369, 0.0002536984, 0.001793415,
  0.0315952, 0.02861645, 9.687263e-06, 0.03925369, 0.0004441041, 
    0.0001927138, 0.0006382657, 0.0005098429, 8.795202e-05, 0.0002442626, 
    0.006346165, 0.0001399644, 0.005929643, 0.0008959979, 4.732385e-05, 
    0.00241277, 7.89256e-05, 8.437345e-06, 7.112853e-05, 7.747441e-05, 
    0.0006061128, 0.00647207, 0.01774277, 5.926147e-05, 1.10388e-06, 
    5.602114e-08, -4.47469e-05, 0.000367649, 0.004542062,
  0.01098592, 0.09214244, 0.0001594805, 0.0007854028, 3.749371e-05, 
    0.0006647903, 0.0005409364, 0.0004563977, 0.02342069, 0.0699326, 
    0.0001752434, 0.001390707, 0.003030504, 8.451708e-05, 2.251871e-05, 
    2.172366e-06, 1.407449e-05, 4.726615e-06, 1.994669e-05, 0.0001139556, 
    0.001853095, 0.03410849, 0.02654575, 0.002854394, 0.001530956, 
    0.0004250385, 0.000276025, 0.0007578628, 0.007938353,
  0.003913717, 0.01759123, 0.000518582, 0.03864427, 5.364412e-09, 
    1.060044e-05, 0.01216051, 0.0001334483, -0.0004730374, 0.000374993, 
    1.162995e-06, 0.001587573, 0.0002942361, 0.0008853254, 0.0001166758, 
    4.753171e-05, 0.001209882, 0.01234211, 0.002336172, 0.005406524, 
    0.0004183143, 0.0001997968, 0.1707741, 0.04236683, 5.235498e-05, 
    0.000517439, 0.0004294172, 0.002395438, 0.01838106,
  6.294461e-08, 2.125421e-08, 1.317281e-08, -1.310008e-10, 4.65871e-08, 
    0.0008317912, -0.000933072, 1.358674e-05, 0.08889995, 9.804705e-05, 
    0.0001727423, 0.0001355199, 2.224011e-05, 0.0008933995, 1.711085e-05, 
    0.0001203812, 0.0003414848, 0.001718945, 0.01231933, 0.04976323, 
    0.004033287, 0.0604698, 6.483811e-06, -0.0009366079, 0.0001535007, 
    0.0009685845, 0.008160696, 0.01273822, 4.178288e-09,
  -1.704998e-09, 2.68378e-07, 0.0002798708, -1.183821e-06, 9.769198e-08, 
    -2.048463e-09, -0.005282034, 0.2746808, 0.1933337, 0.001867967, 
    0.01036689, 0.0005913057, 0.001415644, 0.000962334, 0.003261857, 
    0.00208422, 0.0001348858, 0.003792163, 0.02087952, 0.1424864, 
    -3.109868e-06, 0.009327173, 0.003767739, 0.00206006, 0.001596501, 
    0.002189446, 0.002596015, 0.008162369, -0.0001818364,
  0.001556302, -0.0001353791, -3.000237e-05, 0.2077731, -3.928515e-05, 
    -1.975209e-07, 0.005709487, 6.087983e-07, -8.022076e-05, 0.00865487, 
    0.04401819, 0.1112258, 0.2330813, 0.1914749, 0.1324888, 0.1080664, 
    0.01239497, 0.01327422, 0.03992562, -0.002588552, 4.096647e-06, 
    -6.511581e-06, 0.007173912, 0.048378, 0.03308328, 0.02242886, 0.01547233, 
    0.02733831, 0.06997886,
  0.01196873, 0.0501937, 0.03152561, 0.01382384, 0.0002937763, 0.001749778, 
    8.17218e-05, 0.1024316, 0.1232644, 0.1141881, 0.06513634, 0.06445173, 
    0.4098991, 0.5869526, 0.5526419, 0.4224938, 0.1887506, 0.09620309, 
    0.1402504, 0.03283243, 9.298625e-06, -2.24284e-06, 0.0251953, 0.0607085, 
    0.08911201, 0.3423793, 0.120427, 0.0981304, 0.06547157,
  0.06033167, 0.08008588, 0.01717073, 0.01467256, 0.008459886, 0.06401355, 
    0.08048051, 0.0256444, 0.06553876, 0.1229424, 0.08602753, 0.2819113, 
    0.27856, 0.2739457, 0.1672223, 0.1828238, 0.2045801, 0.2240648, 
    0.2058033, 0.00879615, 0.01814808, 0.1949863, 0.1786273, 0.3134731, 
    0.2620561, 0.08276836, 0.1749481, 0.07792729, 0.06283972,
  0.101143, 0.06898404, 0.175988, 0.09966841, 0.1854847, 0.2667624, 
    0.1733573, 0.2225324, 0.101072, 0.0639564, 0.1997363, 0.1603088, 
    0.1350767, 0.198504, 0.2028352, 0.2040027, 0.1900574, 0.2096136, 
    0.2701274, 0.2920586, 0.3013446, 0.4533423, 0.146442, 0.2060254, 
    0.5129471, 0.1612116, 0.07289734, 0.1556058, 0.1867775,
  0.4631027, 0.4038187, 0.1712752, 0.2816049, 0.3455299, 0.330696, 0.3635961, 
    0.2943248, 0.2301764, 0.2339593, 0.200274, 0.2457545, 0.2140678, 
    0.2327769, 0.2885511, 0.3230245, 0.3602076, 0.3666757, 0.4341118, 
    0.5134634, 0.5319925, 0.2868362, 0.3775854, 0.376669, 0.1605045, 
    0.05426076, 0.02130946, 0.07166918, 0.3428094,
  0.00251772, 0.002610245, 0.002702771, 0.002795297, 0.002887823, 
    0.002980349, 0.003072874, 0.007439569, 0.009584879, 0.01173019, 
    0.0138755, 0.01602081, 0.01816612, 0.02031143, 0.02308439, 0.02318056, 
    0.02327674, 0.02337291, 0.02346908, 0.02356525, 0.02366142, 0.01587232, 
    0.01353831, 0.0112043, 0.008870291, 0.006536283, 0.004202275, 
    0.001868266, 0.002443699,
  0.02413257, 0.01362237, 0.001610231, 0.001994044, 6.271788e-05, 
    0.002247852, 0.001294923, 0.001417566, -7.201451e-08, 2.231896e-05, 
    0.001194994, 0.01922123, 0.052627, -0.0005582937, 0.3473766, 0.1989453, 
    0.2159666, 0.443215, 0.1995608, 0.3971588, 0.57159, 0.6010036, 0.2068193, 
    0.1491499, 0.2404572, 0.3695017, 0.2368624, 0.05181314, 0.05192043,
  0.1548069, 0.05981247, 0.1316558, 0.01982953, 0.0378407, 0.1000297, 
    0.003915902, 0.1091584, 0.05914097, 0.1335454, 0.1378228, 0.08277874, 
    0.07983862, 0.08144537, 0.4174607, 0.3871186, 0.3204322, 0.2880497, 
    0.3844919, 0.3232054, 0.3347097, 0.3414311, 0.4157644, 0.2379998, 
    0.191627, 0.403122, 0.3923418, 0.3238436, 0.2925253,
  0.2948301, 0.2627243, 0.1422395, 0.0556166, 0.0666393, 0.1371654, 
    0.2291609, 0.2091007, 0.04559918, 0.02549914, 0.0449307, 0.07958332, 
    0.1686804, 0.1898754, 0.1346563, 0.1379974, 0.1679381, 0.182772, 
    0.117713, 0.03970866, 0.03819112, 0.06417644, 0.07342658, 0.0682907, 
    0.178787, 0.2095608, 0.2864258, 0.3503492, 0.3537256,
  0.08548409, 0.08331092, 0.08458756, 0.1336644, 0.1623672, 0.1545331, 
    0.1455764, 0.07405267, 0.07756082, 0.05802305, 0.03426846, 0.03708941, 
    0.01678496, 0.04513952, 0.05218281, 0.03230871, 0.01350968, 0.03696458, 
    0.0452396, 0.03251455, 0.02888005, 0.04103025, 0.032798, 0.1219083, 
    0.03031193, 0.04244018, 0.08759976, 0.09966604, 0.09206702,
  0.03787005, 0.01019642, 0.01583887, 0.02690212, 0.02948437, 0.02135183, 
    0.02167268, 0.0124829, 0.009593373, 0.001073557, 0.002950394, 
    0.002576441, 0.0005547538, 0.005325146, 0.08204552, 0.01554743, 
    0.01241152, 0.03309793, 0.02787722, 0.02260125, 0.03645723, 0.05629104, 
    0.01887457, 0.2344375, 0.008056356, 0.02554546, 0.0222178, 0.008804473, 
    0.06957389,
  0.003758746, 0.002044239, 0.001427558, 0.0004618182, 0.0121273, 
    0.007224244, 0.005352741, 0.005316753, 0.005345774, 0.001024942, 
    3.358686e-07, -0.0001951786, 0.004858272, 0.0002443462, 0.004908608, 
    0.008381683, 0.007793383, 0.01406352, 0.008566121, 0.002630982, 
    0.006971386, 0.007110579, 0.003053483, 0.0004755844, 0.06735875, 
    0.006293558, 0.004266297, 0.004119995, 0.006255601,
  0.009350574, 0.01276958, -9.029225e-06, 0.0002974088, -0.0003868925, 
    3.258766e-05, 7.671538e-05, 0.0001748738, 0.0007049391, 9.833032e-05, 
    2.619213e-08, -4.382852e-06, 0.002223254, 0.0004161661, 0.003586891, 
    0.003569601, 0.002920125, 0.001268573, 0.0004594545, 0.0006210259, 
    0.0002128737, 0.002820402, 0.01617391, 0.001273411, -3.56604e-06, 
    0.02339302, 0.001211425, 0.0002188184, 0.001486893,
  0.02610676, 0.02052554, 8.303704e-06, 0.03109789, 0.0003617068, 
    0.0001224369, 0.0005070097, 0.000327903, 6.923491e-05, 0.0001805341, 
    0.004379731, 0.0001182236, 0.003634322, 0.0006633806, 3.949525e-05, 
    0.001405295, 7.004795e-05, 7.293814e-06, 6.102496e-05, 6.630522e-05, 
    0.0005036846, 0.005304026, 0.01464322, 0.0004771075, 2.957256e-07, 
    7.155653e-08, -4.771582e-05, 0.0003040265, 0.003758109,
  0.009000781, 0.1611914, 0.001871167, 0.0005181127, 3.019718e-05, 
    0.000417336, 0.0004372592, 0.0003513607, 0.03804984, 0.09403976, 
    0.0001400831, 0.0008173565, 0.001960103, 5.943514e-05, 1.840784e-05, 
    1.923083e-06, 1.155452e-05, 3.69783e-06, 1.647009e-05, 8.505203e-05, 
    0.001471542, 0.0265661, 0.02201442, 0.03491353, 0.04545336, 0.0003570957, 
    0.0002337538, 0.0006257682, 0.006319559,
  0.0200651, 0.0211114, 0.0003826352, 0.03871886, 1.791095e-08, 8.806719e-06, 
    0.008573242, 9.841767e-05, -0.001275446, 0.000311243, 1.08782e-06, 
    0.001285694, 0.0001993247, 0.0006780296, 9.103526e-05, 4.042058e-05, 
    0.0007082815, 0.006935151, 0.001502079, 0.003340923, 0.0002768329, 
    0.0001517233, 0.236228, 0.04454385, 4.135871e-05, 0.0003653983, 
    0.0003192737, 0.001530932, 0.01836646,
  6.155516e-08, 2.110518e-08, 1.316759e-08, -1.299974e-10, 4.705262e-08, 
    0.0006452436, -0.001014026, -4.885117e-06, 0.1555363, -0.0006442457, 
    0.0001404776, 9.444966e-05, 1.788701e-05, 0.0006424912, 1.456997e-05, 
    9.855009e-05, 0.0002874284, 0.001419359, 0.009758247, 0.03930058, 
    0.003048742, 0.05730137, 5.427153e-06, -0.001594503, 0.0001279338, 
    0.0007957161, 0.006516635, 0.009623515, 4.095308e-09,
  -1.678999e-09, 2.659764e-07, 0.0008363627, -8.079367e-07, 9.502278e-08, 
    -1.997317e-09, -0.004955373, 0.2812352, 0.1966867, 0.001782132, 
    0.006820245, 0.000435891, 0.001030135, 0.0006646012, 0.002031653, 
    0.001725185, 0.0001014273, 0.002644669, 0.01647192, 0.1280987, 
    -2.636102e-06, 0.03419846, 0.0184285, 0.001699375, 0.00130668, 
    0.001768131, 0.002084409, 0.00662155, -0.0001537726,
  0.001924418, -0.0001939003, -0.0001301281, 0.2025385, -5.57064e-05, 
    -1.689193e-07, 0.005093263, 5.999786e-07, -6.969806e-05, 0.007284335, 
    0.07589346, 0.07637186, 0.1699851, 0.1429133, 0.09004801, 0.06986239, 
    0.008204821, 0.008797213, 0.0225246, -0.003037678, 3.930386e-06, 
    0.0002763623, 0.02748546, 0.03732208, 0.02501594, 0.0149877, 0.01091071, 
    0.0171413, 0.05320453,
  0.007778344, 0.06424566, 0.04127526, 0.01169779, 0.0002021329, 0.00118453, 
    5.879516e-05, 0.1165231, 0.1305036, 0.1270171, 0.160685, 0.07956099, 
    0.340954, 0.4783461, 0.4594554, 0.3453732, 0.1385516, 0.07263625, 
    0.1017757, 0.03370296, 6.899691e-06, -1.971473e-06, 0.03339836, 
    0.1019091, 0.08724506, 0.2857254, 0.09250827, 0.07631671, 0.04661389,
  0.04091773, 0.09438886, 0.03350297, 0.01476824, 0.02184696, 0.08548821, 
    0.08803369, 0.03846458, 0.1012358, 0.1349301, 0.1036019, 0.3231288, 
    0.2782285, 0.24085, 0.114838, 0.1426595, 0.2089746, 0.2040125, 0.2008622, 
    0.01305688, 0.01567861, 0.2291368, 0.1373574, 0.3180656, 0.2146599, 
    0.07076719, 0.1372526, 0.05409785, 0.04558471,
  0.072253, 0.04396041, 0.1693096, 0.07776784, 0.1453563, 0.2402429, 
    0.1764914, 0.2198751, 0.0999937, 0.05941672, 0.1879192, 0.1637146, 
    0.1392508, 0.1857055, 0.1854392, 0.1666828, 0.1806544, 0.1933675, 
    0.2642766, 0.314489, 0.2525932, 0.4614947, 0.1426676, 0.1975265, 
    0.4590755, 0.1468557, 0.1140348, 0.142925, 0.1544996,
  0.4063033, 0.3516046, 0.1499672, 0.2247386, 0.2906412, 0.2746036, 
    0.3126978, 0.2560959, 0.1999191, 0.1971035, 0.1693098, 0.2075167, 
    0.1734633, 0.1832475, 0.2306126, 0.2707394, 0.3080624, 0.3214787, 
    0.3613315, 0.4575265, 0.4778801, 0.254878, 0.344133, 0.3695568, 
    0.1472706, 0.04823688, 0.01756029, 0.06503953, 0.3045586,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -9.781895e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -9.885714e-06, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.43997e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0.0001514288, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -8.355161e-05, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001253358, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.000810859, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.000238726, -3.81824e-05, 0, 0, 0, 0, 0, 0, 
    0, 0, -1.487063e-05, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.415689e-05, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0.0003479914, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -9.050902e-05, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0006095336, -3.235338e-05, 0, 0, 
    -3.316172e-05, 0, 0, -7.500415e-06, 0, 0.005095, -2.26638e-05, 0, 
    0.0002422386, 0, -4.364201e-05, 0.0002868087, 0,
  0, 0, 0, 0, 0, 0, -1.74537e-05, 0, 0, 0, 0.004059867, -9.442141e-05, 
    -3.837243e-07, 0, 0, 0, 0, 0, 0, 0, -0.0001768327, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.973796e-10, 0, 0, 0, 0, 0, 0, 0, 0, 
    -6.262018e-05, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0004337995, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0.001233235, 0, 0, 0, 0, 0, 0, 5.138428e-05, 
    -4.78798e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0.0006657381, -1.610592e-05, 0, 0, -4.373563e-06, -2.153974e-05, 
    1.965432e-05, -1.387993e-05, -3.728524e-05, 0, -8.308553e-06, 
    -9.813235e-05, 3.272267e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  -6.610934e-05, 0, 0, 0, 0, 0, 0, 0, 0, 3.935179e-06, 0, 0, 0.002504257, 
    0.0004726522, 0.0007227199, -1.303952e-06, -9.653578e-05, 0.000344757, 0, 
    0.00131345, 0, 0.010941, 0.0002540387, -4.298045e-07, 0.001293074, 0, 
    -0.0002123452, 0.0007198182, 0.0006097128,
  0, 0, 0, 0, 0, 0, -9.04902e-05, -8.90617e-06, 0, -1.331032e-05, 
    0.008458287, 8.612727e-06, 0.0002503446, 0, 0, 0, 0, 0, 0, -1.741212e-06, 
    0.0001259312, -0.000219726, 0, 0, 0, -5.057812e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.000201177, 0.001651591, -8.003853e-05, 0, 
    9.122416e-05, -1.657848e-05, 0, -1.781441e-05, 0, 0, 0, 0, 0, 
    -0.000110207, 0, 0, 0, 0, -7.207611e-06, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001543228, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -3.918361e-07, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0.001983645, 0, 0, 0, 0, 0, 0.007056042, 0.001448675, 
    -6.870827e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0.001419238, -6.336319e-05, 0, 0, -1.312071e-05, -7.513326e-05, 
    -0.0002686432, -9.420764e-05, -0.000111076, 3.452051e-05, -3.819416e-05, 
    -0.0002187346, 7.131127e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.117189e-05, 0, 
    0, 0, 0, 0,
  -9.152051e-05, 0, 0, 0, 0, 0, 0, 0, 0, -1.171252e-05, 0, 0, 0.009056948, 
    0.003039004, 0.001995071, 0.004223988, 0.000148776, 0.0005454406, 0, 
    0.01283345, -7.037379e-05, 0.02224298, 0.0003635887, -2.915038e-05, 
    0.002213437, 3.464592e-07, 0.00183402, 0.001295546, 0.00129986,
  0, 0, 0, 0, 0, 0, -3.954801e-05, -8.899254e-06, 0, -7.320675e-05, 
    0.01685633, 0.002637776, 0.001889014, -2.16438e-05, -1.022657e-06, 0, 0, 
    0, 0, -2.176515e-06, 0.001145471, -0.0004740151, 0, 0, -2.853336e-08, 
    -0.0002311228, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.001071485, 0.003305552, 4.520986e-05, 9.977557e-05, 
    0.0002155102, -9.078297e-05, 2.261364e-05, -7.551741e-05, -1.685627e-05, 
    0, 0, 0, 0, 0.0002414956, 0, 0, 0, 0, -3.939225e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -5.002381e-05, 0, 0.01157395, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -1.564226e-05, -8.228149e-06, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -4.241067e-05, -1.827434e-06, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -4.912456e-06, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0.002609965, 3.432697e-05, 0, 0, 0, 0, 0.01098061, 
    0.006281023, -5.840028e-05, -2.051602e-05, 0, 0, 0, 0, 0, 0, 0, 
    4.555988e-05, 0, 0, 0, 0, 0,
  0, 0.005841359, 0.0001715, 0, 0, -1.749431e-05, -3.271816e-05, 0.001084648, 
    -0.0002683986, 0.0006171967, 0.003469847, 8.542775e-06, -0.0002283165, 
    8.200066e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, -5.181261e-05, 0, 0, 0, 0, 0,
  -2.11705e-05, 0, 0, 0, 0, 0, 0, -2.915672e-05, -4.651621e-05, 
    -4.262479e-05, 0, -1.87429e-07, 0.01573729, 0.009119095, 0.00372278, 
    0.008244063, 0.002935754, 0.001020362, 0.002065616, 0.0276611, 
    0.001904426, 0.04091876, 0.003513187, -1.197321e-06, 0.00417755, 
    -1.989365e-05, 0.005666357, 0.002439415, 0.001263087,
  0, 0, 0, 0, 0, 0, 0.0001609081, -2.267595e-05, 0.0001617404, -0.0001561232, 
    0.0230761, 0.004167772, 0.003000721, -5.256681e-05, -2.447822e-06, 
    -1.358438e-05, 0, 0, 0, -4.982088e-06, 0.006603483, 0.002063659, 
    -3.792061e-05, 0, -6.522172e-08, -0.0002961998, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.002601018, 0.004137632, 0.001523999, 0.00242607, 
    0.0003434146, 0.0003503288, 4.208576e-05, -0.0002370008, -8.740127e-05, 
    0, 0, 0, 0, 0.0005555562, 0, -8.969643e-06, 0, 0, -7.880887e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -5.274376e-08, 0, -0.0002039078, -2.097016e-05, 
    0.01801882, 0.0005361389, -1.568354e-05, -5.251681e-06, 0, 0, 0, 0, 
    -2.789908e-05, 0.000583426, 0, 0, -9.393273e-08, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -1.726657e-05, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0005866437, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.002089471, 0.001695142, 0, 0,
  0, 0, -2.257389e-05, 3.762706e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -8.03917e-07, 0.0007002749, 0, 0, 0, 0, 0, 0, 0, 0, 4.307236e-06, 
    -8.98681e-05, -6.350978e-05, 0.001177977, 0,
  0, 0, 0, 0, 0, 0, -4.060869e-05, 0, 0, 0, 0, 0, 0, 0, 0, -2.90109e-05, 
    2.160598e-05, 0, 0, 0, 0, 0, 0, -9.287453e-08, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0.004847053, 0.000232425, -1.861995e-05, 0, 0, 
    -0.000133966, 0.01514778, 0.0173499, 0.0002787148, -8.508545e-05, 0, 0, 
    0, 0, 0, 0, 0, 0.001498652, 4.984418e-05, 0, 0, 0, 0,
  0, 0.01172126, 0.0007938537, 0, 0, 1.853242e-05, -0.0001217558, 
    0.003366782, -0.0005036614, 0.004181312, 0.008823357, 0.002259003, 
    0.0001125188, 0.0001274211, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0001110065, 0, 
    0, 0, 0, 0,
  -5.510286e-05, 0, 0, 0, 0, 0, 0, 0.0002626573, -0.0002568876, 0.001608647, 
    5.09556e-08, -0.0001081243, 0.03180072, 0.01945211, 0.006678612, 
    0.01673266, 0.008296935, 0.003795568, 0.007750482, 0.04015012, 
    0.006116313, 0.06258518, 0.01041213, 0.000102647, 0.00486993, 
    0.0005644854, 0.009270643, 0.007812337, 0.001135583,
  0, 0, 0, 0, 0, 0, 0.002472179, -0.0001158087, -3.051548e-05, -0.0002698479, 
    0.03736287, 0.01287635, 0.009614972, -5.583945e-05, -4.688327e-06, 
    0.0007322857, 0, 0, 0, -8.653232e-05, 0.01310628, 0.00470697, 
    -7.298674e-05, -2.193821e-05, -6.835789e-07, 0.00258829, 0.0003296851, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.004207053, 0.004615531, 0.01017303, 0.008236018, 
    0.001697425, 0.008540226, -5.818083e-05, -0.0005243531, 0.001718946, 
    -1.147764e-05, 0, 0, 0, 0.001781341, 0.0001073609, 0.0004656807, 
    -4.665671e-06, 0, -0.0001272332, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -1.739246e-05, -4.601426e-05, 0.001364178, 
    0.001440807, 0.0304426, 0.006191449, 0.0007774742, 0.0003747437, 0, 0, 0, 
    0, 0.0004864227, 0.0009613805, -9.0941e-05, 0, 0.0002644317, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001392021, 0, 0.002281927, 
    -3.368898e-06, 7.589472e-06, 0, 0, 0, 0, -2.449964e-05, 0.009535934, 
    1.012176e-06, 0, 0.0002685376, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, -1.152221e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001608351, 0, 
    0, 0.001553583, -7.249587e-06, 0, 0, 0, -6.942182e-06, 0.003790163, 
    0.003426642, 0, 0,
  0, -4.49067e-05, 9.204796e-05, 0.001210957, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0001757115, 0.01177528, 0, 0, -2.579516e-09, 0, 0, 0, 0, 0, 
    0.001187286, 0.008922822, 0.003411999, 0.003782317, 0,
  0, 0, 0, 0, -2.429828e-05, -3.340113e-05, -0.0002738876, 0, 0, 0, 0, 0, 0, 
    0, 3.030915e-06, 0.0008634378, 0.00113931, 0.002697033, 0, 0, 0, 0, 0, 
    -1.857491e-07, 0, -5.668935e-05, 0, 0, 0,
  0, -1.664752e-05, 0, 0, 0, 0, 0.007144061, 0.003456509, 0.003484938, 0, 0, 
    -0.0002850353, 0.01824227, 0.03951813, 0.001770899, 0.0002521914, 0, 0, 
    0, 0, 0, 0, 0, 0.002885957, 0.0001323915, 0, 0, 0, 0,
  0, 0.01626659, 0.002295826, 0, 0, 0.002197282, 0.00513566, 0.01452331, 
    -0.0004922912, 0.01306155, 0.01320583, 0.02170056, 0.0007585455, 
    0.00478151, 0, 0, 0, 0, 0, -1.642343e-09, 0, -2.975207e-06, 
    -2.417258e-05, 0.001537849, -8.312682e-06, 0, 0, -7.407288e-06, 0,
  0.002528193, -1.606619e-05, -7.435376e-07, 0, 0, 3.651586e-08, 0, 
    0.0004662951, -0.0003802091, 0.007154718, 0.0003267124, 0.0009792149, 
    0.05794233, 0.04600804, 0.02239989, 0.03504936, 0.01917174, 0.008277388, 
    0.01006854, 0.06856853, 0.01948326, 0.1265183, 0.01736204, 0.001838697, 
    0.008520728, 0.004742875, 0.01214191, 0.02383994, 0.001453095,
  0, 0, 0, 0, 0, -2.549039e-10, 0.008637235, 0.0002713871, 0.0003484967, 
    -0.0003619637, 0.05206694, 0.02517694, 0.02717919, -5.991453e-05, 
    0.0003851481, 0.001933333, 0, 0, 0, -0.0001351325, 0.02335877, 
    0.01356906, 0.00178869, -7.866944e-05, -2.031376e-06, 0.008704366, 
    0.001630504, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.008830072, 0.006484339, 0.020254, 0.02354565, 
    0.006065949, 0.02086892, 0.007080658, -0.0004819957, 0.007408199, 
    0.0003560103, 0, 0, 0, 0.002985924, 0.004864013, 0.004546701, 
    -5.839358e-05, 0, 0.001392116, 0.0002455346, 0, 0,
  -4.822997e-05, 0, 0, 0, 0, 0, 0, 0, 0, -4.448614e-05, 9.225982e-05, 
    0.008769211, 0.00747145, 0.04573502, 0.01272681, 0.005846427, 
    0.0007885216, 7.994716e-07, 0, 0, 0, 0.001772422, 0.01221018, 
    0.0006959179, 0, 0.02787725, 0.001076214, 0, 0,
  0, -4.782423e-06, 0, -9.610899e-05, 0, 0, 0, 0, 0, 0, 0.001810985, 0, 0, 
    0.005941036, -2.251169e-07, 0.008778214, 0.001061657, 0.0009122181, 0, 0, 
    9.314293e-05, 0.001918684, 0.0003372963, 0.02295977, -7.611265e-06, 
    -7.901977e-05, 0.003912198, -4.593157e-06, 0,
  -0.0001015303, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.400162e-06, 0, 0, 
    0, 0, 0, 0, 0, 0, 7.953724e-05, -0.0002282226, -4.509073e-05, 0, 0, 
    0.0001203066,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, -1.645808e-05, 0, 0.001122706, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, -3.636863e-05, 8.173844e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.004500388, 0, 3.922916e-05, 0.003090102, 0.003175895, 0, 0, 0, 
    7.459193e-06, 0.008187052, 0.008292169, 0.0001791131, 2.16499e-06,
  0, -0.0001092053, 0.0007495228, 0.004400383, 0, -1.890842e-06, 0, 0, 0, 0, 
    0, -5.156893e-08, 0, 0, 0.01784469, 0.03325906, -1.516797e-05, 
    -0.000162745, 0.002114955, 0.004107872, 0.0001364218, -2.028414e-06, 0, 
    0, 0.003533429, 0.02635732, 0.0149418, 0.005605023, 1.717185e-05,
  0, -2.219403e-10, 6.140093e-05, 5.957904e-09, 5.922464e-05, 0.000106764, 
    -0.0001976492, 3.999945e-08, 0, 0, 0, 0, 0, 0, 0.0003122584, 0.00782494, 
    0.00802089, 0.006347543, 0, 0, 0, 0, 0, -2.087652e-06, 0.0002972858, 
    0.00022418, -1.026717e-06, 0, 0,
  0, -1.234402e-05, 5.063643e-05, -6.573477e-07, 0, 0, 0.01149735, 
    0.008857847, 0.007154816, 0, -1.322011e-05, -8.000488e-05, 0.0229218, 
    0.07670309, 0.01606822, 0.001065353, 0, 0, 0, 0, 0, 0, 0, 0.009331354, 
    0.0005409045, 0, 0, 0, 0,
  9.24996e-07, 0.02999467, 0.006673079, 0, 0, 0.004305054, 0.02861732, 
    0.04357098, 0.00575551, 0.02569504, 0.02076055, 0.05510927, 0.01416962, 
    0.0140539, 2.580284e-06, 0.0004511682, 0, 0, 0, -1.246931e-06, 
    1.807331e-09, 0.001005872, 0.002044175, 0.01002378, -2.696222e-05, 
    -1.594953e-05, 0, -2.280094e-05, -1.007776e-06,
  0.01565019, 0.0003306642, -1.789237e-06, 9.318296e-06, 0, 8.007867e-05, 
    0.0006061658, 0.01253241, 0.006556711, 0.02688361, 0.0004990405, 
    0.01373344, 0.1021275, 0.08322516, 0.04860292, 0.05747265, 0.02984068, 
    0.01205728, 0.01464196, 0.1044602, 0.04441098, 0.2083733, 0.04158721, 
    0.006842055, 0.01980191, 0.01507122, 0.02841404, 0.0365794, 0.008075035,
  0, 0, 0, 0, 2.119019e-07, 4.696594e-05, 0.02369689, 0.004404914, 
    0.01127735, 0.003154384, 0.06879716, 0.03582728, 0.05808266, 
    -0.000281789, 0.004033742, 0.002913108, 0.001802831, -3.737134e-08, 0, 
    -1.08896e-05, 0.04487002, 0.04512285, 0.004551253, 0.0006958916, 
    -1.424118e-05, 0.02086826, 0.003206865, 0, 0,
  0, 0, 0, 0, 0, 0, -2.820191e-08, 0.01992368, 0.009993506, 0.02356676, 
    0.04654703, 0.008162831, 0.03852918, 0.02276097, -0.0006846486, 
    0.01654015, 0.001450551, -9.193462e-08, 0, 0, 0.006739598, 0.01351436, 
    0.02791243, 0.001026908, 0.0001919183, 0.01064364, 0.003482279, 0, 
    -5.759725e-06,
  6.25463e-06, 0, -3.477086e-05, 0, 0, 0, 0, 0, 4.760515e-05, -3.646068e-05, 
    0.00280827, 0.02556172, 0.02383007, 0.06182907, 0.02189273, 0.01711096, 
    0.007151959, -1.986671e-05, 0, 0, 0, 0.00303717, 0.01765425, 0.003681912, 
    1.942869e-05, 0.06183925, 0.001973885, 0, -6.562739e-06,
  0, 0.001180165, 0, 0.001118722, -1.661874e-07, -7.108452e-05, 0, 0, 0, 
    -3.433193e-05, 0.007363665, 0, -1.788485e-05, 0.01449528, 0.0002431129, 
    0.01556275, 0.003856189, 0.005797517, -1.682073e-10, 0, 0.0008563458, 
    0.002984956, 0.002759357, 0.03965739, 0.005311573, 0.002078095, 
    0.008562854, 0.002719369, -2.626796e-05,
  9.524312e-05, -1.16431e-06, 0, -1.903805e-05, 0.004227682, 0, 0, 0, 0, 0, 
    0, 0, 0, 6.527681e-05, 0.006246218, -2.77653e-05, 0.001442337, 0, 
    0.0009739827, -8.616473e-11, -1.235578e-09, -1.976801e-10, 0, 
    0.004129256, 0.003189943, 0.001334809, -5.038086e-05, 0, 0.001404512,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.001939088, -7.600936e-06, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -4.131926e-09, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0.0008725772, 0, -4.14609e-05, -0.0001452975, 0.001786552, 0.002965569, 
    0, 0, 0, 0, 0, 0, -3.626838e-06, -6.960699e-06, 0, 0, 0, 0, 
    -1.320232e-05, 0, 0.0005951063, 2.366842e-07, 0, 0, 0, 0, 0, 0,
  0, -0.000212244, 4.024229e-06, 0.0001568153, 0.001331761, 1.188808e-05, 
    0.0001213705, 0, 0, 0, 0, 0.001790054, 0.0007359316, 3.074282e-05, 0, 0, 
    0.006724316, 0, 0.001983273, 0.01216576, 0.01365948, 0.0005022628, 
    0.0003626853, 0, 0.003954867, 0.01188501, 0.01430278, 0.005103887, 
    0.006693348,
  6.861805e-05, 0.001121369, 0.001427845, 0.008932107, 0, 3.24242e-05, 0, 
    5.240645e-09, 5.423284e-08, -3.844954e-08, -2.591106e-10, 0.0004783301, 
    0, 0, 0.03565358, 0.06514537, 0.003072449, 0.006421079, 0.02479143, 
    0.00508352, 0.0007201855, 0.002531176, 3.176756e-05, 6.936576e-09, 
    0.009297855, 0.04559592, 0.0283432, 0.007297894, 3.386635e-05,
  0, 1.259794e-05, 0.009491317, 5.477596e-07, 0.001377094, 0.004039528, 
    0.0006993245, 0.0003272257, 5.666486e-08, 1.422198e-06, 0, 2.24681e-08, 
    2.058252e-08, -2.446131e-07, 0.004964566, 0.03313636, 0.03664198, 
    0.02255308, 0.003315928, -1.491992e-08, 0, -1.344332e-09, 0, 
    0.0003198152, 0.00111272, 0.004465561, 0.0001201964, 2.789568e-07, 
    -4.224208e-07,
  -6.948535e-11, -1.400548e-05, 0.0002913961, 0.0002015571, -9.177233e-11, 
    -7.603288e-10, 0.02140651, 0.04195994, 0.007698529, -2.988989e-05, 
    -7.254703e-05, 0.001355903, 0.05482536, 0.1896626, 0.1468805, 
    0.004441677, -1.798079e-05, -1.472763e-06, -1.078093e-09, 1.322053e-05, 
    3.809613e-06, 7.743822e-05, 4.427724e-07, 0.02895688, 0.02241882, 
    7.408274e-05, 0, -4.767138e-10, 0,
  3.667933e-05, 0.07376056, 0.02461835, 0.0002490722, -8.664547e-12, 
    0.01717106, 0.051157, 0.1169906, 0.04854549, 0.07369952, 0.07992545, 
    0.1681496, 0.0785025, 0.03838981, 0.0002025713, 5.287905e-05, 
    -1.177236e-05, 0, 9.523569e-09, 5.580832e-05, 0.000488901, 0.002870806, 
    0.01673841, 0.07773181, 0.003319387, 5.783884e-05, -4.757804e-10, 
    0.0002391186, -3.29449e-05,
  0.06120208, 0.004112876, 0.0005556771, 0.0002867908, -3.043333e-07, 
    0.0001530545, 0.03441484, 0.2047147, 0.4034996, 0.3638491, 0.2316609, 
    0.2935253, 0.2650338, 0.1994767, 0.1429655, 0.1112511, 0.04735129, 
    0.01536672, 0.01753738, 0.1352882, 0.2332805, 0.4063745, 0.07595796, 
    0.03163847, 0.05437447, 0.02571106, 0.06655107, 0.07306163, 0.01901295,
  -2.597019e-07, 8.95365e-06, 0, 1.890842e-07, 0.0001102008, 0.02148897, 
    0.2503071, 0.1218783, 0.1704847, 0.05381058, 0.1275051, 0.1356729, 
    0.1655368, 0.006355453, 0.008756956, 0.009060838, 0.007239896, 
    0.002199758, 3.522541e-07, 0.01909485, 0.1601001, 0.1563239, 0.03279355, 
    0.02734538, 0.0001125714, 0.03412525, 0.01253659, 0.004130303, 
    1.725069e-06,
  -8.437714e-06, 0, 0, -4.042883e-10, 0, 0, -1.777245e-05, 0.02474244, 
    0.01417759, 0.04302162, 0.08961098, 0.03951184, 0.1332528, 0.1597951, 
    0.04006131, 0.03929574, 0.02471266, -3.180613e-05, 0, -1.098634e-08, 
    0.01796971, 0.09365842, 0.09550796, 0.003957429, 0.0005480588, 
    0.04063243, 0.008083553, 2.064142e-05, 0.0005168817,
  0.000944986, -6.343469e-05, 0.0008064572, 0, -1.97496e-06, 1.793157e-05, 
    -1.371607e-08, 2.922997e-06, 0.0006988527, 0.004704025, 0.02492471, 
    0.03980597, 0.06335934, 0.1208128, 0.06930175, 0.05159536, 0.01934103, 
    0.001001332, 0.0005099092, 0, 0, 0.004997242, 0.02865376, 0.00946553, 
    0.001585955, 0.07772677, 0.004928365, -1.018674e-05, 2.235213e-05,
  0, 0.006705887, 0.001867335, 0.004596033, -8.705648e-05, -2.778389e-05, 0, 
    0, 0, -3.923649e-05, 0.01622304, -3.273751e-05, 0.0008968209, 0.02271388, 
    0.01310803, 0.02139471, 0.01325783, 0.01302374, 0.0002257118, 0, 
    0.003400742, 0.00882555, 0.0091228, 0.05234106, 0.009128892, 0.01144398, 
    0.02425977, 0.01498562, -0.0001919065,
  0.005794088, 2.690049e-05, -2.518372e-05, -6.713808e-05, 0.009117389, 
    -0.0001339194, 0, 0, 0, 0, -1.606106e-05, 0, 0, 0.004504856, 0.01405375, 
    0.003793717, 0.005592282, -3.603274e-05, 0.004922381, -1.16897e-05, 
    -4.28025e-10, -2.225126e-05, 0, 0.004155871, 0.01723991, 0.01032044, 
    0.0008233587, 0, 0.006982683,
  0, 4.727401e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, -1.799819e-05, 0.006617347, -3.303066e-05, 0, 0.0003558002, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, -2.573234e-06, 0, 0, -2.151633e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, -7.461312e-06, 0, 0, 0, 0.002799994, 0, 0, 0, 0,
  0.001516851, 0.004352494, 0, -0.0002993616, 0.002967157, 0.005526523, 
    0.004698166, 2.774344e-07, 0, 0, 0, 0, 0, 0.001487641, 0.0003544267, 
    5.351043e-05, 0, 0, 0, 0.0005498354, 3.689437e-05, 0.004745112, 
    0.008244332, 0.0006555502, 0.0001085562, 0, -8.919832e-07, 0.0002140747, 
    -8.165475e-06,
  -0.0001108237, 0.002629978, 0.003867642, 0.001444055, 0.01066049, 
    0.0006621666, 0.004919372, 0, 7.521744e-08, -2.14542e-08, -5.556248e-07, 
    0.005817895, 0.00909102, 0.00436041, 0, 0.00110009, 0.00761067, 
    0.001989955, 0.003765395, 0.02772425, 0.02588185, 0.007631854, 
    0.004827545, 0.002641332, 0.00788359, 0.01871058, 0.0190054, 0.01462748, 
    0.0219411,
  0.0005037358, 0.003060085, 0.003966005, 0.01879293, 0.0003680136, 
    0.001667849, 5.668726e-08, 6.836003e-07, 0.0004948188, -2.560048e-05, 
    -5.691941e-07, 0.001553824, -6.577417e-06, -6.269126e-09, 0.0581596, 
    0.1023748, 0.03461718, 0.02796299, 0.07235663, 0.033424, 0.01070495, 
    0.01554056, 0.006467844, 0.001506212, 0.01537538, 0.1039585, 0.07231573, 
    0.01473311, 0.0009472028,
  3.018038e-06, 0.0002848801, 0.01828721, 0.0002029233, 0.01235094, 
    0.01586931, 0.007140816, 0.003496831, 1.060559e-05, 1.318923e-06, 
    4.614402e-08, 7.965366e-08, 2.782487e-08, 5.150676e-06, 0.02509387, 
    0.07646876, 0.08317091, 0.07595623, 0.01753025, -1.142565e-06, 
    6.18541e-07, 9.965642e-07, 3.620348e-06, 0.04044962, 0.192697, 
    0.03115632, 0.003694218, 0.0002163793, 0.002779223,
  3.088446e-06, -0.0007773667, 0.02648923, 0.007912273, 8.784863e-06, 
    8.880498e-05, 0.06088402, 0.1120246, 0.02469148, 0.0001879568, 
    0.0001100274, 0.001805775, 0.05329019, 0.2028545, 0.2161961, 0.1100575, 
    0.00781438, 1.776527e-06, 3.107739e-06, 0.0001266232, 4.469495e-06, 
    0.0001537981, 0.0002332277, 0.2194352, 0.2806474, 0.004103807, 
    1.358654e-06, 7.098067e-05, 3.112022e-05,
  0.05524296, 0.4119256, 0.4181103, 0.01171475, 3.214119e-05, 0.1221077, 
    0.233553, 0.323259, 0.2470497, 0.2773297, 0.1077651, 0.1672759, 
    0.08907752, 0.05293262, 0.0006845074, 0.002934414, -4.0031e-05, 
    3.357316e-05, 2.250856e-05, 0.03550509, 0.002142199, 0.03031215, 
    0.06839759, 0.2556576, 0.03865566, 0.002880629, 0.002361359, 0.04543114, 
    0.01989713,
  0.2506035, 0.1474837, 0.1387942, 0.000827016, 0.001433314, 0.008985242, 
    0.1114293, 0.1839605, 0.3441515, 0.2733256, 0.1484648, 0.2434001, 
    0.2573469, 0.1964385, 0.1824077, 0.1854059, 0.1081718, 0.0239576, 
    0.02178068, 0.2028924, 0.3055274, 0.4886021, 0.227974, 0.1616402, 
    0.08942987, 0.06954668, 0.1785304, 0.1791894, 0.1535803,
  0.002340928, 0.02951826, 0.009336075, -1.506047e-06, 0.003275607, 
    0.02282115, 0.2398242, 0.07531302, 0.1572133, 0.02782194, 0.1007622, 
    0.09065462, 0.1441615, 0.03038027, 0.02919567, 0.08797454, 0.08867346, 
    0.01748299, 1.358256e-07, 0.008114488, 0.1189549, 0.1731002, 0.04533328, 
    0.1166483, 0.06759728, 0.06353896, 0.08448116, 0.1128432, 0.05222454,
  0.001005785, -9.048429e-06, 0.0002145113, 0.001060201, 0, -1.136218e-08, 
    -9.440725e-06, 0.03018828, 0.02383978, 0.03878098, 0.07968818, 
    0.04203045, 0.1322459, 0.1812701, 0.06932286, 0.09737822, 0.07611437, 
    0.08316307, 0.0001101356, 1.006391e-05, 0.06004957, 0.1950061, 0.2549603, 
    0.1084163, 0.1072067, 0.1451869, 0.06973325, 0.02675426, 0.004555951,
  0.002268728, 0.001917659, 0.002221572, -2.451574e-06, 0.0007678627, 
    0.002033351, 8.826527e-08, 0.001288663, 0.005056971, 0.04573964, 
    0.05595292, 0.1037907, 0.1552496, 0.2608246, 0.1904829, 0.2236381, 
    0.04453805, 0.02549488, 0.0310028, 0.0004117432, 4.082523e-05, 
    0.007194079, 0.08488762, 0.04150203, 0.06323986, 0.129586, 0.04731572, 
    0.00423272, 0.01174678,
  0.0001554619, 0.02019355, 0.004218793, 0.00776908, 0.003845002, 
    0.0003548753, -2.165753e-06, -2.026814e-05, 0.0003350409, 0.0001048021, 
    0.02933811, 0.0005214853, 0.01506832, 0.07116394, 0.03817683, 0.04002263, 
    0.05685769, 0.03372463, 0.0206465, 0.0004364441, 0.007742003, 0.01709761, 
    0.01879378, 0.06379676, 0.01920426, 0.03077625, 0.0815184, 0.03961893, 
    0.001697905,
  0.0232137, 0.00310649, -9.048192e-05, 0.0003447301, 0.01132944, 
    -0.0001758144, -2.695383e-09, 0, 0, -2.078065e-05, 0.0009065717, 
    -1.972395e-06, -0.0001046695, 0.008663917, 0.02635412, 0.02945479, 
    0.01454432, 0.0001153231, 0.009431949, 0.0005327932, 0.0009570807, 
    0.0008902011, 0, 0.004904736, 0.04493847, 0.03632667, 0.01326731, 0, 
    0.01801126,
  -4.815727e-05, 0.003137488, 0.0001402465, 0.001622775, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.000540616, -2.309643e-05, 0, 0, 0, 0, -3.135176e-05, 
    0.01310894, 9.541075e-05, 1.549736e-05, 0.005446964, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -2.259028e-05, -6.909158e-08, 0, 0, -1.386659e-13, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0.0006760372, -1.406661e-05, 0, -2.231673e-06, 0, 0, 
    -7.83875e-06, -0.000103569, -5.888257e-05, 0.0009279374, -4.392544e-05, 
    -1.367401e-07, 0, 0, 0, 0, -4.537053e-05, 0, 2.090976e-05, 0, 
    0.004065834, -6.923798e-05, 0, 0, 0,
  0.008095167, 0.01410246, -8.466774e-06, 0.00351022, 0.008867174, 
    0.01532354, 0.009535013, 0.001573358, -0.0002450033, 0.001536158, 
    0.001866044, 0.0001821578, 2.969793e-07, 0.00925338, 0.00750484, 
    0.002691243, -5.890622e-06, 0.0005279623, 0, 0.002532994, 0.008527495, 
    0.01523479, 0.01694154, 0.006882973, 0.005101373, 0.0003516398, 
    -3.42703e-05, 0.004985381, 0.006036427,
  0.0511441, 0.04797908, 0.01681557, 0.007841481, 0.0320981, 0.02915773, 
    0.01155213, -1.985951e-05, 4.996885e-06, -2.826501e-05, 0.0001972329, 
    0.01044727, 0.01527125, 0.01360837, -1.54832e-06, 0.003891843, 0.014513, 
    0.009514243, 0.01370967, 0.03578391, 0.07312292, 0.05353241, 0.01875901, 
    0.01108672, 0.01444067, 0.02968891, 0.04028958, 0.04529391, 0.0654792,
  0.03765809, 0.0393702, 0.01024576, 0.09156011, 0.03694425, 0.01227851, 
    0.004457145, -4.57711e-05, 0.02199979, 0.008143228, 0.01065098, 
    0.01816769, 0.01310563, 0.002703771, 0.06847878, 0.150545, 0.1024272, 
    0.06553151, 0.1462909, 0.1222125, 0.03406705, 0.02462947, 0.02568989, 
    0.02000892, 0.03149622, 0.1312593, 0.1134125, 0.09327576, 0.04429642,
  4.445328e-07, 0.005009303, 0.1086546, 0.0219672, 0.02672327, 0.01562443, 
    0.003230011, 0.005235771, 9.29569e-06, 3.115699e-07, 3.400879e-08, 
    2.813926e-08, 2.667036e-08, 5.994156e-06, 0.02897456, 0.1093318, 
    0.09373511, 0.1071841, 0.01042227, -2.307032e-06, 1.226872e-08, 
    3.291135e-08, 7.615989e-07, 0.0445294, 0.1487185, 0.1349585, 
    0.0002160033, 0.003005887, 0.0003070929,
  1.512032e-06, -0.0001514456, 0.02153767, 0.001101178, 2.025195e-06, 
    0.001856818, 0.02915131, 0.1109929, 0.02262726, 1.74818e-05, 
    -8.363016e-05, 0.0006082169, 0.03589872, 0.1621145, 0.1522689, 0.0813022, 
    0.006439243, 6.50471e-06, 5.275059e-08, 3.943406e-06, 1.212998e-06, 
    8.886653e-06, 4.293079e-06, 0.1788172, 0.1929151, 8.063993e-05, 
    6.059257e-07, 5.440103e-06, 6.805275e-07,
  0.01176618, 0.3837976, 0.2993493, 0.003758618, 1.359173e-05, 0.08855357, 
    0.1679118, 0.2400402, 0.2013611, 0.203916, 0.08215262, 0.145291, 
    0.05802292, 0.03578116, 0.0002733489, 0.0005950994, 3.76775e-05, 
    5.858189e-06, 5.269143e-06, 0.0108775, 9.955074e-05, 0.01214551, 
    0.06352522, 0.209311, 0.01768245, 0.002418811, 0.0001748968, 0.009306278, 
    0.00746269,
  0.2081532, 0.1053512, 0.08488443, 0.01364748, 0.000972521, 0.004970196, 
    0.06725123, 0.1367053, 0.2592035, 0.1786285, 0.09463122, 0.1669492, 
    0.2027886, 0.1786443, 0.1610793, 0.1504581, 0.08557725, 0.01819434, 
    0.0210616, 0.1675832, 0.2168733, 0.459901, 0.1991591, 0.1085311, 
    0.06793054, 0.04015009, 0.1225199, 0.1591816, 0.09876635,
  0.0001749396, 0.02131538, 0.004815829, 0.0001056764, 0.009475616, 
    0.02641437, 0.2085915, 0.0676985, 0.1011377, 0.02495675, 0.09650671, 
    0.0779902, 0.1321262, 0.02042166, 0.01344934, 0.08271603, 0.07989287, 
    0.01028205, 7.368919e-08, 0.01196332, 0.09086637, 0.1362096, 0.02460932, 
    0.08623383, 0.03074135, 0.04948786, 0.068914, 0.1435903, 0.1064415,
  0.1054997, 0.01336474, 0.0001282635, 0.0002645694, 0, 3.229787e-08, 
    -2.874149e-06, 0.03455052, 0.05520908, 0.04511972, 0.06875115, 
    0.03651101, 0.1129562, 0.13932, 0.04041663, 0.08357025, 0.05837723, 
    0.09815658, 0.02220064, 4.551508e-06, 0.06487954, 0.1327369, 0.2103174, 
    0.06963506, 0.09075251, 0.0972169, 0.06384979, 0.06613215, 0.07897185,
  0.09541996, 0.04105048, 0.01023368, 0.0003363571, 0.00321715, 0.02741656, 
    0.001408177, 0.01293617, 0.04506965, 0.08704944, 0.1235256, 0.1167842, 
    0.2127628, 0.238166, 0.1869988, 0.2519127, 0.1023412, 0.1347531, 
    0.09008171, 0.002537037, 0.002717554, 0.05035877, 0.1113373, 0.08531531, 
    0.1140797, 0.1733025, 0.1084874, 0.06567217, 0.08065993,
  0.04675009, 0.03052681, 0.01153565, 0.02565642, 0.03396456, 0.003321737, 
    0.003523734, -5.362518e-05, 0.001937406, 0.001985924, 0.03673492, 
    0.01762774, 0.04114875, 0.1177205, 0.06155989, 0.08540149, 0.08631223, 
    0.1055145, 0.1077795, 0.02929583, 0.02869909, 0.06952247, 0.03549423, 
    0.08520401, 0.0581023, 0.0792171, 0.1522696, 0.08121514, 0.06718268,
  0.0497926, 0.01960189, 0.0005366886, 0.005022397, 0.01333683, 0.00053613, 
    1.763354e-05, 0.0001828423, 0, 0.001363896, 0.005494862, -1.151751e-05, 
    0.001507093, 0.07814681, 0.03792935, 0.02059361, 0.02722298, 0.01707907, 
    0.01939933, 0.01494808, 0.01710093, 0.0170747, -3.45821e-05, 0.008789666, 
    0.06559082, 0.0467455, 0.06885913, 0.00777012, 0.03803707,
  0.003487279, 0.01308819, 0.0004337469, 0.004754583, 0, 0, 0, 0, 0, 
    -7.636868e-06, 5.941738e-05, -3.987258e-05, 0, 0, 0.0001071152, 0, 
    -1.572608e-05, 0.004999769, -7.251883e-05, -3.079828e-05, -2.97968e-05, 
    0.0003122264, 0, 1.047599e-05, 0.02782755, 0.0008505926, 0.002856897, 
    0.02678283, 0.01850714,
  0, 0, -1.093182e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -5.487416e-05, 
    -8.764776e-05, 0, 2.640497e-05, 0, 3.463278e-06, 0.0001525665, 
    -3.090734e-07, -3.684231e-05, -0.0002295225, 2.000067e-05, -3.16794e-10, 
    -5.033446e-05, 2.909437e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, -1.823854e-05, -8.122645e-06, 0, 0.002084943, 9.884e-05, -1.321309e-05, 
    -3.665641e-05, -3.058281e-06, 0, -2.438529e-05, -0.00030626, 0.001352062, 
    0.002290255, 0.0006261951, 0.0003032894, -4.391996e-05, 0, 0, 0, 
    0.004458278, 0.00109383, 0.002087728, -2.704699e-06, 0.004895203, 
    0.002981239, -1.257377e-05, 0.001051027, 0,
  0.02440376, 0.04864612, 0.01814774, 0.02478013, 0.03209614, 0.04170712, 
    0.03449965, 0.009849236, 0.005385921, 0.007432404, 0.005456863, 
    0.001613634, 0.003393383, 0.02701678, 0.01521476, 0.01002595, 
    0.001610251, 0.002812167, 0.002029881, 0.008629377, 0.03103009, 
    0.0364529, 0.05353537, 0.03605397, 0.0516515, 0.01198772, 0.001938066, 
    0.007281002, 0.0315104,
  0.1085362, 0.07570712, 0.1068816, 0.1273087, 0.2507493, 0.1323018, 
    0.07844432, 0.03968281, 0.03800214, 0.02141517, 0.00552981, 0.02220904, 
    0.04514246, 0.03755858, 0.0062762, 0.0371615, 0.05595215, 0.03430239, 
    0.02492182, 0.06751344, 0.1607927, 0.1394068, 0.1161914, 0.03219094, 
    0.09940507, 0.08026201, 0.08943938, 0.07851315, 0.121333,
  0.03862131, 0.03109048, 0.07712628, 0.1410146, 0.04490277, 0.01559359, 
    0.0002596584, -0.0002425815, 0.02304758, 0.009800116, 0.01167069, 
    0.0173289, 0.01257903, 0.003288442, 0.07112048, 0.151805, 0.09163914, 
    0.10442, 0.2355822, 0.1337857, 0.03026463, 0.04450259, 0.0576843, 
    0.04503924, 0.0564871, 0.1318708, 0.132753, 0.1091542, 0.04843682,
  1.020204e-07, 0.008270652, 0.1433169, 0.0153062, 0.02930614, 0.01550179, 
    0.0003748066, 0.01621956, 3.080768e-06, 1.253238e-07, 9.440301e-09, 
    1.007401e-08, 1.86407e-07, 1.056069e-05, 0.03207092, 0.1114887, 
    0.09812088, 0.07828172, 0.004865051, -5.609644e-08, -3.106448e-11, 
    -2.898968e-10, 1.261036e-08, 0.05059927, 0.130016, 0.1211216, 
    -0.0005247686, 0.001078595, 5.064786e-06,
  4.560754e-07, -7.925805e-05, 0.01331225, 0.002212505, 7.18624e-08, 
    0.001054263, 0.02194881, 0.1120353, 0.02279986, 2.307004e-06, 
    1.293028e-05, 0.004075414, 0.03643244, 0.1455996, 0.1277342, 0.06696831, 
    0.003319334, 6.359975e-06, 3.18175e-07, 5.491476e-07, 3.984205e-07, 
    1.081295e-06, 5.126631e-07, 0.1561899, 0.1633054, 3.789522e-06, 
    2.733572e-07, 1.96713e-06, 4.288227e-07,
  0.002881865, 0.3563524, 0.2124247, 0.0001420927, 0.0001978828, 0.06344829, 
    0.143371, 0.2013069, 0.1800423, 0.1558266, 0.07118133, 0.1326777, 
    0.04706947, 0.03825225, 0.001086812, 5.20657e-05, 6.849263e-05, 
    7.634455e-06, 1.767315e-06, 0.0006737362, 1.436582e-05, 0.004671913, 
    0.04760744, 0.1855562, 0.01177109, 0.00238285, 0.0001533206, 0.001357774, 
    0.0001377846,
  0.1877892, 0.09050556, 0.05758924, 0.004693497, 0.0003065472, 0.003531163, 
    0.05258452, 0.1066432, 0.203104, 0.1304583, 0.06423011, 0.1180802, 
    0.1842051, 0.1663523, 0.1554722, 0.1323374, 0.07903784, 0.02064532, 
    0.02283673, 0.144991, 0.1632323, 0.402434, 0.1813196, 0.08531347, 
    0.06631269, 0.03297708, 0.09611846, 0.1496306, 0.1021892,
  -5.30852e-05, 0.01049333, 0.0004960105, 1.374719e-05, 0.0007381261, 
    0.02504393, 0.1798612, 0.06265116, 0.07907263, 0.02413767, 0.08565108, 
    0.0686733, 0.1333335, 0.02537661, 0.01103993, 0.0667805, 0.07777179, 
    0.0003602726, 2.007876e-07, 0.006091348, 0.07576441, 0.1247781, 
    0.02758421, 0.07697598, 0.02538219, 0.05047559, 0.06188559, 0.1273778, 
    0.09280258,
  0.1033506, 0.006902059, 2.231815e-05, 2.907117e-05, 0, 9.670453e-08, 
    -2.441688e-06, 0.07478124, 0.1290484, 0.07284132, 0.05753041, 0.03238244, 
    0.09255876, 0.1192206, 0.02750783, 0.06858011, 0.03959882, 0.06757901, 
    0.01130424, -5.37081e-06, 0.04541853, 0.107237, 0.1946929, 0.07120943, 
    0.08123054, 0.06892083, 0.06346597, 0.04458411, 0.0912048,
  0.1456517, 0.08249489, 0.01579791, 0.006929414, 0.00141685, 0.03321862, 
    0.002821858, 0.1104571, 0.1625394, 0.1711514, 0.1744443, 0.1362421, 
    0.2099689, 0.2142337, 0.1751992, 0.2398158, 0.09292804, 0.1368756, 
    0.0958335, 0.04798137, 0.08250258, 0.03213521, 0.09367377, 0.08664735, 
    0.08666512, 0.1567473, 0.10607, 0.05954389, 0.1041548,
  0.1043796, 0.124247, 0.1302732, 0.1673457, 0.1467091, 0.1185109, 
    0.03588349, 0.0005790966, 0.002181114, 0.004474551, 0.04608793, 
    0.06574022, 0.07779585, 0.1549737, 0.1107763, 0.1254212, 0.1254054, 
    0.1274628, 0.1354172, 0.04041234, 0.05738412, 0.1066915, 0.08052406, 
    0.1141304, 0.06675909, 0.09782826, 0.1772986, 0.1309998, 0.1396165,
  0.1511977, 0.0946178, 0.04696681, 0.06998219, 0.05633078, 0.01731238, 
    0.00576119, 0.001357312, 0.0008159872, 0.01489333, 0.01886649, 
    0.02285237, 0.07429506, 0.1001823, 0.03343314, 0.05990521, 0.04790016, 
    0.08590323, 0.05900973, 0.08099633, 0.06867778, 0.06594221, 0.007060942, 
    0.03450438, 0.128945, 0.1352923, 0.1902401, 0.06267066, 0.1335895,
  0.01556308, 0.0315574, 0.02166433, 0.06447604, 0.01940604, 0.01180574, 
    8.657054e-05, -5.699361e-09, 0, 0.001346667, 0.004453682, -0.0003943056, 
    0.03609462, 0.04321975, 0.04522654, 0.03767489, 0.005274408, 0.02511259, 
    0.05242082, 0.06104558, 0.03649922, 0.02649854, 0.03608171, 0.002395891, 
    0.04447173, 0.005783226, 0.01021654, 0.04069238, 0.02277388,
  -0.0001842443, 0.0001230506, -0.0003786436, 0.0003086943, 0.0006933554, 
    0.0008649475, 4.420407e-05, 0, 0, 0, 0, 0, 0, -2.855088e-05, 
    -3.052782e-05, 0.0001061215, -0.0001631266, 0.01055114, 0.02363876, 
    0.01591658, 0.001668052, 0.0003372089, -3.304083e-05, 0.0002875909, 
    0.003648616, 0.0003401537, -0.00074115, 0.006095942, 0.002042236,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0.0001105272, -7.859999e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.006483078, 0.006293155, 0.0006354065, 0, 0, 0, 7.919124e-05, 0, 
    4.989892e-05, 0, 0, 0, 0, 0, 0,
  -4.622279e-05, -7.228284e-05, 2.603357e-05, -1.379298e-05, 0.008077858, 
    0.005972483, 0.01074582, 0.001880518, 0.0032673, 0.001196043, 
    -2.827507e-05, 0.005846807, 0.00351451, 0.006202494, 0.01088355, 
    0.0184492, 0.01531432, 0.00215148, -3.913255e-05, 0.0001065741, 
    0.007779766, 0.00576836, 0.01491296, 0.01024666, 0.02906579, 0.01608448, 
    0.002960399, 0.003804196, 0,
  0.1053776, 0.1112528, 0.09975202, 0.09411145, 0.1076647, 0.1217017, 
    0.1105944, 0.09408183, 0.08275691, 0.05525736, 0.07625221, 0.07582219, 
    0.07516826, 0.1344488, 0.1106335, 0.06508956, 0.04551339, 0.03474614, 
    0.02864088, 0.0449737, 0.0677715, 0.06075433, 0.10399, 0.07218536, 
    0.09619068, 0.06531332, 0.03763326, 0.08078732, 0.09863149,
  0.1693758, 0.1216015, 0.1246596, 0.1591823, 0.2424479, 0.1369519, 
    0.1109417, 0.08069701, 0.0678717, 0.04481117, 0.03623587, 0.07597993, 
    0.06621248, 0.1064363, 0.02243724, 0.06139519, 0.1229482, 0.1068912, 
    0.07746746, 0.097233, 0.1825403, 0.172915, 0.1547351, 0.06437846, 
    0.1831184, 0.127602, 0.1667486, 0.1372261, 0.1900963,
  0.04550297, 0.0148644, 0.07295588, 0.113708, 0.05558793, 0.02742831, 
    0.001067306, -9.074021e-05, 0.002091904, 0.001142434, 0.003924657, 
    0.01573072, 0.0126952, 5.426518e-05, 0.07411072, 0.1518831, 0.07994673, 
    0.1057351, 0.2179881, 0.1232961, 0.02793546, 0.04094868, 0.05899522, 
    0.04253124, 0.06130048, 0.1269908, 0.1239137, 0.07862977, 0.03350809,
  7.066146e-08, 0.01068918, 0.1226499, 0.009438972, 0.02558749, 0.01468745, 
    -0.0002898346, 0.02498806, 7.860872e-06, -8.884041e-07, -3.453501e-07, 
    -5.953487e-08, 8.510866e-08, 0.0003824556, 0.0526586, 0.09650861, 
    0.1049982, 0.05213965, 0.003209234, -1.011112e-07, 0, 3.342052e-11, 0, 
    0.06591415, 0.1128807, 0.1105328, -7.170262e-06, 0.007127867, 2.82825e-06,
  5.182416e-08, -5.183064e-05, 0.01151471, 0.001114203, 1.43661e-06, 
    0.0006508522, 0.02010396, 0.1117684, 0.02605165, 3.718119e-06, 
    0.0001725213, 0.007659399, 0.03960843, 0.1311023, 0.08990246, 0.04449346, 
    0.001799385, -1.202867e-06, 4.123567e-07, 1.733386e-07, 2.92629e-07, 
    1.086599e-06, 2.889203e-07, 0.1108009, 0.1298, 1.963696e-06, 
    3.166749e-07, 2.058692e-07, 7.967692e-07,
  0.0004810807, 0.2955885, 0.1354043, 1.34301e-05, 0.0007023176, 0.04105646, 
    0.111479, 0.1578618, 0.1546557, 0.1322675, 0.06081866, 0.119464, 
    0.03213424, 0.0355728, 0.004139919, 2.026149e-05, 3.299776e-05, 
    1.406978e-06, 3.10079e-06, 2.412794e-05, 1.440251e-05, 0.006086804, 
    0.04216709, 0.1519625, 0.007469545, 1.203751e-05, 5.583148e-05, 
    0.0001433971, 2.42679e-06,
  0.1435588, 0.07523711, 0.05429818, 0.002105371, 8.410337e-05, 0.006369498, 
    0.03265022, 0.07821752, 0.1478471, 0.09629983, 0.04699646, 0.07151405, 
    0.159557, 0.1515878, 0.1357685, 0.1310082, 0.06753894, 0.02457429, 
    0.02851092, 0.1504648, 0.1146154, 0.3591691, 0.1582597, 0.06405784, 
    0.06021676, 0.02871669, 0.07679202, 0.1292591, 0.09802929,
  -1.285729e-05, 0.0009800012, 2.431663e-05, 2.884755e-06, 3.405795e-06, 
    0.01523455, 0.1611055, 0.04930502, 0.0685633, 0.01720512, 0.08114104, 
    0.05332422, 0.12718, 0.02321454, 0.008981361, 0.05418814, 0.05722122, 
    7.185098e-07, 2.947695e-08, 0.0238967, 0.06499144, 0.1186525, 0.02608761, 
    0.05539601, 0.01861521, 0.05021143, 0.05773773, 0.1118341, 0.040309,
  0.07716397, 0.002264047, 1.194743e-05, 1.484683e-06, -7.57696e-08, 
    1.441662e-08, -1.472829e-05, 0.07432902, 0.1347931, 0.08640233, 
    0.04890678, 0.02428826, 0.0855452, 0.1093441, 0.02092884, 0.06640363, 
    0.02905276, 0.03530543, 0.007047384, -3.079584e-05, 0.0320963, 
    0.09347054, 0.165975, 0.06059695, 0.06607185, 0.04850812, 0.05351965, 
    0.02854211, 0.08527528,
  0.1283202, 0.07703674, 0.01415339, 0.009968495, 0.002999034, 0.02027741, 
    0.006147666, 0.1552106, 0.1721086, 0.2213743, 0.1730296, 0.130021, 
    0.2021611, 0.2041766, 0.1760277, 0.2220149, 0.09124782, 0.1224387, 
    0.09905707, 0.02847971, 0.1007993, 0.02821845, 0.0780338, 0.07536245, 
    0.06324996, 0.1495827, 0.1036389, 0.04265881, 0.09021555,
  0.113256, 0.183278, 0.1342876, 0.1918015, 0.1628844, 0.1789074, 0.1186657, 
    0.008646239, 0.004281426, 0.03120235, 0.09798935, 0.07960898, 0.1269927, 
    0.1952625, 0.1000208, 0.1366013, 0.1401793, 0.1394769, 0.1426218, 
    0.04557967, 0.1031535, 0.1108931, 0.1338908, 0.1375806, 0.08278847, 
    0.105584, 0.1750372, 0.1314647, 0.1248931,
  0.1790768, 0.1580655, 0.1241579, 0.106043, 0.09834845, 0.09099761, 
    0.1186565, 0.07704704, 0.07013533, 0.1535662, 0.05749397, 0.08584588, 
    0.09289791, 0.09964728, 0.02802468, 0.07574122, 0.09694967, 0.2084951, 
    0.1824493, 0.1333244, 0.1180526, 0.1708838, 0.09399559, 0.1209097, 
    0.2441412, 0.2591712, 0.2228699, 0.1266412, 0.1991715,
  0.09614106, 0.1112062, 0.1497199, 0.08897888, 0.1274874, 0.1308124, 
    0.1183132, 0.1065893, 0.01191983, 0.02393799, 0.03416603, 0.06639611, 
    0.06056685, 0.0745258, 0.05941693, 0.06293195, 0.06531101, 0.1794313, 
    0.1185521, 0.1885821, 0.1022083, 0.06260423, 0.07142931, 0.05192422, 
    0.1095969, 0.03283807, 0.02746093, 0.1322254, 0.09443846,
  0.03841753, 0.03950712, 0.07237664, 0.08510326, 0.08142205, 0.03450944, 
    0.003328423, 0.004621934, 0.0002725919, 0.005331518, 0.01604011, 
    0.02744339, 0.03525207, 0.04251073, 0.03541344, 0.03215851, 0.05551466, 
    0.04536576, 0.05247084, 0.04663371, 0.009188371, 0.01427232, 0.005288381, 
    -6.621228e-05, 0.005124596, 0.00841057, 0.008555846, 0.006695222, 
    0.04673808,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0.001665481, 0.006497986, 0.0001110562, 0, 0, 0, 0, 0, 0, 0, 0, 
    -3.74662e-05, -7.770991e-05, 0.01156027, 0.01335373, 0.01441413, 
    0.005479305, -1.467839e-05, 0, 0.0001733713, 0, 0.0002053303, 
    3.567099e-05, 0.0001578324, -1.505592e-05, -2.575796e-07, 0, 0,
  0.003646403, 0.01515054, 0.01397728, 0.01837311, 0.04184015, 0.03382904, 
    0.03647117, 0.03431899, 0.02308535, 0.009005896, 0.009140503, 0.02365163, 
    0.0339165, 0.07794052, 0.07611805, 0.07680155, 0.06787837, 0.04696645, 
    0.03239722, 0.02023903, 0.03471801, 0.03194181, 0.05696547, 0.05923915, 
    0.1075735, 0.06030285, 0.04526216, 0.01645931, 0.00264381,
  0.176716, 0.1609, 0.167648, 0.1642697, 0.2074724, 0.204464, 0.1905534, 
    0.1872442, 0.1729847, 0.1537029, 0.1476854, 0.1940919, 0.16535, 
    0.1882695, 0.1331832, 0.1319283, 0.1168075, 0.1466852, 0.1245876, 
    0.1403838, 0.1227954, 0.1120578, 0.1529595, 0.1370544, 0.1473811, 
    0.09430511, 0.1169009, 0.1743692, 0.1729116,
  0.1515098, 0.1043138, 0.1193874, 0.1438746, 0.1933356, 0.1002131, 
    0.1164703, 0.07833008, 0.04208825, 0.03434794, 0.03965985, 0.0962937, 
    0.07230955, 0.1048297, 0.01929909, 0.05656107, 0.1209419, 0.123187, 
    0.07140738, 0.09734324, 0.189624, 0.1959663, 0.1635587, 0.09277972, 
    0.1526008, 0.125735, 0.1546483, 0.1288339, 0.1771822,
  0.0388226, 0.009144113, 0.05025925, 0.09791359, 0.05763264, 0.02342178, 
    0.004048176, -1.844159e-06, -1.852451e-05, -1.323187e-05, 0.0002176428, 
    0.02434907, 0.01409487, 0.003307286, 0.06842801, 0.1533526, 0.06008324, 
    0.06696894, 0.2024667, 0.108419, 0.02590802, 0.03424528, 0.03010417, 
    0.03025106, 0.06020065, 0.1205397, 0.09795915, 0.06553125, 0.0297402,
  6.16689e-08, 0.01115919, 0.1011297, 0.008317111, 0.02197814, 0.01515589, 
    0.001150939, 0.01928466, 2.013196e-06, -5.944177e-10, -6.126944e-06, 
    5.756481e-08, -5.775764e-08, 0.005431116, 0.06186699, 0.1004234, 
    0.07743274, 0.0380358, 0.001862655, -8.236935e-08, 0, 1.153467e-08, 
    2.605392e-09, 0.07400607, 0.08859423, 0.1010078, -0.0006398573, 
    0.005598856, -1.221778e-06,
  2.051243e-08, -2.719186e-05, 0.01009095, 9.494153e-05, 7.857521e-05, 
    0.0006113992, 0.02106162, 0.114261, 0.0282636, 1.701337e-05, 
    0.0003075156, 0.003623484, 0.04097855, 0.1398588, 0.07091236, 0.02906309, 
    0.001475605, -4.230583e-07, 3.569994e-07, 5.735322e-09, 2.400139e-08, 
    5.512046e-07, 2.911158e-07, 0.09243531, 0.09388757, 1.18836e-06, 
    3.202365e-08, 2.776233e-08, 1.094658e-07,
  0.001333857, 0.2491175, 0.09133645, 2.605421e-06, 0.000973227, 0.03157583, 
    0.08995514, 0.1236602, 0.1280992, 0.1221501, 0.0630023, 0.1068498, 
    0.0233051, 0.02984647, 0.007515262, 0.0001622168, 9.608115e-06, 
    7.254634e-07, 1.084047e-06, 5.734463e-06, 5.590766e-06, 0.006454921, 
    0.03265821, 0.09598032, 0.007943222, -0.0001481705, 9.495468e-06, 
    2.39474e-05, 1.596921e-06,
  0.1149189, 0.06521723, 0.04817744, 0.006557402, 0.0001718059, 0.005941661, 
    0.02182809, 0.04303606, 0.09721717, 0.06357566, 0.02675529, 0.04432452, 
    0.1375019, 0.1431406, 0.1150287, 0.1170984, 0.05812492, 0.02133831, 
    0.04266934, 0.1549284, 0.07247888, 0.3196973, 0.13065, 0.03918087, 
    0.05244529, 0.02458197, 0.06604714, 0.1154952, 0.09080546,
  -9.56382e-05, 6.151099e-05, 2.383796e-06, 1.035186e-06, 7.666606e-07, 
    0.002640935, 0.1323256, 0.03273151, 0.05261422, 0.01321506, 0.0767655, 
    0.04033551, 0.1206498, 0.01715266, 0.008847371, 0.05878117, 0.02726847, 
    -1.541262e-05, 4.396728e-08, 0.003877907, 0.06255717, 0.1063857, 
    0.01929462, 0.03402334, 0.01381027, 0.05381169, 0.07792979, 0.1154978, 
    0.007335782,
  0.06713249, 0.002923877, 2.626989e-06, 8.973369e-07, -1.058453e-06, 
    -2.531385e-10, 0.0001632516, 0.08067789, 0.1534965, 0.08932357, 
    0.04484399, 0.01293956, 0.06510401, 0.09302108, 0.01655281, 0.05539398, 
    0.03745532, 0.01535448, 0.0003161492, 0.01479218, 0.01756696, 0.07789392, 
    0.1306585, 0.0453782, 0.0535138, 0.03667777, 0.04427075, 0.01615313, 
    0.093279,
  0.1284072, 0.07814001, 0.01707768, 0.01225562, 0.003549827, 0.0208626, 
    0.02379978, 0.1435589, 0.1646451, 0.2083716, 0.1629854, 0.1199268, 
    0.1823664, 0.1852935, 0.1848298, 0.2165472, 0.07681804, 0.1054334, 
    0.06947447, 0.02329578, 0.08001672, 0.01861729, 0.09170962, 0.0598255, 
    0.05338148, 0.1451243, 0.1085344, 0.03558697, 0.08277873,
  0.09116615, 0.1920266, 0.1247451, 0.1819542, 0.126183, 0.1547977, 
    0.1412251, 0.06730326, 0.05711397, 0.09259317, 0.1411371, 0.1022863, 
    0.2060594, 0.2314051, 0.1155804, 0.159961, 0.1667948, 0.1450733, 
    0.1252846, 0.05118232, 0.1002111, 0.1008389, 0.1325976, 0.161827, 
    0.08484297, 0.1125858, 0.1452446, 0.1359568, 0.09581557,
  0.1809939, 0.1713749, 0.126977, 0.1229849, 0.1448451, 0.1176489, 0.1080128, 
    0.2050285, 0.1246637, 0.2378747, 0.1060566, 0.1194898, 0.1195038, 
    0.1233755, 0.05183664, 0.1317279, 0.1693308, 0.2807421, 0.2622997, 
    0.1819184, 0.1680616, 0.1904678, 0.1327661, 0.1482965, 0.2884365, 
    0.2514272, 0.2128143, 0.1520688, 0.182034,
  0.2224747, 0.2043043, 0.1798591, 0.08172859, 0.1464425, 0.1759668, 
    0.1596517, 0.160651, 0.07420889, 0.1018101, 0.1477646, 0.1150289, 
    0.142774, 0.1398679, 0.05687871, 0.09088484, 0.1559546, 0.2177694, 
    0.1559893, 0.2697896, 0.1699657, 0.2104601, 0.1618275, 0.1155856, 
    0.1405306, 0.04326006, 0.03301794, 0.1895788, 0.2086562,
  0.0966699, 0.07348852, 0.08293358, 0.1518672, 0.1736197, 0.1362632, 
    0.1166448, 0.08906913, 0.08365844, 0.08442368, 0.07117583, 0.06420395, 
    0.0479103, 0.06781632, 0.07760199, 0.1326108, 0.1723145, 0.1901798, 
    0.2376022, 0.1681275, 0.07866634, 0.09452865, 0.03687594, -0.005698027, 
    0.02264418, 0.00858927, 0.007969439, 0.00713607, 0.1201284,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0003945547, -5.913019e-05, 0, 0, 0, 0,
  0.002830535, 0.01466665, 0.01381115, 0.005517603, -1.84707e-05, 0, 
    -3.389049e-05, 0, 0, 0, 0, 0, 0.0005025529, 0.008154538, 0.03383303, 
    0.02138069, 0.01617233, 0.01477085, 0.01055332, 0.001242558, 0.009524498, 
    0.005953109, 0.009928228, 0.01461325, 0.02702, 0.0568931, 0.03296849, 
    0.001181322, 0,
  0.05691278, 0.06512037, 0.05543577, 0.0685795, 0.1201104, 0.1061506, 
    0.09191363, 0.0739151, 0.0571017, 0.01825305, 0.05651582, 0.1118762, 
    0.1778767, 0.1715175, 0.1625515, 0.1699246, 0.1939109, 0.1449245, 
    0.095032, 0.1225832, 0.1006754, 0.1312391, 0.1538033, 0.1322098, 
    0.1941058, 0.1369189, 0.09311458, 0.06413618, 0.0517075,
  0.2091613, 0.1861367, 0.20635, 0.1834534, 0.2200508, 0.2151698, 0.2100745, 
    0.2198648, 0.2049903, 0.225918, 0.1975655, 0.2505331, 0.1854136, 
    0.1955066, 0.1492144, 0.140778, 0.1181316, 0.1604346, 0.1655887, 
    0.2049074, 0.1882, 0.1777274, 0.1979479, 0.1922088, 0.1813449, 0.156847, 
    0.2033026, 0.2315145, 0.2237491,
  0.139761, 0.1012788, 0.1014496, 0.1124993, 0.1396901, 0.07544945, 
    0.1128114, 0.07223526, 0.02530574, 0.02804062, 0.0455879, 0.09655574, 
    0.06359697, 0.0978198, 0.0152454, 0.06043104, 0.1135278, 0.1279488, 
    0.0822801, 0.09997538, 0.1833483, 0.1888731, 0.1685121, 0.1180653, 
    0.1085102, 0.1230986, 0.1335419, 0.1189135, 0.1713705,
  0.0283114, 0.008970227, 0.04154268, 0.0792999, 0.05560498, 0.0218902, 
    1.704922e-05, -5.62062e-06, -3.314344e-06, 4.413198e-06, 0.003575724, 
    0.05082241, 0.02008228, 0.009606564, 0.05034628, 0.1437986, 0.06128904, 
    0.0478295, 0.1895709, 0.08633845, 0.02535409, 0.02569992, 0.02374538, 
    0.02058368, 0.05900165, 0.1152478, 0.08859055, 0.05770925, 0.03027456,
  -1.273848e-09, 0.007836474, 0.08962404, 0.004451544, 0.01435204, 
    0.006409078, 0.001631215, 0.02049508, 7.05268e-07, 6.007241e-09, 
    0.0001531115, 8.570544e-08, -2.371471e-07, 0.005269486, 0.06147394, 
    0.1112206, 0.06734609, 0.02702444, 0.001015756, -1.433614e-08, 0, 
    7.254589e-08, 2.089331e-08, 0.07683588, 0.06344341, 0.08515002, 
    0.005101032, 0.0001777777, 1.171229e-07,
  -4.743343e-09, -0.0001471457, 0.007001095, 8.813959e-05, 0.000184849, 
    0.0006113608, 0.02086853, 0.1267873, 0.02816122, 0.0001359476, 
    0.0006452436, 0.01419598, 0.06665932, 0.1603513, 0.05236672, 0.02435519, 
    0.0011948, -3.116651e-07, 1.141701e-07, -8.532496e-11, -1.233613e-09, 
    3.752497e-08, 7.930958e-05, 0.08344711, 0.06018432, 8.661887e-06, 
    -2.375931e-09, 8.771265e-10, 1.443087e-08,
  0.01472059, 0.2125553, 0.06831576, 4.65192e-06, 0.001340095, 0.02857837, 
    0.08313429, 0.1028051, 0.07947861, 0.1315824, 0.07467978, 0.09599564, 
    0.01945824, 0.02723057, 0.008351337, 0.001110574, -2.186693e-06, 
    4.906513e-07, 6.967284e-07, 2.197417e-06, 1.280118e-06, 0.00696778, 
    0.02179933, 0.06011819, 0.01017124, 4.422065e-05, 2.737058e-06, 
    -0.0001112187, 1.388039e-05,
  0.09686599, 0.05522849, 0.0458561, 0.004671501, 0.0004178095, 0.00497845, 
    0.01639011, 0.02741603, 0.06390207, 0.0677324, 0.01742217, 0.02858326, 
    0.1156808, 0.1354637, 0.1042725, 0.1187477, 0.05417677, 0.01876799, 
    0.05532709, 0.1884674, 0.05569096, 0.2816816, 0.1261706, 0.02942342, 
    0.0573935, 0.02046157, 0.06761108, 0.1033916, 0.07993924,
  0.0003487703, 3.571287e-05, 2.320068e-06, -6.960872e-07, 4.400274e-07, 
    -4.899674e-05, 0.1189874, 0.02431669, 0.05442821, 0.01217221, 0.07143868, 
    0.03732971, 0.1065869, 0.01595855, 0.007368268, 0.05975763, 0.006238562, 
    -3.606333e-05, 9.763183e-08, 0.004666646, 0.06242967, 0.09733105, 
    0.01300495, 0.02594731, 0.0102066, 0.05064828, 0.08150902, 0.09850663, 
    0.001153684,
  0.04544021, 0.00157597, 9.68144e-07, 1.91104e-07, -3.327874e-07, 
    8.109999e-05, 0.0004315102, 0.08772559, 0.1722404, 0.1128308, 0.04634593, 
    0.01552392, 0.04526269, 0.0967474, 0.01720058, 0.0450913, 0.01417, 
    0.006986462, 7.36031e-05, 0.01844376, 0.01368648, 0.0666266, 0.1040535, 
    0.028589, 0.03922015, 0.02599086, 0.03517189, 0.005224343, 0.1004524,
  0.1078312, 0.08129637, 0.01776794, 0.01372921, 0.008690442, 0.02597382, 
    0.05591067, 0.1177819, 0.1424917, 0.1696632, 0.152944, 0.1009572, 
    0.1578728, 0.1744224, 0.1762536, 0.215462, 0.07561974, 0.09005194, 
    0.07271554, 0.02506231, 0.06564151, 0.0152072, 0.09313335, 0.0595018, 
    0.05716562, 0.1416505, 0.1083907, 0.02550007, 0.06157345,
  0.08349067, 0.1772575, 0.1303095, 0.1636949, 0.1158285, 0.1275866, 
    0.1286308, 0.1376744, 0.1178142, 0.1749424, 0.1469214, 0.1187226, 
    0.2020918, 0.2249994, 0.1118998, 0.1736551, 0.1722195, 0.1513232, 
    0.1057858, 0.04786517, 0.09278622, 0.0939692, 0.1323165, 0.1655675, 
    0.08575747, 0.1011716, 0.1449653, 0.1323315, 0.09183482,
  0.1570705, 0.2399547, 0.1160617, 0.1293802, 0.1578281, 0.1135055, 
    0.1019344, 0.2170872, 0.1797052, 0.2659624, 0.1033321, 0.1309275, 
    0.1458739, 0.1442164, 0.08870626, 0.2271176, 0.2568878, 0.3407071, 
    0.3198972, 0.2380797, 0.1551058, 0.172306, 0.1403783, 0.1802984, 
    0.3412973, 0.2474449, 0.2082444, 0.1348988, 0.1575416,
  0.2665653, 0.217798, 0.2422153, 0.1918072, 0.1968729, 0.1853846, 0.1877551, 
    0.2282721, 0.126951, 0.1853256, 0.1805936, 0.1881601, 0.1900625, 
    0.190898, 0.0934078, 0.09973861, 0.1858987, 0.2425814, 0.199147, 
    0.2472508, 0.1716979, 0.191255, 0.1733499, 0.1252634, 0.175801, 0.111309, 
    0.03634754, 0.1691044, 0.3030868,
  0.2052532, 0.1662178, 0.142913, 0.235379, 0.2391613, 0.1440362, 0.1308563, 
    0.1436178, 0.1347297, 0.1865915, 0.1715346, 0.127387, 0.09408338, 
    0.1213127, 0.1915152, 0.2336433, 0.2246112, 0.284127, 0.2448419, 
    0.2455286, 0.1932377, 0.1704085, 0.1040703, 0.07668338, 0.07607693, 
    0.03043619, 0.01614271, 0.07162787, 0.2050383,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0006221674, 0.009894222, 
    0.01246836, -0.0003257772, 0, 0, 0, 0, 2.432515e-06, 0.01816609, 
    0.02122493, -0.00209801, 0, 0, 0,
  0.01911864, 0.02967228, 0.03746058, 0.013054, -0.0002862806, -2.326257e-05, 
    0.009424954, 0, 0, 0, 0, 0, 0.01049508, 0.06532964, 0.1014256, 
    0.08924621, 0.07413227, 0.06045419, 0.08236003, 0.07394987, 0.1264323, 
    0.1237082, 0.1746768, 0.1491834, 0.2136264, 0.1634729, 0.09947067, 
    0.03633438, 0.02531421,
  0.1106078, 0.1204498, 0.1153019, 0.1533815, 0.1372684, 0.1481735, 
    0.1271116, 0.09625421, 0.1010936, 0.09924089, 0.1188149, 0.1795889, 
    0.252371, 0.2403406, 0.2086899, 0.2127157, 0.2546011, 0.235064, 
    0.1546547, 0.169848, 0.2046709, 0.217974, 0.3000932, 0.2178931, 
    0.2740302, 0.1910277, 0.1553595, 0.09881951, 0.1409358,
  0.2288162, 0.2508863, 0.2261794, 0.1939505, 0.1974197, 0.1974806, 
    0.2084972, 0.2284087, 0.1950303, 0.2632116, 0.2289684, 0.2528588, 
    0.1950387, 0.1897441, 0.150538, 0.136391, 0.1250419, 0.153144, 0.1720158, 
    0.2484435, 0.2312209, 0.2162579, 0.2258729, 0.2091233, 0.1909467, 
    0.1666069, 0.2139347, 0.2376334, 0.2406055,
  0.1268418, 0.08903645, 0.09194123, 0.09192293, 0.1009891, 0.06520941, 
    0.108946, 0.07261185, 0.02638366, 0.02637365, 0.04929265, 0.0941118, 
    0.0612746, 0.09106065, 0.01409573, 0.06896718, 0.110378, 0.1165032, 
    0.09279878, 0.1076516, 0.1828674, 0.1845952, 0.1522174, 0.120619, 
    0.0704288, 0.1187765, 0.1328175, 0.1080176, 0.1643851,
  0.01637193, 0.009453892, 0.05131555, 0.06534939, 0.0449523, 0.005725294, 
    -4.490324e-05, -0.0002639282, 0.001156519, 5.603285e-06, 0.01002217, 
    0.06294086, 0.03060392, 0.02686096, 0.04718356, 0.1272778, 0.07765582, 
    0.04749491, 0.1914555, 0.09249086, 0.02837223, 0.01084683, 0.005910534, 
    0.0211212, 0.05364975, 0.1208564, 0.08170867, 0.0576578, 0.02270151,
  -4.972477e-10, 0.004889738, 0.08124286, 0.001740273, 0.009845812, 
    0.0008704889, 0.006243653, 0.03396863, -1.167939e-05, 9.592428e-07, 
    1.007641e-05, 6.36221e-07, -5.386105e-07, 0.000485791, 0.0709713, 
    0.09946219, 0.05377553, 0.03975341, 0.002392245, -1.313388e-09, 0, 
    7.670469e-08, -1.151478e-07, 0.05052848, 0.04786193, 0.0684212, 
    0.01107944, -3.858347e-06, 4.579461e-08,
  4.376792e-08, -0.0001692129, 0.005604059, 7.194752e-06, 0.0001074786, 
    0.0006078703, 0.01977926, 0.1085317, 0.02451143, 0.0003711249, 
    0.0005002555, 0.03877765, 0.07366201, 0.15459, 0.0516496, 0.02605005, 
    0.002148221, 1.059394e-05, 3.27239e-08, 0, 2.284495e-09, 1.460691e-09, 
    0.002742801, 0.07536761, 0.03913547, 1.226367e-05, 7.882051e-09, 
    3.153132e-09, 1.848697e-08,
  0.01665686, 0.1886498, 0.06020479, 0.0001280971, 0.01220524, 0.04870319, 
    0.07924979, 0.09118413, 0.05805874, 0.1457121, 0.06855672, 0.0912798, 
    0.02315581, 0.03007241, 0.009501612, 0.004467319, 0.0001026083, 
    -4.115897e-06, 6.879907e-07, 1.664081e-06, 5.328417e-07, 0.0112413, 
    0.03091393, 0.05248701, 0.01989309, 0.0007652068, 0.0008316398, 
    8.169514e-06, 0.003169714,
  0.08158189, 0.04535376, 0.04705212, 0.005711269, 0.0001767936, 0.004643092, 
    0.01499019, 0.02152344, 0.06756788, 0.06207528, 0.01176044, 0.01875083, 
    0.1012378, 0.1264371, 0.1097897, 0.116308, 0.05248587, 0.01978386, 
    0.04904268, 0.2095821, 0.06615921, 0.2503993, 0.117067, 0.02673474, 
    0.05680081, 0.02048667, 0.08304778, 0.1012612, 0.0695563,
  0.01101599, 1.244389e-05, 4.304486e-06, 1.119276e-05, 1.041802e-07, 
    -4.743223e-07, 0.1109333, 0.01857677, 0.05467284, 0.01359875, 0.07666727, 
    0.0364088, 0.1017081, 0.01735914, 0.006190205, 0.04672021, 0.002307236, 
    -1.549223e-06, -4.585963e-08, 0.008859262, 0.06105516, 0.1015274, 
    0.01065316, 0.02263866, 0.008291737, 0.05035951, 0.08707385, 0.0589418, 
    0.0006086453,
  0.03851922, 0.003322992, 3.133901e-05, 6.18346e-08, -3.494867e-06, 
    0.005087956, 0.000184109, 0.1061283, 0.1891625, 0.1353174, 0.04885122, 
    0.02366568, 0.04070651, 0.08848648, 0.02620181, 0.03724933, 0.0132655, 
    0.002331898, 0.0005495053, 0.002606407, 0.01373681, 0.04883011, 
    0.09134932, 0.02357376, 0.02924159, 0.01880483, 0.03532524, 0.003091557, 
    0.1035252,
  0.08915804, 0.09195979, 0.01254053, 0.01249137, 0.02173845, 0.02909328, 
    0.07629405, 0.09172527, 0.1172281, 0.1232556, 0.1306246, 0.09304038, 
    0.1352372, 0.1583324, 0.1545792, 0.1851211, 0.06575672, 0.07491039, 
    0.05362685, 0.0250716, 0.05656092, 0.02052089, 0.08470759, 0.05518209, 
    0.03963117, 0.1389837, 0.1000299, 0.01268347, 0.05081712,
  0.07788865, 0.1562209, 0.1394423, 0.1518509, 0.1148398, 0.1162059, 
    0.1089227, 0.1638101, 0.2053689, 0.1652982, 0.1288231, 0.1110204, 
    0.2006712, 0.2192701, 0.110536, 0.1643829, 0.1585634, 0.1705979, 
    0.0881902, 0.04206812, 0.08892847, 0.07990836, 0.1254287, 0.1620819, 
    0.09259846, 0.1104747, 0.1453612, 0.1255689, 0.09640251,
  0.169273, 0.2443238, 0.1174821, 0.1098993, 0.1511278, 0.1081052, 
    0.08695856, 0.2067917, 0.1947738, 0.2480556, 0.1099734, 0.1387012, 
    0.14345, 0.1555363, 0.1243497, 0.24226, 0.2430033, 0.3709829, 0.3732179, 
    0.2163105, 0.1259551, 0.1579155, 0.1457439, 0.2010631, 0.3362441, 
    0.2511678, 0.22315, 0.1363138, 0.1326005,
  0.2482042, 0.2100568, 0.2524469, 0.2073976, 0.2480982, 0.237372, 0.2087324, 
    0.2375073, 0.1706502, 0.2270076, 0.1839418, 0.1883325, 0.1914446, 
    0.2303366, 0.1287893, 0.08773284, 0.1953999, 0.2364393, 0.1863057, 
    0.2233011, 0.1481709, 0.1852013, 0.1560047, 0.1363062, 0.156514, 
    0.1336301, 0.05831983, 0.1496045, 0.2933029,
  0.2272304, 0.2057678, 0.1844337, 0.2140631, 0.2522022, 0.1805187, 
    0.1569436, 0.186301, 0.1919083, 0.256191, 0.2480538, 0.2433121, 
    0.1870876, 0.1501122, 0.2113194, 0.2687799, 0.279413, 0.2967407, 
    0.2380129, 0.2549623, 0.226732, 0.1857026, 0.1483359, 0.1399462, 
    0.1489713, 0.08630453, 0.07243743, 0.1068974, 0.2389906,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01101346, 0.07396509, 0.08156186, 
    0.06361921, 0.02466682, 0.001100985, 2.635689e-05, 0, 0, 0.00405192, 
    0.1012879, 0.1253427, 0.01970686, 0.06047835, -0.0012504, 0,
  0.0669033, 0.07756995, 0.1596124, 0.06443169, -0.0006392789, -0.00054435, 
    0.03397123, -0.0001474808, -1.408183e-08, -2.251903e-05, 1.00424e-05, 
    -4.506805e-05, 0.02613871, 0.1158888, 0.1379064, 0.1328792, 0.1554851, 
    0.2108308, 0.2661105, 0.2328767, 0.2669865, 0.2647299, 0.2798488, 
    0.3087005, 0.3116802, 0.2895496, 0.2489916, 0.094054, 0.1180556,
  0.1537169, 0.1808916, 0.1966998, 0.2069498, 0.242425, 0.2198863, 0.1894811, 
    0.1569836, 0.1329488, 0.1430247, 0.1676894, 0.2722865, 0.3129692, 
    0.286516, 0.2531433, 0.2304616, 0.2796178, 0.3269228, 0.2143779, 
    0.2231043, 0.2559362, 0.2580102, 0.337983, 0.237454, 0.2877424, 
    0.2251088, 0.1945457, 0.1802852, 0.2306596,
  0.2255466, 0.2474906, 0.2172487, 0.1757077, 0.170716, 0.1876086, 0.20075, 
    0.2257538, 0.1967137, 0.2774971, 0.2413054, 0.2524002, 0.2071446, 
    0.1896356, 0.1447892, 0.1238073, 0.1189612, 0.1458896, 0.1812913, 
    0.2665616, 0.2289297, 0.2114086, 0.2292788, 0.2014639, 0.1667738, 
    0.1432525, 0.2065792, 0.2220868, 0.2232035,
  0.1160861, 0.08890778, 0.08479237, 0.08626986, 0.086936, 0.06624696, 
    0.1042638, 0.0660621, 0.03576535, 0.02775118, 0.05002981, 0.08040197, 
    0.05866169, 0.08488473, 0.02453822, 0.07329883, 0.09709274, 0.104262, 
    0.07917646, 0.09755123, 0.1575891, 0.1708403, 0.1284754, 0.1133114, 
    0.05753242, 0.1103915, 0.1186269, 0.123787, 0.1621512,
  0.005098387, 0.01019554, 0.07431482, 0.05730509, 0.04300814, 0.0009923918, 
    1.639248e-06, -0.0001014675, -3.187124e-05, 2.604173e-06, 0.03072627, 
    0.07671279, 0.04340904, 0.04548604, 0.05780246, 0.1142655, 0.07668525, 
    0.04511688, 0.1686614, 0.08730797, 0.01101733, 0.003737773, 0.0001830983, 
    0.02524605, 0.05300996, 0.1251089, 0.08032726, 0.05888281, 0.01383077,
  2.534814e-09, 0.001999732, 0.07986397, 0.007111342, 0.013813, 0.01094976, 
    0.02355358, 0.04233946, -5.298217e-06, 0.0006060962, 3.007691e-08, 
    0.000339012, -2.526419e-07, -1.723586e-05, 0.0754288, 0.0883932, 
    0.02818549, 0.05841309, 0.0009563023, -3.176883e-10, 0, 9.479549e-10, 
    -1.17374e-06, 0.01873386, 0.03551333, 0.05245974, 0.0151945, 
    9.733578e-06, 5.771778e-08,
  7.545287e-08, -2.378319e-05, 0.005891978, 0.0001261854, 0.0001652472, 
    0.0008120104, 0.01890802, 0.09650281, 0.01703955, 0.0002315583, 
    0.0002359947, 0.03158156, 0.085757, 0.123286, 0.05521055, 0.02622225, 
    0.006253532, 3.495486e-06, -5.567712e-10, -2.031803e-10, -4.669564e-11, 
    5.378297e-09, 0.0002922121, 0.05762148, 0.02588356, 3.359251e-05, 
    4.010098e-09, 4.612481e-08, 2.616614e-08,
  0.03623626, 0.1688652, 0.05842264, 0.006591523, 0.0369586, 0.0552783, 
    0.08211497, 0.09090018, 0.04799899, 0.1533388, 0.06169239, 0.08124959, 
    0.01873961, 0.01785641, 0.009165493, 0.004996791, 0.004483268, 
    0.0002398065, 0.004814546, 1.448204e-05, 1.012717e-06, 0.006954161, 
    0.05094261, 0.04113294, 0.01118998, 0.002758582, 0.0002444092, 
    0.005705421, 0.01264219,
  0.07240597, 0.03486664, 0.05593528, 0.009866502, 0.001253384, 0.007382536, 
    0.0184701, 0.01725725, 0.07160011, 0.06813243, 0.01117123, 0.01237878, 
    0.09652982, 0.1184661, 0.106792, 0.116169, 0.05681666, 0.02604221, 
    0.05116053, 0.2516901, 0.09816444, 0.2227933, 0.1183754, 0.02105867, 
    0.05699882, 0.02144501, 0.08309435, 0.09972903, 0.06612218,
  -0.0001302887, 7.379556e-06, 2.011763e-06, 7.467913e-05, 5.922168e-08, 
    0.0002998608, 0.07805456, 0.01803065, 0.05691133, 0.0170799, 0.08115725, 
    0.03841898, 0.09623052, 0.02722308, 0.005282393, 0.03704168, 0.001857312, 
    2.860737e-06, -7.215602e-05, 0.01154489, 0.05193182, 0.1067804, 
    0.008453167, 0.02142938, 0.007136775, 0.05463266, 0.07873252, 0.03640586, 
    0.003370212,
  0.02743774, 0.001022293, 1.060598e-05, 8.931898e-09, -1.343747e-05, 
    0.007894056, 0.0004146069, 0.1219033, 0.2121071, 0.1527562, 0.06176693, 
    0.02858713, 0.03974134, 0.08301143, 0.02184776, 0.03306459, 0.009066288, 
    0.0002681346, 0.0006935063, 0.0002787923, 0.01625284, 0.04389942, 
    0.07974891, 0.02003603, 0.02613402, 0.0190285, 0.03159722, 0.003088297, 
    0.09178793,
  0.09086055, 0.09707637, 0.01282974, 0.013098, 0.04289164, 0.02347665, 
    0.08794698, 0.07536569, 0.09152186, 0.09578463, 0.10647, 0.08456601, 
    0.1107084, 0.1502158, 0.1259182, 0.1622604, 0.08040387, 0.07767351, 
    0.05018786, 0.02919067, 0.06520938, 0.05471847, 0.08254799, 0.05150334, 
    0.03549871, 0.134672, 0.09058864, 0.02178937, 0.05070049,
  0.05542342, 0.1364879, 0.1418394, 0.1515567, 0.1130502, 0.1090434, 
    0.1020942, 0.1575753, 0.2144356, 0.1489323, 0.1239994, 0.1013764, 
    0.1955521, 0.2247754, 0.1071123, 0.1452447, 0.1566873, 0.1753775, 
    0.08541259, 0.0403409, 0.0845804, 0.06913719, 0.1181353, 0.1534089, 
    0.1003958, 0.1051839, 0.1304072, 0.1255626, 0.1073583,
  0.1690532, 0.2291616, 0.1117427, 0.09966579, 0.1380186, 0.109789, 
    0.07520141, 0.1752669, 0.2000235, 0.2285545, 0.09622606, 0.1591911, 
    0.1293381, 0.155039, 0.1297007, 0.2475868, 0.2347138, 0.4207001, 
    0.3611161, 0.1880136, 0.1276427, 0.1635774, 0.1568049, 0.2183182, 
    0.3208438, 0.2624927, 0.2372654, 0.1313946, 0.1274112,
  0.2442247, 0.193372, 0.2644394, 0.2116415, 0.2328784, 0.2557705, 0.2244895, 
    0.3172231, 0.2520569, 0.2724894, 0.1773448, 0.1790627, 0.1904172, 
    0.2381268, 0.1430109, 0.1028588, 0.2308001, 0.2465584, 0.1775612, 
    0.1931945, 0.1537999, 0.1798797, 0.1517082, 0.1499823, 0.1541924, 
    0.1636251, 0.06461154, 0.1400466, 0.2621682,
  0.2184969, 0.2174922, 0.1924317, 0.1847975, 0.2616608, 0.212176, 0.1907759, 
    0.2189664, 0.2076361, 0.2648311, 0.2574466, 0.2466505, 0.200613, 
    0.1519835, 0.2025044, 0.338448, 0.3387267, 0.3041128, 0.2165136, 
    0.2529997, 0.2222461, 0.1756028, 0.1584086, 0.1541157, 0.1570827, 
    0.1606642, 0.1534566, 0.09315137, 0.2498566,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002004698, 0.07834487, 0.114068, 
    0.1697503, 0.1809707, 0.1059613, 0.01244422, 9.909963e-06, 0, 
    -9.433498e-06, 0.0302825, 0.1816014, 0.1846623, 0.1713521, 0.1265238, 
    0.004912191, 0,
  0.1378718, 0.1705835, 0.1825389, 0.127192, -0.001380393, -0.003199937, 
    0.05890749, -0.001731099, 0, -0.0001124005, 2.409733e-05, -0.001095872, 
    0.07274657, 0.2075343, 0.2229754, 0.1662464, 0.195435, 0.2471014, 
    0.3345391, 0.3271593, 0.3156994, 0.2917016, 0.3102527, 0.3438317, 
    0.3591954, 0.3186103, 0.2895312, 0.1291488, 0.181244,
  0.1551291, 0.2243618, 0.2311936, 0.2268675, 0.2907026, 0.285796, 0.2609017, 
    0.2121668, 0.2475716, 0.2655818, 0.2533196, 0.3206559, 0.3110274, 
    0.2750823, 0.2535688, 0.2296128, 0.2891856, 0.3216145, 0.2013395, 
    0.2393672, 0.2687632, 0.2524358, 0.3372325, 0.2465413, 0.2830411, 
    0.2055267, 0.1695791, 0.1612522, 0.2206991,
  0.2266879, 0.253606, 0.1975757, 0.1593432, 0.1622712, 0.1853229, 0.1900793, 
    0.2280756, 0.2153937, 0.2923294, 0.2508365, 0.2581262, 0.2042985, 
    0.1823643, 0.1417037, 0.1257041, 0.09350243, 0.132811, 0.1743025, 
    0.2433772, 0.2100047, 0.2062486, 0.2158659, 0.1870383, 0.1387241, 
    0.1634928, 0.194387, 0.2044835, 0.2016747,
  0.1088511, 0.09933508, 0.06520866, 0.07671324, 0.07411946, 0.06073047, 
    0.08142888, 0.05286955, 0.02988602, 0.02018566, 0.04931026, 0.06444934, 
    0.05599957, 0.08023534, 0.03044927, 0.07045034, 0.09404551, 0.08064602, 
    0.08369564, 0.07033537, 0.1380957, 0.1535947, 0.1344671, 0.1060427, 
    0.05389177, 0.09755939, 0.1023818, 0.1216866, 0.1451093,
  0.006799352, 0.01170686, 0.1081396, 0.056394, 0.03159909, 0.0001037719, 
    1.330604e-06, -2.281567e-05, 2.946941e-05, 2.323747e-07, 0.05989609, 
    0.0932099, 0.04511696, 0.04320144, 0.0594419, 0.09544162, 0.07783885, 
    0.04635753, 0.1473539, 0.08161478, 0.002497898, 0.005814431, 
    -9.014862e-05, 0.02960135, 0.06186447, 0.1273762, 0.07198159, 0.057204, 
    0.01466356,
  3.114269e-08, 0.001521257, 0.08722859, 0.002749479, 0.01119046, 0.04020159, 
    0.0526142, 0.05570808, -1.251939e-06, 4.880972e-06, 1.006298e-07, 
    0.007299447, -7.862425e-06, -0.0002067993, 0.0727024, 0.07388698, 
    0.02021219, 0.06389675, 0.0005077602, 4.435821e-09, 4.241483e-11, 
    2.839955e-10, -3.1171e-06, 0.01688651, 0.0357648, 0.03640289, 0.01871358, 
    -2.628733e-05, 6.447734e-08,
  9.640767e-08, 0.002102397, 0.004869336, 6.044111e-05, 0.0002013082, 
    0.0006562095, 0.02514986, 0.09581944, 0.0111522, 0.0007415649, 
    0.0003800607, 0.02256595, 0.0827983, 0.1176896, 0.04661709, 0.02199306, 
    0.008051537, 0.0001419208, 1.636585e-07, 6.494818e-09, 8.36617e-09, 
    3.069866e-08, 0.007479364, 0.05241129, 0.02487889, 0.0004347352, 
    1.240096e-06, 1.611496e-07, 3.375107e-08,
  0.03358351, 0.1747259, 0.06582638, 0.005111217, 0.03412464, 0.0702924, 
    0.08160704, 0.1117938, 0.06519225, 0.1438165, 0.06376603, 0.07337472, 
    0.02577934, 0.01956679, 0.009298655, 0.005269287, 0.0005178115, 
    0.003994629, 0.01843203, 0.001476431, 0.002245164, 5.745709e-06, 
    0.0530526, 0.04904343, 0.007509794, 0.005614045, 0.002578107, 0.01949947, 
    0.004086979,
  0.0782408, 0.03055602, 0.05811936, 0.02062275, 0.005627143, 0.01005039, 
    0.02243014, 0.03188626, 0.09736793, 0.08419929, 0.01117243, 0.01076503, 
    0.100932, 0.1120195, 0.1048881, 0.1374682, 0.06806002, 0.05684251, 
    0.05337744, 0.2810391, 0.1081394, 0.2153973, 0.1271437, 0.02640042, 
    0.05720885, 0.02061159, 0.09970753, 0.1135444, 0.06312132,
  0.005405259, -1.884302e-05, 1.481555e-06, 0.000221301, -7.472519e-06, 
    0.002393122, 0.08816469, 0.02706347, 0.06145237, 0.02274583, 0.08485238, 
    0.04279657, 0.1024745, 0.0333591, 0.005834017, 0.02487073, 0.002075965, 
    5.021173e-06, -1.384893e-06, 0.01180124, 0.05467134, 0.1030024, 
    0.009166392, 0.02582598, 0.007157865, 0.06288909, 0.07280654, 0.01488584, 
    0.005897327,
  0.02223805, 0.001307336, 5.834966e-06, 3.599074e-10, 0.00469676, 
    0.002281537, 0.000633061, 0.1253676, 0.2289006, 0.1785697, 0.07639542, 
    0.04116215, 0.04283005, 0.0866019, 0.023683, 0.03215078, 0.007583934, 
    0.0002541268, 0.000578251, -2.226002e-05, 0.01947102, 0.02993638, 
    0.08308372, 0.02194778, 0.03018995, 0.02005612, 0.03159378, 0.003059331, 
    0.05112423,
  0.0830962, 0.1242116, 0.0146448, 0.0139312, 0.04266011, 0.01579546, 
    0.1014747, 0.0622755, 0.06741368, 0.07260739, 0.09068594, 0.06923688, 
    0.0864194, 0.144289, 0.1113338, 0.1638409, 0.08053281, 0.08239413, 
    0.03911013, 0.037003, 0.1010962, 0.07943085, 0.1020285, 0.04833907, 
    0.03002015, 0.142057, 0.08451579, 0.02776984, 0.06005702,
  0.03840957, 0.1288705, 0.1419202, 0.1722367, 0.1094661, 0.09774136, 
    0.09490514, 0.1594255, 0.2138675, 0.1352469, 0.1114834, 0.07706288, 
    0.1817595, 0.1921433, 0.1175358, 0.1446117, 0.175532, 0.1848091, 
    0.09828707, 0.04045054, 0.07658713, 0.05893445, 0.1113063, 0.1621016, 
    0.1092248, 0.1204851, 0.1066296, 0.1273494, 0.1106044,
  0.1481803, 0.2227243, 0.1120343, 0.0949718, 0.1459734, 0.1206862, 
    0.06379417, 0.1491678, 0.2138532, 0.2220381, 0.07786409, 0.1575491, 
    0.122205, 0.1697214, 0.1270514, 0.2406799, 0.2270374, 0.4472787, 
    0.3565525, 0.1759125, 0.1114884, 0.1608905, 0.1566388, 0.2871703, 
    0.3057702, 0.2891948, 0.2441948, 0.1344796, 0.1128122,
  0.2752699, 0.2059068, 0.3158559, 0.2255913, 0.1896874, 0.2569157, 
    0.2348472, 0.3284916, 0.2930799, 0.2851469, 0.177944, 0.1790902, 
    0.1857127, 0.2372602, 0.1597452, 0.1005219, 0.2442935, 0.2528518, 
    0.1925228, 0.2213998, 0.1705579, 0.1603024, 0.1788238, 0.1685984, 
    0.1954714, 0.1705607, 0.07534145, 0.1288983, 0.2447007,
  0.2405873, 0.2234711, 0.1925264, 0.2155533, 0.2776149, 0.2241114, 
    0.1798263, 0.2424286, 0.242335, 0.2933748, 0.2820024, 0.2559964, 
    0.2027986, 0.1439092, 0.1993951, 0.3629425, 0.3829402, 0.3135806, 
    0.2169803, 0.2509193, 0.2413598, 0.1982008, 0.1677576, 0.1672679, 
    0.1636213, 0.201665, 0.1749813, 0.08344255, 0.2660829,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.004543521, 0.1172404, 0.2137537, 
    0.2417362, 0.1661263, 0.1557806, 0.06160487, 0.003165253, -0.001134588, 
    -0.0001391634, 0.06968253, 0.1859972, 0.1860633, 0.1738612, 0.1352339, 
    0.027836, 6.477561e-06,
  0.1635917, 0.2551761, 0.2413407, 0.1951836, 0.005838073, 0.01052068, 
    0.07689545, 0.00250993, -0.0003450057, -0.001996513, 0.0007927381, 
    -0.004065052, 0.1525976, 0.2267178, 0.2210722, 0.1960803, 0.2312274, 
    0.2565722, 0.3591867, 0.3451183, 0.3048793, 0.276439, 0.3016299, 
    0.3607627, 0.3768148, 0.2907097, 0.2739096, 0.1142366, 0.184465,
  0.1636288, 0.2436326, 0.2429719, 0.2239197, 0.2982037, 0.3182892, 
    0.2861632, 0.2244398, 0.2737158, 0.299706, 0.268926, 0.3123612, 
    0.2928106, 0.2723992, 0.2500995, 0.2395745, 0.2800002, 0.3045462, 
    0.2040452, 0.2330224, 0.26227, 0.2362178, 0.3071097, 0.2292699, 
    0.2779997, 0.2174179, 0.1882104, 0.1711886, 0.2328025,
  0.2174649, 0.2357814, 0.1863107, 0.1562904, 0.1466663, 0.1833809, 
    0.1977063, 0.226889, 0.2207584, 0.2731052, 0.2608835, 0.2343413, 
    0.2034798, 0.1868258, 0.1395361, 0.120035, 0.08533038, 0.1442072, 
    0.1721378, 0.2299275, 0.222313, 0.1904571, 0.2086365, 0.1711782, 
    0.1172139, 0.1324683, 0.1733647, 0.2100202, 0.1903959,
  0.105849, 0.08358642, 0.07182215, 0.06765721, 0.07414703, 0.06529947, 
    0.07959605, 0.055804, 0.03036327, 0.02575215, 0.05207411, 0.07066307, 
    0.05723887, 0.07734562, 0.03119351, 0.062746, 0.08251385, 0.07141763, 
    0.06512203, 0.05507241, 0.1197867, 0.1472677, 0.1423311, 0.1062483, 
    0.05276963, 0.08766016, 0.0934068, 0.1144115, 0.1343205,
  0.008734897, 0.01884867, 0.1163408, 0.05982888, 0.03166524, 0.002571488, 
    7.42199e-05, -3.413934e-05, 0.0001615038, 3.544876e-07, 0.07254162, 
    0.09606855, 0.04576542, 0.03659943, 0.05850857, 0.09378485, 0.08802838, 
    0.05654139, 0.1485106, 0.06931778, 0.004093932, 0.01099767, 5.173011e-05, 
    0.03575908, 0.09481981, 0.1254734, 0.0693454, 0.06828929, 0.01979313,
  1.008831e-07, 0.001001211, 0.07476605, 0.001188241, 0.01261657, 0.05987082, 
    0.06987701, 0.07685707, -4.752461e-06, 6.078825e-08, 0.0004038161, 
    0.02120896, 0.002353746, -0.0005541802, 0.08898669, 0.07280461, 
    0.01930813, 0.07711811, 0.00033703, 2.227184e-08, 5.463306e-10, 
    1.887097e-09, -3.872338e-08, 0.009417388, 0.03856109, 0.04016274, 
    0.01690007, -2.023449e-05, 1.466702e-07,
  1.894297e-06, 0.01089501, 0.01951325, 6.605389e-05, 0.0002982303, 
    0.00192908, 0.04141592, 0.1207373, 0.007239463, 0.0007800474, 0.00024795, 
    0.02341506, 0.1006111, 0.1286961, 0.06607359, 0.03071126, 0.01017399, 
    0.0006763614, 4.132471e-06, 5.23147e-08, 5.11544e-08, 1.209876e-07, 
    7.48499e-05, 0.06222536, 0.03407022, 0.01085669, -1.107607e-05, 
    1.668018e-06, 2.608376e-07,
  0.03070647, 0.1964467, 0.1037795, 0.001885694, 0.02789744, 0.07965771, 
    0.09331533, 0.1300832, 0.1112996, 0.1385802, 0.08092929, 0.08045038, 
    0.03512182, 0.02138542, 0.009872994, 0.006556048, 0.001188381, 
    0.01209098, 0.01969745, 0.008484785, 0.0004140557, -0.0001275933, 
    0.05457804, 0.067646, 0.008137644, 0.009413224, 0.004152138, 0.01757618, 
    0.003399674,
  0.0901437, 0.03979567, 0.0644078, 0.03642206, 0.01038146, 0.01251597, 
    0.03377397, 0.0516196, 0.1705877, 0.1315705, 0.02363423, 0.01633044, 
    0.1152806, 0.1123485, 0.1256432, 0.1715584, 0.07168348, 0.07185839, 
    0.05986182, 0.3190586, 0.1574628, 0.2451486, 0.152409, 0.03451883, 
    0.06473505, 0.0301518, 0.1224416, 0.1305263, 0.08039156,
  0.008702842, 0.001050383, 8.66225e-07, 0.0002470745, -5.048087e-05, 
    0.0003087036, 0.1380445, 0.0544754, 0.0905779, 0.02412257, 0.0879372, 
    0.04556715, 0.1229438, 0.0419012, 0.008509584, 0.02397116, 0.002523709, 
    3.1167e-06, 9.13705e-07, 0.01636313, 0.07055794, 0.1186467, 0.01375995, 
    0.04193653, 0.0105104, 0.06975792, 0.06831991, 0.01669795, 0.003422575,
  0.02275667, 0.01669255, 4.679999e-06, 2.854904e-10, 0.0009268796, 
    0.0001263818, 0.0009409161, 0.1422668, 0.2567361, 0.189907, 0.08722878, 
    0.04941507, 0.06048089, 0.1009549, 0.02792671, 0.03513212, 0.008798315, 
    0.0002797742, 0.006752421, 5.261428e-05, 0.03182952, 0.02941998, 
    0.0860574, 0.0262629, 0.03655079, 0.0239279, 0.03945069, 0.004473556, 
    0.03394721,
  0.05791153, 0.09114243, 0.01231056, 0.02295571, 0.02953987, 0.01176131, 
    0.1144002, 0.05255598, 0.05048358, 0.05767721, 0.0758011, 0.05588226, 
    0.07583326, 0.1450377, 0.1133381, 0.1656602, 0.08376114, 0.0790736, 
    0.03703867, 0.03110077, 0.09684609, 0.0693497, 0.09583526, 0.04287212, 
    0.02095507, 0.1474678, 0.09109423, 0.04497932, 0.0538392,
  0.04611087, 0.1269292, 0.1398491, 0.1623043, 0.1040583, 0.0870831, 
    0.08608814, 0.1486253, 0.2137862, 0.1327431, 0.1082728, 0.09360191, 
    0.2012969, 0.199483, 0.1253731, 0.1680677, 0.1619154, 0.1798465, 
    0.1134344, 0.04204854, 0.06819663, 0.06737339, 0.1313158, 0.1601089, 
    0.1110503, 0.1097598, 0.08729278, 0.1275371, 0.1123909,
  0.172543, 0.214183, 0.1207382, 0.1061511, 0.1833063, 0.1257383, 0.06872949, 
    0.126924, 0.2214674, 0.2053259, 0.07006092, 0.1736049, 0.09657204, 
    0.1481808, 0.1375343, 0.224009, 0.2347817, 0.4488882, 0.3462457, 
    0.153711, 0.102169, 0.1501015, 0.1636684, 0.2866778, 0.3422682, 
    0.3046105, 0.2006955, 0.1194823, 0.1090182,
  0.3070761, 0.2248137, 0.3441812, 0.241018, 0.1650665, 0.2619221, 0.2420494, 
    0.3358269, 0.311258, 0.2705988, 0.1972159, 0.1843904, 0.1833458, 
    0.215191, 0.1683286, 0.1126228, 0.274541, 0.2630132, 0.2043563, 
    0.2276159, 0.1608792, 0.1807216, 0.1877084, 0.1816342, 0.203077, 
    0.1892005, 0.1150292, 0.1162123, 0.2454955,
  0.2477552, 0.2231117, 0.2150164, 0.1885585, 0.2474684, 0.2203029, 
    0.1729289, 0.297994, 0.2966121, 0.3228413, 0.2867184, 0.2637723, 
    0.2459777, 0.1377852, 0.2093878, 0.4001459, 0.431487, 0.3405414, 
    0.2578014, 0.2822984, 0.266367, 0.1878973, 0.1985303, 0.1835677, 
    0.1857036, 0.1918239, 0.1611989, 0.09130574, 0.2668045,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  -0.0005570832, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01692027, 0.1623898, 
    0.2040262, 0.2109015, 0.1530037, 0.1502126, 0.1050384, 0.1181186, 
    0.02900444, 0.01280251, 0.1922966, 0.1904521, 0.1890518, 0.1669859, 
    0.1332399, 0.0621181, 0.01247951,
  0.1973523, 0.3193837, 0.2496545, 0.2326527, 0.02394811, 0.02632768, 
    0.101619, 0.007661106, -0.0008890003, -0.007273511, 0.005950481, 
    0.0002785411, 0.2083704, 0.2332321, 0.2130768, 0.2032589, 0.2541122, 
    0.2658127, 0.3682061, 0.3785056, 0.3229443, 0.2538976, 0.2989451, 
    0.3605773, 0.4026634, 0.3012253, 0.2626201, 0.1207145, 0.1795593,
  0.1484758, 0.2453373, 0.242379, 0.2122274, 0.3025715, 0.312036, 0.3003308, 
    0.2216254, 0.2765636, 0.2908409, 0.2751719, 0.310371, 0.278636, 
    0.2567807, 0.2434984, 0.2409768, 0.2661613, 0.2680873, 0.2014446, 
    0.234063, 0.2787075, 0.2363543, 0.2862535, 0.233583, 0.275046, 0.2042196, 
    0.1834401, 0.1494417, 0.2334774,
  0.2086642, 0.2298885, 0.1798078, 0.1517657, 0.1447503, 0.1896618, 
    0.1996937, 0.2230443, 0.2206921, 0.2557093, 0.256207, 0.2424611, 
    0.2173203, 0.1711057, 0.1498254, 0.1348691, 0.08463875, 0.1491437, 
    0.1500397, 0.2150666, 0.2180666, 0.1780149, 0.2064466, 0.1624954, 
    0.09267811, 0.1363352, 0.1449319, 0.1811935, 0.1780243,
  0.1144555, 0.08319327, 0.08656547, 0.06961887, 0.08233921, 0.06849009, 
    0.07684381, 0.06888233, 0.03908662, 0.02741695, 0.05526216, 0.06833176, 
    0.05242487, 0.07188509, 0.02972745, 0.05360764, 0.08532142, 0.06280755, 
    0.06295555, 0.04851589, 0.1045796, 0.1360699, 0.139967, 0.1137696, 
    0.04999318, 0.07863097, 0.0760056, 0.1101246, 0.1248421,
  0.006835034, 0.02353477, 0.0971382, 0.05648816, 0.04817514, 0.01029193, 
    7.896403e-05, 4.928192e-05, 0.0006253857, 9.382943e-08, 0.0550372, 
    0.06779933, 0.05810362, 0.04425225, 0.05876028, 0.1112058, 0.08290248, 
    0.0552034, 0.1502845, 0.06580233, 0.006816951, 0.01404705, 0.00939722, 
    0.04657891, 0.1149668, 0.1166136, 0.06088499, 0.0583316, 0.02388981,
  1.690229e-07, 0.00681548, 0.08372876, 0.0008100033, 0.01334826, 0.06746586, 
    0.07467651, 0.06167147, 1.095549e-06, -6.410112e-09, 0.01880907, 
    0.01708468, 0.000906986, 0.01416237, 0.09378529, 0.07846929, 0.02752963, 
    0.0895215, 0.004649818, 2.942998e-08, 4.210639e-09, 1.238946e-08, 
    9.662687e-09, 0.005525505, 0.04089037, 0.07494639, 0.02619589, 
    0.0001933271, 2.599091e-07,
  3.511526e-05, 0.02635651, 0.1214041, 0.0001956129, 0.0003284934, 
    0.005636842, 0.04728894, 0.1302472, 0.009241664, 0.001053751, 
    0.0007576325, 0.03700272, 0.1141252, 0.1499339, 0.08723713, 0.03652877, 
    0.007814556, 0.002048504, 9.577668e-05, 9.091723e-08, 8.24078e-08, 
    1.451389e-07, 0.001720973, 0.07228135, 0.04639795, 0.08119678, 
    2.582808e-05, 2.691973e-06, 3.424518e-07,
  0.03378442, 0.2439662, 0.1681521, 0.001704532, 0.01833321, 0.0782431, 
    0.1093256, 0.1645639, 0.1397278, 0.1646779, 0.08785329, 0.08411702, 
    0.04010001, 0.02623614, 0.005931395, 0.004650693, 0.0004699049, 
    0.002211828, 0.01571316, 0.0003550605, 0.0001588372, 0.001536187, 
    0.0599106, 0.09503096, 0.01266591, 0.003894721, 0.001885672, 0.005315273, 
    0.01535675,
  0.1140238, 0.06324208, 0.07437497, 0.08087684, 0.006941554, 0.007461076, 
    0.043908, 0.05884835, 0.2071725, 0.1456833, 0.04534745, 0.02516969, 
    0.1276452, 0.1070177, 0.1556389, 0.1848874, 0.07552794, 0.09485602, 
    0.07110523, 0.3436519, 0.1939268, 0.2740133, 0.1797301, 0.04194754, 
    0.06363884, 0.03627774, 0.1394785, 0.157702, 0.1121461,
  0.0008538531, 0.0001876896, 2.540817e-06, -7.601637e-08, 0.004387491, 
    2.492787e-06, 0.1893855, 0.07839298, 0.1480689, 0.03100426, 0.09078179, 
    0.04951918, 0.1329802, 0.04648183, 0.01030686, 0.02570572, 0.00341918, 
    7.477811e-07, 7.612746e-07, 0.01971039, 0.07851772, 0.1352834, 
    0.01491777, 0.06041212, 0.01156663, 0.07132794, 0.08189793, 0.01060604, 
    0.01233494,
  0.00500271, 0.004851322, 2.112905e-05, 8.720816e-09, 0.001910207, 
    -2.21156e-05, 0.0004394186, 0.1911482, 0.2591277, 0.2087464, 0.102106, 
    0.05976345, 0.06511959, 0.09511638, 0.02959712, 0.04282411, 0.01260331, 
    0.0006778405, 0.0002014141, 0.0002139263, 0.0516958, 0.03652306, 
    0.09032422, 0.02710091, 0.03703682, 0.02823785, 0.04396769, 0.005140994, 
    0.02245452,
  0.03907455, 0.0635457, 0.01073519, 0.03157645, 0.02537938, 0.01128226, 
    0.1243276, 0.03561068, 0.03516968, 0.06346747, 0.06160495, 0.05477899, 
    0.07108197, 0.1609621, 0.1259103, 0.1792112, 0.09124856, 0.08013956, 
    0.03917378, 0.01268715, 0.06758113, 0.06956771, 0.09201407, 0.04868809, 
    0.01724927, 0.1491202, 0.1079337, 0.06439862, 0.04970962,
  0.041969, 0.1240745, 0.1483267, 0.1753972, 0.1187934, 0.07363879, 
    0.0815564, 0.1410666, 0.2078423, 0.1426181, 0.1121597, 0.0897717, 
    0.1711739, 0.1922593, 0.1317801, 0.1738341, 0.1443922, 0.1758662, 
    0.1023182, 0.04605149, 0.06902223, 0.0681996, 0.1331585, 0.132629, 
    0.1095566, 0.1059458, 0.09347996, 0.1287097, 0.1171833,
  0.1560866, 0.2087582, 0.117258, 0.115042, 0.1631453, 0.1292314, 0.08287615, 
    0.1304186, 0.2373, 0.2083002, 0.06930799, 0.1646276, 0.07098501, 
    0.1715044, 0.1109281, 0.2160455, 0.2448714, 0.4618749, 0.3342313, 
    0.1433712, 0.09951311, 0.1566317, 0.1938962, 0.3426133, 0.3550428, 
    0.3309868, 0.2208427, 0.1179943, 0.1166633,
  0.3130877, 0.2589948, 0.2914768, 0.1817653, 0.154126, 0.2338575, 0.2743402, 
    0.3620726, 0.3222833, 0.2685822, 0.2210265, 0.200232, 0.1929788, 
    0.2238428, 0.1961997, 0.1116397, 0.3374173, 0.2625462, 0.213199, 
    0.2606885, 0.2187088, 0.1392898, 0.1742877, 0.2545564, 0.1741007, 
    0.1715485, 0.1336705, 0.1623682, 0.2284191,
  0.2319986, 0.2292397, 0.2058535, 0.2203877, 0.2985965, 0.2727433, 
    0.2036923, 0.3491271, 0.315426, 0.3396053, 0.2711369, 0.2702153, 
    0.2197465, 0.1897231, 0.2438767, 0.4681285, 0.4983529, 0.4331554, 
    0.304523, 0.3385501, 0.2831077, 0.2087062, 0.23735, 0.2139591, 0.2119349, 
    0.1846767, 0.1331625, 0.1054729, 0.2702278,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0.002879241, -0.0003239195, 0, 0, 0, 0, 0, 0, 0, 0, 0, -7.300912e-06, 
    0.01724504, 0.2159359, 0.157343, 0.1690706, 0.141106, 0.1478283, 
    0.121247, 0.1457795, 0.111696, 0.1269714, 0.1718466, 0.1809255, 
    0.1979163, 0.1624601, 0.1123992, 0.07845632, 0.0373401,
  0.2300213, 0.3226455, 0.2268556, 0.2215019, 0.04603687, 0.04374039, 
    0.1071022, 0.01695665, 0.004223095, 0.03061308, 0.02168561, 0.04235755, 
    0.280617, 0.2571158, 0.2357538, 0.2228637, 0.2872662, 0.238013, 
    0.3659561, 0.3924099, 0.2904858, 0.2491133, 0.3012855, 0.3825775, 
    0.4158379, 0.2917798, 0.2719601, 0.1373042, 0.1804769,
  0.1693519, 0.2696297, 0.2531583, 0.2138117, 0.3104526, 0.3151239, 
    0.3265559, 0.2242056, 0.2723146, 0.2791231, 0.2453111, 0.3120802, 
    0.2670025, 0.2421027, 0.2461112, 0.2445735, 0.2745892, 0.2913726, 
    0.2343746, 0.2295129, 0.2853838, 0.2677241, 0.3015429, 0.238076, 
    0.2683847, 0.2305217, 0.2060288, 0.1700826, 0.2635792,
  0.1964662, 0.2116597, 0.1777893, 0.1476285, 0.1386017, 0.1704733, 
    0.1861014, 0.2320608, 0.22935, 0.2595539, 0.262674, 0.2582086, 0.2242593, 
    0.1686685, 0.1325984, 0.1139011, 0.08316595, 0.1501696, 0.1693594, 
    0.2288944, 0.232213, 0.1732145, 0.2032009, 0.1601294, 0.07574234, 
    0.1163768, 0.1488007, 0.1917947, 0.1671021,
  0.1060717, 0.08982318, 0.09417126, 0.06757901, 0.07994968, 0.0791931, 
    0.07099467, 0.06089596, 0.04755042, 0.04401501, 0.04982238, 0.0541403, 
    0.05455783, 0.08454934, 0.03761571, 0.05390962, 0.06362439, 0.057275, 
    0.06581725, 0.05243379, 0.09819308, 0.1351668, 0.1421959, 0.1238207, 
    0.05338312, 0.08556957, 0.06359055, 0.1067651, 0.1222454,
  0.005018848, 0.01025969, 0.06379755, 0.06323158, 0.07074347, 0.0223933, 
    0.0007055236, 0.001436562, 0.002509088, -7.759035e-06, 0.02586189, 
    0.04931965, 0.06920525, 0.06339823, 0.06448948, 0.1156813, 0.0867006, 
    0.04681715, 0.1504711, 0.08125404, 0.01288928, 0.02460739, 0.01154312, 
    0.03435006, 0.1316282, 0.1119889, 0.05674338, 0.05002544, 0.04313643,
  1.210653e-07, 0.006872704, 0.09724414, 0.007544121, 0.01606289, 0.06656828, 
    0.0898528, 0.05620059, 6.140357e-07, -7.711395e-06, 0.07495293, 
    0.07840751, 0.003900863, 0.02277626, 0.08222853, 0.08456481, 0.04765242, 
    0.100022, 0.0180026, 1.565665e-07, 2.979743e-08, 1.88505e-08, 
    5.088083e-09, 0.0001553438, 0.03758341, 0.1184665, 0.01310178, 
    4.440135e-05, 1.781878e-07,
  6.140212e-07, 0.02307822, 0.1825557, 0.002648162, 0.001496702, 0.01341987, 
    0.06140136, 0.1151447, 0.007509132, 0.0016027, 0.002511446, 0.006525555, 
    0.1084496, 0.1101588, 0.08037295, 0.03955221, 0.007571153, 0.001436918, 
    3.607071e-05, 8.829079e-08, 1.115728e-07, 1.804605e-07, 0.01090757, 
    0.08510187, 0.04921928, 0.3051488, 0.0001519514, 1.227225e-06, 
    3.481218e-07,
  0.04653901, 0.2706259, 0.1951954, 0.001744208, 0.01363508, 0.06653092, 
    0.1130618, 0.1304377, 0.1359043, 0.1629757, 0.07749352, 0.05448798, 
    0.03127591, 0.02579311, 0.00486951, 0.003199758, 0.0003510004, 
    5.4557e-05, 0.01516441, 0.003695823, 6.475156e-05, 0.01373046, 
    0.04988253, 0.1123146, 0.01832878, 0.002997213, 0.0006395671, 
    0.0007111849, 0.003754857,
  0.1007159, 0.07389325, 0.06165129, 0.1431019, 0.006056599, 0.005823422, 
    0.04870851, 0.05056033, 0.1197102, 0.1168977, 0.03353272, 0.01536636, 
    0.09789418, 0.09212458, 0.1229016, 0.178393, 0.08882578, 0.109312, 
    0.06667153, 0.3221825, 0.1862649, 0.2510948, 0.2153524, 0.0417558, 
    0.05542809, 0.03202169, 0.129025, 0.1324189, 0.1339372,
  0.000130248, 1.233164e-05, 6.464562e-06, 1.629955e-07, 0.0001259983, 
    1.257973e-06, 0.1858815, 0.06318074, 0.1928163, 0.03610903, 0.0878815, 
    0.04139922, 0.09050006, 0.04327277, 0.01067732, 0.01996185, 0.002239885, 
    6.288342e-07, -2.343558e-06, 0.03355438, 0.0534629, 0.118834, 0.01191688, 
    0.06090612, 0.0112554, 0.06890172, 0.08150289, 0.002632764, 0.002024046,
  0.0002064465, 0.01377841, 4.172396e-05, 4.48699e-09, 0.0001485662, 
    -2.167882e-06, 0.0003310602, 0.2027869, 0.2894646, 0.242012, 0.09507195, 
    0.06226747, 0.05926254, 0.06848131, 0.03711219, 0.04517898, 0.01290725, 
    0.003213041, -5.457756e-06, 0.0001473289, 0.08337604, 0.03617523, 
    0.09355164, 0.02271562, 0.03912365, 0.03114942, 0.05023216, 0.005544378, 
    0.02034684,
  0.03422961, 0.02299009, 0.009557024, 0.03846227, 0.02216255, 0.01459255, 
    0.1056156, 0.01735323, 0.02751836, 0.05763623, 0.05662102, 0.05584436, 
    0.08085751, 0.1693822, 0.138666, 0.1914016, 0.1010557, 0.08867727, 
    0.0296911, 0.003570464, 0.05954111, 0.04141494, 0.107991, 0.05698581, 
    0.02420847, 0.1480859, 0.1141912, 0.08986315, 0.05525437,
  0.04408798, 0.1256891, 0.1545091, 0.1848422, 0.08927404, 0.05286636, 
    0.07872818, 0.1602714, 0.2031018, 0.1523148, 0.1114003, 0.0983787, 
    0.2050115, 0.1676211, 0.1385967, 0.1873792, 0.1328287, 0.1621029, 
    0.08898536, 0.04880088, 0.07589434, 0.04989811, 0.1386137, 0.1489034, 
    0.121894, 0.09076133, 0.1009521, 0.122962, 0.1013626,
  0.1586178, 0.2058599, 0.145663, 0.1407643, 0.1825648, 0.1358688, 
    0.09620218, 0.142376, 0.2883313, 0.2001687, 0.07319599, 0.1602888, 
    0.08323014, 0.1750398, 0.1047446, 0.2230737, 0.2330909, 0.4885195, 
    0.3269763, 0.151291, 0.09839188, 0.1965027, 0.2342638, 0.3662543, 
    0.3164641, 0.3188305, 0.2256144, 0.1435514, 0.12925,
  0.3381713, 0.2592607, 0.2786577, 0.2442926, 0.1935148, 0.2345739, 
    0.2915588, 0.3817952, 0.3315016, 0.2397644, 0.2397274, 0.1989303, 
    0.203405, 0.2327629, 0.1914768, 0.1359225, 0.3838313, 0.3015943, 
    0.2062952, 0.2941905, 0.1943306, 0.1451919, 0.1412184, 0.2620125, 
    0.1513377, 0.1883059, 0.1410674, 0.1684287, 0.214525,
  0.1741044, 0.2011874, 0.1720744, 0.2033524, 0.294458, 0.2723018, 0.2818365, 
    0.39946, 0.4011014, 0.3632851, 0.2884207, 0.2942808, 0.2916091, 
    0.1892178, 0.2391098, 0.4164539, 0.4608684, 0.368792, 0.2937279, 
    0.3258539, 0.255594, 0.1839372, 0.2658855, 0.2405192, 0.2450307, 
    0.2067242, 0.156397, 0.1489628, 0.2176956,
  0, 0, 0, 0, 0, 0, 0, -7.144712e-07, -4.722776e-07, -2.30084e-07, 
    1.210968e-08, 2.543033e-07, 4.96497e-07, 7.386906e-07, -0.0002083428, 
    -0.0001621147, -0.0001158866, -6.965856e-05, -2.343049e-05, 2.279758e-05, 
    6.902565e-05, 0.0001522427, 0.0001057725, 5.930221e-05, 1.283195e-05, 
    -3.363832e-05, -8.010858e-05, -0.0001265788, 0,
  0.01253692, 0.00167431, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.813885e-05, 
    0.04286562, 0.2155251, 0.1324699, 0.1654923, 0.1225865, 0.1688684, 
    0.1232484, 0.1418245, 0.168682, 0.2263457, 0.1597975, 0.1708272, 
    0.1867128, 0.1416433, 0.1063737, 0.08004363, 0.1074397,
  0.2395806, 0.3450722, 0.2214209, 0.2262395, 0.08834197, 0.04698767, 
    0.1322894, 0.04260911, 0.006233814, 0.1225831, 0.07718437, 0.09625766, 
    0.2933735, 0.2925886, 0.2632481, 0.3051814, 0.3116001, 0.3805228, 
    0.457235, 0.4129462, 0.3516743, 0.3558234, 0.3492723, 0.400986, 
    0.4094566, 0.2759975, 0.3334994, 0.1525208, 0.2051943,
  0.1784989, 0.2831555, 0.2638564, 0.2259796, 0.3270456, 0.3208339, 0.313117, 
    0.242934, 0.2866544, 0.2844219, 0.2533901, 0.3180889, 0.2466409, 
    0.2437688, 0.2844518, 0.245026, 0.2815048, 0.2936143, 0.3077723, 
    0.2593246, 0.2747003, 0.2659633, 0.3153672, 0.2123243, 0.252977, 
    0.2395755, 0.207032, 0.1682697, 0.2515188,
  0.2097192, 0.2096486, 0.1799424, 0.1466404, 0.1383498, 0.1773994, 
    0.2024539, 0.2491509, 0.2365571, 0.2858737, 0.2812195, 0.2453383, 
    0.209953, 0.1677011, 0.128324, 0.1174648, 0.09220636, 0.1563573, 
    0.1625888, 0.2312951, 0.2243059, 0.1531237, 0.1665522, 0.1660338, 
    0.06908122, 0.1208054, 0.145288, 0.193974, 0.1955206,
  0.1145261, 0.09578026, 0.1068442, 0.08683016, 0.08814767, 0.09445102, 
    0.06748676, 0.07733724, 0.05862094, 0.04642669, 0.05866583, 0.06618656, 
    0.05290611, 0.1004289, 0.03265376, 0.06540987, 0.06540558, 0.06035524, 
    0.06662828, 0.05267287, 0.1092763, 0.1358619, 0.1354381, 0.1310096, 
    0.0445246, 0.08872104, 0.05797332, 0.1187369, 0.133027,
  0.005275201, 0.006254755, 0.04419966, 0.0695923, 0.05962595, 0.03558135, 
    0.006022705, 0.003932469, 0.004815873, 0.000340712, 0.006237211, 
    0.04610872, 0.0912937, 0.07100344, 0.0676, 0.1217072, 0.08494753, 
    0.03570791, 0.1467835, 0.08385383, 0.02765662, 0.03897997, 0.01319565, 
    0.0164669, 0.1367573, 0.1171876, 0.06030906, 0.06238834, 0.05057536,
  7.765693e-08, 0.001646167, 0.1060139, 0.02089883, 0.0210318, 0.07094297, 
    0.1113864, 0.04007217, 0.001431689, -1.91203e-07, 0.05867929, 0.0489581, 
    0.005842662, 0.03855436, 0.06856171, 0.08655292, 0.04908328, 0.1038881, 
    0.04107682, 1.204048e-05, 1.827795e-07, 2.216354e-08, -2.641542e-07, 
    3.030764e-06, 0.0337481, 0.1419633, 0.006043265, -1.376353e-05, 
    1.828891e-06,
  -6.080755e-06, 0.01030388, 0.1477431, 0.02145269, 0.002125268, 0.01336082, 
    0.06610584, 0.1074175, 0.002350935, 0.001365023, 0.00567746, 0.002576188, 
    0.09505797, 0.07096716, 0.07521975, 0.04361446, 0.01073598, 0.00136864, 
    3.336342e-05, 6.693452e-08, 1.051259e-07, 4.267267e-08, 0.004148578, 
    0.05873923, 0.03576814, 0.1828904, 0.0002600798, 3.84308e-07, 3.265055e-07,
  0.009214538, 0.2355791, 0.1222698, 0.001345813, 0.01268761, 0.04351633, 
    0.09988678, 0.09371074, 0.1005557, 0.1365191, 0.06756502, 0.03242073, 
    0.03099966, 0.02779523, 0.006219358, 0.004045546, 0.0002193883, 
    0.0002337701, 0.01115281, 0.003396964, 0.0006101765, 0.01731922, 
    0.05078396, 0.06979703, 0.02228269, 0.001880824, 0.0008309108, 
    0.0005571194, 0.001308645,
  0.05452762, 0.02821242, 0.01622181, 0.1975412, 0.01934278, 0.006147055, 
    0.06514476, 0.0487302, 0.07789966, 0.1053882, 0.02207641, 0.01261299, 
    0.07422579, 0.07625458, 0.1027494, 0.1622431, 0.09162466, 0.1095438, 
    0.05583365, 0.2849815, 0.1783115, 0.2269373, 0.2013983, 0.03529818, 
    0.04580071, 0.02218826, 0.1099526, 0.09206212, 0.09627473,
  1.954976e-06, 8.493222e-06, 3.608719e-06, 4.932404e-08, 9.50637e-06, 
    3.594706e-07, 0.1549345, 0.06113458, 0.1603958, 0.03913136, 0.0904384, 
    0.03633405, 0.06775731, 0.04048005, 0.01147993, 0.01648679, 0.001895122, 
    -4.559918e-05, -1.543361e-05, 0.03782336, 0.0373476, 0.108039, 
    0.01093974, 0.04701958, 0.01140989, 0.06297331, 0.07036683, 0.000194178, 
    0.0002908938,
  4.747969e-05, 0.01022771, 9.348265e-05, 2.691304e-09, 1.424518e-05, 
    1.080182e-06, 0.0001889838, 0.2675394, 0.3393873, 0.2545859, 0.08391098, 
    0.07576253, 0.05618022, 0.05487918, 0.03104736, 0.04154537, 0.007029162, 
    0.01155291, -3.996284e-07, 7.621482e-05, 0.08572294, 0.02893585, 
    0.07480212, 0.019855, 0.03218467, 0.02749417, 0.03345306, 0.006380203, 
    0.01332548,
  0.02526738, 0.006918193, 0.01515817, 0.03954857, 0.01884086, 0.007606782, 
    0.0836525, 0.006598998, 0.0266489, 0.07736807, 0.05059801, 0.06578457, 
    0.08185864, 0.1694742, 0.1262617, 0.1716443, 0.118292, 0.1051567, 
    0.04071981, 0.00131154, 0.05173191, 0.03163724, 0.1015331, 0.05503796, 
    0.02297327, 0.126691, 0.1151784, 0.09888162, 0.07591758,
  0.05066225, 0.1327341, 0.1984349, 0.2273949, 0.08398118, 0.03333135, 
    0.1084021, 0.2011444, 0.201106, 0.1563306, 0.1490471, 0.1644821, 
    0.2232706, 0.1845863, 0.1744764, 0.201253, 0.1475404, 0.1692496, 
    0.09732217, 0.04721391, 0.08951046, 0.03599843, 0.1378962, 0.1785192, 
    0.1196816, 0.0919705, 0.1121847, 0.1444835, 0.0976491,
  0.1688803, 0.2034714, 0.1460609, 0.1453664, 0.1816136, 0.1335846, 
    0.1589832, 0.1661311, 0.2553023, 0.2048919, 0.0976612, 0.2148158, 
    0.1059915, 0.2127776, 0.1237726, 0.2228414, 0.2321671, 0.5138751, 
    0.3622111, 0.1377599, 0.1097045, 0.2252889, 0.2068758, 0.3854846, 
    0.3673304, 0.3238846, 0.2574905, 0.130132, 0.1189703,
  0.2664938, 0.2354956, 0.2924026, 0.2032492, 0.2166965, 0.2663957, 
    0.2761989, 0.3928342, 0.3337713, 0.246931, 0.2404266, 0.204545, 
    0.2400061, 0.2916135, 0.2557797, 0.2194633, 0.4035399, 0.2818385, 
    0.2424405, 0.2368721, 0.1720529, 0.1141714, 0.1654573, 0.2819868, 
    0.1662424, 0.2163276, 0.1517296, 0.1683673, 0.2176358,
  0.1930903, 0.1674086, 0.1271133, 0.1293056, 0.2405423, 0.221526, 0.2378345, 
    0.3812423, 0.4156462, 0.3798506, 0.3194839, 0.3528571, 0.2697366, 
    0.2192446, 0.3090511, 0.4936598, 0.4836201, 0.3449712, 0.2551737, 
    0.2479116, 0.189748, 0.1841148, 0.2866612, 0.3201987, 0.2689294, 
    0.2227865, 0.2147465, 0.1814779, 0.2276051,
  1.881689e-05, 1.200311e-05, 5.189337e-06, -1.624438e-06, -8.438213e-06, 
    -1.525199e-05, -2.206576e-05, -2.510263e-07, 3.309159e-07, 9.128582e-07, 
    1.4948e-06, 2.076743e-06, 2.658685e-06, 3.240627e-06, -0.0007606444, 
    -0.0006729095, -0.0005851747, -0.0004974398, -0.0004097049, 
    -0.0003219701, -0.0002342352, -0.0006430517, -0.0007245548, 
    -0.0008060578, -0.0008875608, -0.0009690639, -0.001050567, -0.00113207, 
    2.426791e-05,
  0.06458889, 0.006456007, -0.0004724902, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.002178364, 0.08264544, 0.1828716, 0.1395119, 0.1566684, 0.1491674, 
    0.1753924, 0.123353, 0.1377833, 0.1717151, 0.2474314, 0.1689497, 
    0.1838993, 0.1849855, 0.1216982, 0.1040326, 0.08683234, 0.1414526,
  0.2308246, 0.3472365, 0.2379127, 0.2247235, 0.1304852, 0.04935478, 
    0.1382663, 0.103708, 0.08894392, 0.1587057, 0.1714399, 0.1554116, 
    0.2840315, 0.3060523, 0.2962831, 0.3385286, 0.3262744, 0.2939912, 
    0.4567688, 0.3963103, 0.3299937, 0.2878598, 0.3606656, 0.475247, 
    0.4241254, 0.2819097, 0.3368025, 0.2153996, 0.2094088,
  0.2645955, 0.3199721, 0.2951519, 0.2236802, 0.3733969, 0.2927482, 
    0.3031642, 0.2640784, 0.2987973, 0.2866072, 0.2596018, 0.2909488, 
    0.2582315, 0.2562748, 0.2759129, 0.2713115, 0.2890924, 0.3138132, 
    0.3037524, 0.2917122, 0.2855539, 0.2754232, 0.3297623, 0.2354544, 
    0.2599328, 0.252969, 0.1960548, 0.2071729, 0.3244258,
  0.2053028, 0.2334382, 0.1862612, 0.1649387, 0.1521444, 0.1693292, 
    0.1954319, 0.2461145, 0.2493477, 0.3058313, 0.2991746, 0.2497645, 
    0.1858754, 0.1814218, 0.1270068, 0.1119953, 0.1013147, 0.1867877, 
    0.1829573, 0.2337554, 0.2473202, 0.181241, 0.1953606, 0.1698796, 
    0.1215353, 0.127255, 0.1362709, 0.1918704, 0.1814768,
  0.1435596, 0.1119919, 0.1143679, 0.08518439, 0.1193141, 0.1123205, 
    0.093812, 0.1065365, 0.07097414, 0.06545332, 0.0702688, 0.07007866, 
    0.05510163, 0.1083781, 0.03212005, 0.07782063, 0.06958123, 0.0653509, 
    0.08294258, 0.0635417, 0.1178013, 0.1536289, 0.1597291, 0.1443402, 
    0.0498003, 0.09276464, 0.05874154, 0.1348089, 0.1501166,
  0.004475353, 0.002122514, 0.04234307, 0.07608689, 0.0477486, 0.03931938, 
    0.02328681, 0.02004981, 0.004865622, 0.003015568, 0.00493482, 0.03655981, 
    0.1226132, 0.08295603, 0.07455985, 0.1324552, 0.08696309, 0.03221821, 
    0.1576927, 0.1212307, 0.05939477, 0.05892808, 0.01398277, 0.001896909, 
    0.09469514, 0.1170405, 0.06833287, 0.07024236, 0.07357133,
  3.85526e-08, 0.0002742452, 0.08806439, 0.01599278, 0.04458886, 0.08016493, 
    0.1114513, 0.0165224, 0.009216798, -1.871278e-08, 0.009697322, 
    0.01373597, 0.01088275, 0.05384635, 0.09762989, 0.07856219, 0.04306648, 
    0.1079947, 0.07431556, 0.002410245, 0.0001622202, 5.354859e-07, 
    7.875754e-09, 7.5686e-05, 0.0282692, 0.1049298, 0.005015702, 1.79965e-05, 
    1.629982e-06,
  3.944275e-08, 0.005929339, 0.09480303, 0.08463229, 0.005957361, 0.01363136, 
    0.06924095, 0.1085813, 0.002276686, 0.002536469, 0.009553755, 
    0.001795267, 0.09241134, 0.05362404, 0.08231146, 0.05204483, 0.02619161, 
    0.004633995, 0.000192491, 1.228313e-07, 9.386208e-08, -1.085293e-07, 
    0.002047574, 0.05802129, 0.02604705, 0.05383526, 0.001365182, 
    1.002883e-07, 1.106924e-07,
  0.000704083, 0.2056083, 0.0409011, 0.001792201, 0.01139895, 0.02677724, 
    0.09102762, 0.07365765, 0.09171543, 0.1330923, 0.05196585, 0.02298017, 
    0.0343543, 0.02728642, 0.01088349, 0.005694422, 0.0007399809, 
    3.31643e-05, 0.003203031, 0.0004488492, 0.001671513, 0.01308821, 
    0.06084348, 0.06058295, 0.03947372, 0.001649184, 0.002525772, 
    7.519848e-05, 0.001058668,
  0.03689109, 0.008630161, 0.006929998, 0.2386353, 0.05022755, 0.01038113, 
    0.07324509, 0.04633695, 0.05762129, 0.09815805, 0.01822149, 0.01248352, 
    0.05963055, 0.06686135, 0.08861616, 0.1504591, 0.1002417, 0.1190341, 
    0.06119424, 0.2564347, 0.1766109, 0.2108888, 0.195868, 0.03327357, 
    0.03690132, 0.02183498, 0.09340198, 0.07231386, 0.06981181,
  3.056425e-07, 5.554623e-06, 2.806919e-06, -4.18041e-08, 8.269382e-07, 
    1.166217e-07, 0.1490252, 0.05842814, 0.1544222, 0.03962632, 0.1101226, 
    0.04017194, 0.05480572, 0.03963278, 0.01737144, 0.02431936, 0.004299693, 
    0.01581621, 0.0001280352, 0.05273106, 0.03532126, 0.1004821, 0.01231412, 
    0.03412277, 0.01098985, 0.05753335, 0.06038988, 4.644693e-05, 4.441129e-05,
  2.562168e-05, 0.001273437, 0.005428072, 1.900196e-09, 5.60178e-06, 
    6.054004e-07, -1.372675e-05, 0.322457, 0.3247666, 0.2559285, 0.08753717, 
    0.09162134, 0.06486147, 0.05205766, 0.02944256, 0.04208884, 0.008273696, 
    0.0241847, 5.105792e-07, -3.939028e-05, 0.0601873, 0.02707546, 
    0.06834345, 0.02035501, 0.02443109, 0.02738006, 0.02712325, 0.008719301, 
    0.009540047,
  0.02421333, 0.002886273, 0.01366677, 0.04589862, 0.01581562, 0.0112792, 
    0.08226355, -1.514858e-06, 0.02345119, 0.09249191, 0.06394278, 0.0727695, 
    0.08446029, 0.1887943, 0.122849, 0.1498621, 0.1270381, 0.1022885, 
    0.05221777, 0.002806892, 0.01926109, 0.02981518, 0.09294212, 0.05753825, 
    0.01784982, 0.1073621, 0.09204388, 0.1209379, 0.07005277,
  0.0673388, 0.1452194, 0.2100895, 0.2266471, 0.09676103, 0.04933025, 
    0.1107088, 0.2049317, 0.2108, 0.1586309, 0.1788278, 0.1879101, 0.2715755, 
    0.2093447, 0.1733078, 0.2067902, 0.1583131, 0.1739943, 0.1108619, 
    0.04430585, 0.1074553, 0.02820655, 0.2034359, 0.2058012, 0.2161929, 
    0.1333214, 0.1385839, 0.1680675, 0.1119931,
  0.1701699, 0.2282966, 0.1855513, 0.1554986, 0.1826952, 0.157186, 0.1617869, 
    0.2035112, 0.3057423, 0.245355, 0.1361721, 0.1997807, 0.1165703, 
    0.2308363, 0.1461058, 0.2754003, 0.2471059, 0.5552813, 0.3574137, 
    0.1407539, 0.1315179, 0.2301517, 0.2503568, 0.4357589, 0.4098007, 
    0.3318672, 0.2408718, 0.1669482, 0.1787304,
  0.2972559, 0.2647394, 0.3153409, 0.2707257, 0.2297638, 0.3092267, 
    0.3335928, 0.4143596, 0.3628206, 0.2433041, 0.2430106, 0.2993877, 
    0.223207, 0.2770613, 0.3969698, 0.2666956, 0.3868344, 0.3167573, 
    0.2237038, 0.2537065, 0.1511809, 0.1152823, 0.1551278, 0.2812304, 
    0.1813314, 0.278423, 0.1598979, 0.1395023, 0.2538512,
  0.2098216, 0.1756084, 0.1403382, 0.181199, 0.2494888, 0.2809871, 0.3673815, 
    0.3748974, 0.4335397, 0.4218578, 0.350632, 0.3720257, 0.321918, 
    0.2280522, 0.2814542, 0.4986335, 0.4163308, 0.2876768, 0.2227663, 
    0.2791504, 0.2553585, 0.2632563, 0.2742097, 0.337112, 0.3594898, 
    0.3716641, 0.242317, 0.1901949, 0.2565775,
  0.003274292, 0.002119844, 0.0009653963, -0.0001890512, -0.001343499, 
    -0.002497946, -0.003652394, 6.239866e-05, 0.0001538454, 0.0002452921, 
    0.0003367388, 0.0004281855, 0.0005196322, 0.0006110789, -0.009336403, 
    -0.006934186, -0.004531968, -0.002129751, 0.0002724653, 0.002674682, 
    0.005076899, -0.002373186, -0.003712402, -0.005051618, -0.006390834, 
    -0.00773005, -0.009069266, -0.01040848, 0.004197849,
  0.09254536, 0.02910665, 0.00754202, -6.21305e-05, 0, 0, 0, 0, 0, 0, 
    0.0003615627, 0.01981817, 0.1078455, 0.1775926, 0.122493, 0.1340488, 
    0.1367945, 0.1826597, 0.1422357, 0.1397798, 0.1868311, 0.2334268, 
    0.1860097, 0.1871131, 0.1740377, 0.1169324, 0.1135694, 0.1108971, 
    0.1599799,
  0.2158216, 0.2913547, 0.2356786, 0.2126013, 0.1585219, 0.04362791, 
    0.1514582, 0.1748794, 0.2165709, 0.1830238, 0.1905113, 0.2108549, 
    0.283823, 0.2914879, 0.3137317, 0.2888122, 0.2756205, 0.2458113, 
    0.419606, 0.3374994, 0.2883413, 0.247428, 0.3569244, 0.4883628, 
    0.3996975, 0.264674, 0.2610977, 0.1751951, 0.2307273,
  0.2285686, 0.3025942, 0.2990495, 0.2564652, 0.3716263, 0.316555, 0.320708, 
    0.2348511, 0.3184263, 0.2989896, 0.2417388, 0.2927278, 0.242241, 
    0.2773626, 0.3112859, 0.2789497, 0.2832662, 0.3153268, 0.3032188, 
    0.2995646, 0.3033907, 0.3087953, 0.3279599, 0.2593919, 0.2563847, 
    0.2361832, 0.2232915, 0.2118084, 0.3036154,
  0.2057221, 0.2534523, 0.2095838, 0.1775636, 0.1707039, 0.1756346, 
    0.2116315, 0.2590421, 0.2517632, 0.3135864, 0.3075303, 0.2377776, 
    0.1750111, 0.1880489, 0.1417697, 0.1322674, 0.1277741, 0.1996563, 
    0.209604, 0.2278873, 0.2523406, 0.1969551, 0.1954782, 0.1773731, 
    0.0783825, 0.1216386, 0.1167762, 0.268588, 0.2033727,
  0.1717891, 0.1383521, 0.1284017, 0.09435835, 0.1255707, 0.1394225, 
    0.1368668, 0.1179579, 0.08434622, 0.09491665, 0.07676934, 0.07610641, 
    0.0747305, 0.09839456, 0.03696916, 0.08252732, 0.08338933, 0.08259612, 
    0.100232, 0.08585281, 0.1455783, 0.1639407, 0.1855928, 0.164991, 
    0.04802285, 0.1069324, 0.07926051, 0.1542624, 0.1724251,
  0.01087605, 0.002656449, 0.04202349, 0.06632491, 0.04523952, 0.04041707, 
    0.02174623, 0.01953201, 0.005411329, 0.009380329, 0.006332407, 
    0.02723333, 0.1480089, 0.08157896, 0.09932051, 0.1464366, 0.08996087, 
    0.04017958, 0.1670359, 0.1448449, 0.0887734, 0.08131809, 0.01579103, 
    -0.0002057162, 0.05801284, 0.1018021, 0.06548605, 0.0821074, 0.08386442,
  2.835139e-08, 0.0004042468, 0.09403612, 0.01157412, 0.05088498, 0.06594823, 
    0.1096429, 0.01112878, 0.01146018, -7.612019e-08, 0.0002009131, 
    0.01415078, 0.02283933, 0.06875311, 0.1028903, 0.07845845, 0.05098813, 
    0.1085307, 0.08319663, 0.02233884, 0.004393475, 0.0007829104, 
    6.679161e-08, 2.323813e-05, 0.01932525, 0.04447034, 0.01448584, 
    0.0001422578, 1.778199e-06,
  1.420764e-07, 0.0009807459, 0.02542648, 0.1182704, 0.008847054, 0.01655754, 
    0.06340256, 0.1110422, 0.006622847, 0.006117783, 0.01206937, 0.00423383, 
    0.09712525, 0.05114887, 0.07888991, 0.04688109, 0.03177203, 0.01309231, 
    0.003945619, 0.0001866769, 3.365431e-07, -3.129477e-07, 0.002447861, 
    0.04691434, 0.0192876, 0.006814715, 0.002791728, 1.367945e-07, 
    4.244277e-08,
  7.597229e-05, 0.2032266, 0.02010459, 0.004962794, 0.01363113, 0.02383872, 
    0.08243006, 0.05842146, 0.09075134, 0.137128, 0.04263777, 0.02124769, 
    0.03440846, 0.02646021, 0.01266638, 0.00839202, 0.002608363, 
    0.0002865313, 9.979042e-05, 2.987136e-05, 0.0004438551, 0.002288558, 
    0.04639129, 0.04934812, 0.06318079, 0.001814345, 0.0051563, 6.845962e-05, 
    0.0001793222,
  0.02625025, 0.005969493, 0.004428575, 0.1548468, 0.0293009, 0.01534393, 
    0.07592242, 0.0424754, 0.04405123, 0.08981372, 0.02140571, 0.01393276, 
    0.05583823, 0.05166487, 0.07212537, 0.1274862, 0.09898897, 0.1173417, 
    0.06607876, 0.2379709, 0.1833422, 0.2028817, 0.2021013, 0.0333221, 
    0.03233134, 0.0226633, 0.07945855, 0.05323965, 0.05504872,
  2.533973e-07, 2.899673e-06, 2.139485e-06, -5.051317e-08, 8.882915e-08, 
    2.060699e-08, 0.1410728, 0.05311765, 0.1654052, 0.04668373, 0.1201828, 
    0.04386986, 0.04890558, 0.0437106, 0.02394256, 0.04449935, 0.01031051, 
    0.01557717, 0.0004829689, 0.0648589, 0.03477394, 0.1030696, 0.01410692, 
    0.02154064, 0.01351545, 0.05473049, 0.05206939, 1.432524e-05, 1.00744e-05,
  6.462125e-06, 0.0001075056, 0.0009711296, 1.175048e-09, 2.090285e-06, 
    3.098833e-07, 0.0001481527, 0.302397, 0.290121, 0.2651804, 0.09547353, 
    0.09807194, 0.07067851, 0.05062357, 0.03195615, 0.03907701, 0.01330459, 
    0.03449395, -1.270115e-07, 0.0003580332, 0.04480544, 0.02442468, 
    0.06591139, 0.02555933, 0.02063405, 0.03274012, 0.0324026, 0.0170249, 
    0.00367667,
  0.02270084, 0.001853457, 0.0165661, 0.05360867, 0.01156181, 0.008071261, 
    0.05680342, 0.003115897, 0.02063361, 0.08395773, 0.07210699, 0.07708133, 
    0.08937556, 0.1885753, 0.1144382, 0.1543598, 0.1407502, 0.09897573, 
    0.07043306, 0.001133104, 0.003427276, 0.02758379, 0.08586263, 0.05898554, 
    0.01943971, 0.08749258, 0.1057261, 0.1042364, 0.05960643,
  0.08481853, 0.1901592, 0.2364886, 0.2256262, 0.102129, 0.07280008, 
    0.09510533, 0.2043249, 0.2321726, 0.1546914, 0.1826188, 0.2693643, 
    0.3005515, 0.2438937, 0.1856579, 0.2354497, 0.1981122, 0.1821466, 
    0.1109281, 0.07351571, 0.1124745, 0.03289549, 0.1898504, 0.2276227, 
    0.2291025, 0.1299901, 0.1455975, 0.1807993, 0.1033819,
  0.1846888, 0.2502785, 0.2009527, 0.1773655, 0.1896457, 0.1587849, 
    0.2028145, 0.2414527, 0.3459432, 0.2375359, 0.1657235, 0.185311, 
    0.1335526, 0.2297729, 0.1395899, 0.2684745, 0.2935428, 0.5391436, 
    0.3227048, 0.1589669, 0.1204512, 0.2409082, 0.2154205, 0.4775305, 
    0.383775, 0.3440833, 0.2334707, 0.1849845, 0.1969954,
  0.3467098, 0.3085787, 0.3790341, 0.2768131, 0.2498471, 0.276935, 0.3067251, 
    0.3873568, 0.3591206, 0.2395986, 0.3045599, 0.2853027, 0.2757893, 
    0.3536921, 0.4141438, 0.3226384, 0.4389507, 0.324093, 0.2198374, 
    0.2776734, 0.1574654, 0.1254102, 0.1433423, 0.2465648, 0.1577603, 
    0.3237815, 0.1491027, 0.1248158, 0.2522926,
  0.2005927, 0.219365, 0.2263264, 0.2274628, 0.370674, 0.4098069, 0.3006405, 
    0.3634925, 0.4750357, 0.4486865, 0.3047551, 0.2881269, 0.2705024, 
    0.1995236, 0.2899322, 0.4944589, 0.4235036, 0.2999022, 0.2917244, 
    0.2962411, 0.2334965, 0.3061413, 0.3309315, 0.3092891, 0.2593108, 
    0.3841872, 0.2302308, 0.1719241, 0.2480672,
  0.04760399, 0.0384461, 0.02928821, 0.02013032, 0.01097243, 0.001814537, 
    -0.007343354, 0.01748797, 0.01870978, 0.01993159, 0.0211534, 0.02237521, 
    0.02359702, 0.02481883, -0.008470987, 0.001669213, 0.01180941, 
    0.02194961, 0.03208981, 0.04223001, 0.05237021, 0.0923899, 0.09018578, 
    0.08798166, 0.08577754, 0.08357343, 0.08136931, 0.07916519, 0.05493031,
  0.1480272, 0.06183461, 0.02397298, 0.002854783, 0, 0, 0, 0, 0, 
    0.0001808498, 0.01120334, 0.04286439, 0.1807737, 0.1881068, 0.1166049, 
    0.1115192, 0.1393848, 0.1739816, 0.1563843, 0.1542251, 0.2261096, 
    0.2436184, 0.1988914, 0.188864, 0.1981452, 0.1134033, 0.1585397, 
    0.1325124, 0.171092,
  0.2325559, 0.2824143, 0.2173999, 0.2109562, 0.1457561, 0.04215206, 
    0.1608085, 0.236827, 0.2617554, 0.1975945, 0.1936402, 0.2441767, 
    0.2981348, 0.2836178, 0.2605701, 0.2746891, 0.2517835, 0.2293489, 
    0.3817393, 0.3564846, 0.2841534, 0.2886358, 0.3368637, 0.4572433, 
    0.397294, 0.2764367, 0.2636944, 0.2015439, 0.2452565,
  0.2476708, 0.3085496, 0.3372994, 0.2998127, 0.3885977, 0.3330815, 
    0.3645098, 0.2566207, 0.3229289, 0.3190264, 0.2368554, 0.2963485, 
    0.2538529, 0.3116088, 0.3464682, 0.2914518, 0.3165227, 0.3120387, 
    0.3303593, 0.2988064, 0.3171394, 0.2927418, 0.3367928, 0.2280772, 
    0.2666835, 0.2681939, 0.234739, 0.2961385, 0.2994457,
  0.2548106, 0.294919, 0.2414525, 0.1930133, 0.1770818, 0.1853941, 0.259602, 
    0.2907596, 0.2814056, 0.3224827, 0.3256211, 0.2468143, 0.1906836, 
    0.2147581, 0.1769274, 0.183095, 0.1698067, 0.2153079, 0.2288299, 
    0.2351305, 0.2486933, 0.2119344, 0.2008342, 0.1894964, 0.05423135, 
    0.1318205, 0.1155037, 0.2237399, 0.2230784,
  0.1995978, 0.1652652, 0.138533, 0.1241071, 0.1325745, 0.1453712, 0.1472119, 
    0.1347249, 0.1311977, 0.1384975, 0.1134388, 0.0947518, 0.07261083, 
    0.09277882, 0.05388385, 0.0882407, 0.1113178, 0.09655837, 0.1332333, 
    0.1223253, 0.158228, 0.1865437, 0.1957243, 0.1722509, 0.0416465, 
    0.1226438, 0.1029893, 0.1818806, 0.1918114,
  0.01914886, 0.002171158, 0.03677853, 0.05883022, 0.04437889, 0.05648137, 
    0.03394082, 0.02140941, 0.01080222, 0.05150461, 0.008408562, 0.02509735, 
    0.1038559, 0.1054957, 0.111572, 0.1497493, 0.104848, 0.07279217, 
    0.1965611, 0.1453607, 0.09024201, 0.09367757, 0.04268962, -0.0001327384, 
    0.04108344, 0.1030926, 0.08468298, 0.08781823, 0.08942099,
  7.432766e-09, 0.0007350477, 0.04837338, 0.005067809, 0.04590602, 
    0.07764914, 0.1166441, 0.01793618, 0.006596928, 6.454154e-07, 
    5.634722e-06, 0.001630959, 0.02462893, 0.05957936, 0.1030621, 0.0712061, 
    0.05187484, 0.1173881, 0.07438926, 0.03418149, 0.0111819, 0.003672404, 
    2.752746e-05, 1.827854e-05, 0.00968373, 0.01982248, 0.0421553, 
    0.006156664, 7.514836e-05,
  8.467568e-08, 0.0006897033, 0.005126482, 0.06899022, 0.01196739, 
    0.02960717, 0.06380421, 0.1175502, 0.01122572, 0.01312754, 0.01188424, 
    0.007854809, 0.08982473, 0.05295797, 0.06725888, 0.03891253, 0.02887001, 
    0.01662705, 0.01246623, 0.01255648, 0.0001905386, 5.842135e-07, 
    0.0008457069, 0.03905793, 0.01742298, 0.0003683548, 0.01372922, 
    2.047111e-06, 3.468323e-07,
  0.0002234525, 0.1993681, 0.0180751, 0.008372244, 0.01745412, 0.02227658, 
    0.07139232, 0.04958579, 0.08718983, 0.1540395, 0.03943275, 0.02024404, 
    0.02625587, 0.0245163, 0.01304547, 0.008270011, 0.01503301, 0.0014407, 
    0.0004222224, 2.221137e-05, 0.001607078, 0.002480519, 0.03396768, 
    0.04455376, 0.0498112, 0.00192205, 0.007793515, 0.0005415576, 0.0001240364,
  0.01939857, 0.004926473, 0.004044123, 0.07503814, 0.00393578, 0.01203687, 
    0.0746133, 0.03840856, 0.03239335, 0.07006945, 0.03733127, 0.01638916, 
    0.04815825, 0.03984756, 0.06086749, 0.1081276, 0.09039703, 0.1162668, 
    0.07712353, 0.2326141, 0.2005498, 0.179549, 0.2016036, 0.03641515, 
    0.02681739, 0.02405757, 0.06922525, 0.04530782, 0.04246497,
  1.7218e-07, 1.541827e-06, 1.210134e-06, -2.276899e-08, 1.549267e-08, 
    2.384362e-09, 0.1190253, 0.04452604, 0.1736414, 0.05269988, 0.1125274, 
    0.03906823, 0.04213677, 0.03947394, 0.02326392, 0.04098186, 0.03109599, 
    0.01422521, 0.003711522, 0.07266649, 0.03680684, 0.1030699, 0.01465821, 
    0.0153654, 0.01476299, 0.06225686, 0.0359546, 1.04358e-05, 1.431444e-06,
  2.23441e-06, 3.895208e-05, 0.0007205262, 5.500183e-10, 1.129138e-06, 
    1.362214e-07, 4.136655e-05, 0.2579726, 0.2611925, 0.2477876, 0.08900046, 
    0.1007533, 0.07316906, 0.05422028, 0.04141665, 0.03554617, 0.03223103, 
    0.05573934, 4.802911e-06, 0.001003216, 0.03198287, 0.02619693, 
    0.06249887, 0.03152737, 0.02287201, 0.04148192, 0.03904456, 0.0232982, 
    0.0009735663,
  0.013299, 0.001298118, 0.01844616, 0.06646778, 0.003542867, 0.003205083, 
    0.05096491, 0.0005957047, 0.01576404, 0.07486808, 0.0850297, 0.07914267, 
    0.08470516, 0.1810861, 0.1222928, 0.1802727, 0.1732178, 0.1165515, 
    0.06307423, 0.001504751, 0.0003807165, 0.02558978, 0.09627791, 
    0.05972021, 0.0233615, 0.08472378, 0.104554, 0.09648342, 0.0514553,
  0.07838269, 0.2139304, 0.224357, 0.223774, 0.09185408, 0.07189862, 
    0.08793336, 0.197644, 0.2009118, 0.165613, 0.2138381, 0.2945094, 
    0.2749552, 0.2802216, 0.1974435, 0.254233, 0.245222, 0.1892915, 
    0.1291491, 0.09626476, 0.1051624, 0.0747683, 0.1775947, 0.2914348, 
    0.1750496, 0.1361499, 0.1590153, 0.1843403, 0.1126385,
  0.2018494, 0.235684, 0.2259217, 0.1920533, 0.1942113, 0.1750412, 0.2313403, 
    0.2230912, 0.2947413, 0.2832225, 0.1548387, 0.1548763, 0.1887907, 
    0.2510113, 0.1366943, 0.3011342, 0.320114, 0.5561434, 0.3368748, 
    0.178807, 0.1185176, 0.2156153, 0.1956985, 0.4666463, 0.3571479, 
    0.3199689, 0.233315, 0.2105171, 0.227107,
  0.3618889, 0.3771907, 0.3396994, 0.2394722, 0.207838, 0.2516091, 0.2907103, 
    0.3819202, 0.3240957, 0.2116119, 0.3049265, 0.2703179, 0.3076477, 
    0.3561115, 0.2479201, 0.3051613, 0.3839513, 0.3307984, 0.2255608, 
    0.2435296, 0.1717642, 0.1271739, 0.1626002, 0.2174001, 0.1512978, 
    0.3305152, 0.1392969, 0.1019487, 0.2081136,
  0.153692, 0.2054917, 0.1865329, 0.2208741, 0.3631143, 0.291803, 0.290752, 
    0.3440196, 0.4308862, 0.4095785, 0.2695275, 0.2393785, 0.2782218, 
    0.2448097, 0.2429, 0.3937565, 0.4014151, 0.3005208, 0.2667642, 0.2288994, 
    0.2252803, 0.2713549, 0.3498125, 0.2642569, 0.2354292, 0.3516682, 
    0.2279113, 0.1866647, 0.1931442,
  0.168439, 0.1551169, 0.1417949, 0.1284729, 0.1151509, 0.1018289, 
    0.08850683, 0.08526802, 0.08886553, 0.09246305, 0.09606057, 0.09965809, 
    0.1032556, 0.1068531, 0.1091515, 0.1209332, 0.1327148, 0.1444965, 
    0.1562782, 0.1680599, 0.1798415, 0.2215892, 0.2195321, 0.2174749, 
    0.2154177, 0.2133605, 0.2113034, 0.2092462, 0.1790966,
  0.1690663, 0.07180968, 0.065359, 0.03228244, -0.0007493389, 0, 0, 0, 0, 
    0.0002819458, 0.01513186, 0.09801385, 0.2850856, 0.189435, 0.1235034, 
    0.1086576, 0.203754, 0.1609049, 0.1519791, 0.1493893, 0.2880416, 
    0.2791908, 0.2115528, 0.1865474, 0.2145068, 0.1320101, 0.1848413, 
    0.1521784, 0.1718476,
  0.2419821, 0.2907658, 0.2456693, 0.2040157, 0.1329415, 0.03081864, 
    0.1610828, 0.290659, 0.2648373, 0.2108013, 0.1961924, 0.2351837, 
    0.2978434, 0.2778541, 0.2483404, 0.2384624, 0.257012, 0.2499814, 
    0.3758621, 0.3952697, 0.3001734, 0.316611, 0.343278, 0.44734, 0.4147949, 
    0.3068391, 0.3296586, 0.2851917, 0.2240019,
  0.3124943, 0.2735536, 0.3454358, 0.3505038, 0.3990529, 0.3549211, 0.384367, 
    0.324941, 0.3672841, 0.3440609, 0.2877775, 0.3234819, 0.2701925, 
    0.3343755, 0.3349428, 0.3181046, 0.3605607, 0.3637725, 0.3497939, 
    0.3018619, 0.3106331, 0.2909634, 0.369585, 0.2819537, 0.2988731, 
    0.3030252, 0.2733829, 0.2626783, 0.3675939,
  0.2969065, 0.3168992, 0.2738252, 0.2410129, 0.2025812, 0.2167532, 
    0.2692487, 0.3094641, 0.2867126, 0.3085198, 0.3200937, 0.2727724, 
    0.2018381, 0.2874015, 0.2211575, 0.2691588, 0.2626441, 0.3091331, 
    0.2629662, 0.253162, 0.2626786, 0.2489642, 0.2495154, 0.2089161, 
    0.0732142, 0.1307629, 0.145019, 0.2375938, 0.2592278,
  0.2067535, 0.1917562, 0.1470042, 0.1986943, 0.1503295, 0.1346634, 
    0.1371427, 0.1716817, 0.1724074, 0.1958331, 0.1238896, 0.1003432, 
    0.04978362, 0.1279077, 0.07458434, 0.1024712, 0.1565709, 0.1306228, 
    0.2104878, 0.1890382, 0.1817177, 0.2069893, 0.2209209, 0.1886277, 
    0.04319802, 0.1428253, 0.1429559, 0.2218267, 0.2427838,
  0.0374317, 0.02521102, 0.03262018, 0.06751519, 0.0815286, 0.07534127, 
    0.06302572, 0.0603027, 0.04810065, 0.08304907, 0.00626318, 0.01783119, 
    0.06597101, 0.1129908, 0.1351249, 0.1545765, 0.1667041, 0.1278573, 
    0.2281357, 0.1938236, 0.1336467, 0.1259759, 0.06398652, -0.0001078892, 
    0.02668968, 0.1303736, 0.1200361, 0.09857266, 0.1207235,
  -1.553534e-07, 0.0005693274, 0.02777978, 0.003599372, 0.04208982, 
    0.08962964, 0.1187767, 0.0232866, 0.0441404, -6.030346e-07, 2.684607e-07, 
    0.0001649452, 0.02792979, 0.05202874, 0.1144651, 0.08029963, 0.07667757, 
    0.1292669, 0.06797858, 0.0463852, 0.07983482, 0.03268262, 0.0009908694, 
    1.12147e-05, 0.003172186, 0.009032872, 0.05185485, 0.04390889, 0.001118577,
  9.707306e-07, -4.800974e-05, 0.001000872, 0.04762486, 0.01259564, 
    0.03572249, 0.06964216, 0.106753, 0.01399366, 0.01418429, 0.01379822, 
    0.009561697, 0.1048208, 0.07145229, 0.05391382, 0.03373715, 0.0254269, 
    0.02460242, 0.01589052, 0.0327673, 0.01316618, 0.0001119184, 
    2.773644e-07, 0.03927087, 0.01775221, 7.149817e-05, 0.04009468, 
    0.0005643493, 1.895056e-06,
  0.001818206, 0.2013227, 0.01845333, 0.01227201, 0.01877677, 0.02119455, 
    0.05776182, 0.03905431, 0.08660243, 0.1715401, 0.0380777, 0.01826031, 
    0.02374376, 0.02037332, 0.01464445, 0.009978632, 0.02249595, 0.00633235, 
    0.004757712, 0.002447079, 0.002743443, 0.001925169, 0.01979578, 
    0.04521783, 0.03642922, 0.002326549, 0.01564391, 0.003746036, 0.0001225821,
  0.01478851, 0.004326897, 0.002917636, 0.03966627, 0.0005935505, 0.0136255, 
    0.07042374, 0.03136783, 0.02368794, 0.04925877, 0.05800623, 0.01835474, 
    0.03987693, 0.03035489, 0.0491964, 0.08835871, 0.08892059, 0.1133367, 
    0.07622235, 0.22442, 0.2013891, 0.1570031, 0.196072, 0.0408511, 
    0.02440078, 0.02432158, 0.06207423, 0.0441953, 0.04181219,
  1.288124e-07, 6.922699e-07, 4.483562e-07, -5.418802e-09, 6.303611e-09, 
    -1.622617e-08, 0.09729789, 0.03608936, 0.1881253, 0.04795933, 0.1034953, 
    0.03220234, 0.03542895, 0.03814682, 0.0240964, 0.03149816, 0.04576248, 
    0.05710739, 0.01130207, 0.07407695, 0.04548073, 0.1077246, 0.01624851, 
    0.01318632, 0.01586846, 0.06155697, 0.02538042, 9.866289e-06, 1.98815e-08,
  1.108501e-06, -4.477517e-06, 6.443382e-06, 1.608346e-10, 7.339601e-07, 
    5.664047e-08, 0.0001016506, 0.2109637, 0.2815055, 0.2214911, 0.08539111, 
    0.09805126, 0.07297069, 0.05249811, 0.05536371, 0.0433682, 0.04327901, 
    0.07383613, 0.001108798, 0.002452693, 0.03368712, 0.02635208, 0.06226871, 
    0.03559129, 0.03603835, 0.04420422, 0.05652852, 0.03385366, 0.0001736789,
  0.01011476, 0.001020489, 0.01266422, 0.07819085, 0.001377953, 0.0002748314, 
    0.04883566, 4.119029e-06, 0.008778019, 0.06932441, 0.07925606, 
    0.08021738, 0.0717844, 0.1808198, 0.1624839, 0.1879454, 0.219438, 
    0.1310943, 0.07594141, 0.001100287, 0.0002322217, 0.02424357, 0.1009397, 
    0.08807231, 0.04784462, 0.09247706, 0.1189811, 0.08986554, 0.04717814,
  0.07874564, 0.1730242, 0.2503404, 0.2558872, 0.07156099, 0.08298437, 
    0.08110572, 0.2343537, 0.1952522, 0.1631291, 0.2151496, 0.2439531, 
    0.2718251, 0.3257542, 0.2375001, 0.2869173, 0.280531, 0.1842321, 
    0.1552341, 0.09894724, 0.09104109, 0.06627966, 0.1771913, 0.3591463, 
    0.1808711, 0.1661868, 0.172664, 0.1916181, 0.139952,
  0.2058565, 0.2168407, 0.2089598, 0.1865685, 0.1598746, 0.1743498, 
    0.2017853, 0.2147407, 0.2623688, 0.2674785, 0.1830587, 0.2121635, 
    0.2373992, 0.2093977, 0.1408675, 0.3246342, 0.3657713, 0.5648173, 
    0.3437022, 0.1691454, 0.1479559, 0.3009647, 0.2172167, 0.5413055, 
    0.3964413, 0.2811773, 0.2892693, 0.2635258, 0.2097064,
  0.4185604, 0.4190503, 0.3166989, 0.2399761, 0.2109489, 0.2286765, 
    0.3494759, 0.4074616, 0.3248242, 0.2199201, 0.3323262, 0.3626423, 
    0.2796801, 0.434163, 0.2553368, 0.2623329, 0.3934495, 0.3718551, 
    0.2045092, 0.2568564, 0.1959185, 0.2066463, 0.2520169, 0.2490148, 
    0.155231, 0.2958528, 0.1697571, 0.09119616, 0.2481228,
  0.145045, 0.1762595, 0.1280334, 0.201316, 0.3059506, 0.2441619, 0.306978, 
    0.3700284, 0.3848647, 0.3543828, 0.3177693, 0.2689982, 0.3848859, 
    0.3631054, 0.2707094, 0.3661171, 0.3313846, 0.270693, 0.3257809, 
    0.2833256, 0.159777, 0.2171689, 0.3486421, 0.309314, 0.2793906, 
    0.3499553, 0.2589789, 0.1774278, 0.1699811,
  0.2528341, 0.2436806, 0.2345271, 0.2253736, 0.2162201, 0.2070666, 
    0.1979131, 0.2108992, 0.2170321, 0.2231649, 0.2292978, 0.2354306, 
    0.2415635, 0.2476963, 0.2258062, 0.2285735, 0.2313408, 0.2341081, 
    0.2368755, 0.2396428, 0.2424101, 0.2449083, 0.2451616, 0.2454149, 
    0.2456683, 0.2459216, 0.2461749, 0.2464283, 0.2601569,
  0.1832339, 0.08408518, 0.094083, 0.03996529, 0.006547013, -0.0001371469, 0, 
    0, 0, 0.005602987, 0.01162574, 0.1849934, 0.3216917, 0.1814503, 
    0.1328634, 0.1358276, 0.2159156, 0.1634022, 0.1553188, 0.1446955, 
    0.2767054, 0.2921492, 0.2200567, 0.1779057, 0.2131184, 0.153016, 
    0.1870897, 0.1705836, 0.1792089,
  0.2570284, 0.2811323, 0.2372062, 0.1762137, 0.1185899, 0.02549384, 
    0.144899, 0.311111, 0.2503561, 0.2113459, 0.1934141, 0.2175423, 
    0.2979075, 0.2613088, 0.2672699, 0.2309887, 0.2419327, 0.267514, 
    0.3873203, 0.4634648, 0.294029, 0.3693324, 0.3557245, 0.4781892, 
    0.4130175, 0.321301, 0.3507846, 0.2706307, 0.263888,
  0.3178132, 0.269055, 0.3769247, 0.4434163, 0.4615095, 0.389628, 0.3634394, 
    0.3695267, 0.4875119, 0.3589599, 0.3461245, 0.3567992, 0.2898772, 
    0.3647678, 0.3463797, 0.3555446, 0.3642245, 0.4405613, 0.3796253, 
    0.2845372, 0.3310559, 0.3162392, 0.414071, 0.3870936, 0.312959, 0.329576, 
    0.2923401, 0.241335, 0.3729333,
  0.3341479, 0.3029608, 0.3256746, 0.2580238, 0.2173229, 0.2209643, 
    0.2807581, 0.3055721, 0.3075345, 0.2831911, 0.2597538, 0.2619957, 
    0.1882978, 0.2778442, 0.2067958, 0.2722846, 0.2430182, 0.3098261, 
    0.3099661, 0.2770517, 0.3004535, 0.2812063, 0.2761658, 0.2171776, 
    0.07863988, 0.2076572, 0.2620828, 0.3661928, 0.3110879,
  0.2740124, 0.2532298, 0.1737745, 0.2269028, 0.1963517, 0.1623026, 
    0.1653499, 0.2451834, 0.2295704, 0.1864337, 0.17436, 0.1033052, 
    0.04612692, 0.2027778, 0.1089687, 0.1791051, 0.148396, 0.2262826, 
    0.3193461, 0.2067683, 0.1942019, 0.2046676, 0.2651033, 0.2210629, 
    0.05468944, 0.1677531, 0.2019248, 0.2640182, 0.3257911,
  0.06116373, 0.02197616, 0.03229536, 0.0769218, 0.09648116, 0.1035736, 
    0.08300464, 0.1428993, 0.1309287, 0.09925922, 0.005549384, 0.0123708, 
    0.05662362, 0.09221401, 0.1706797, 0.187505, 0.2101805, 0.1196847, 
    0.2342748, 0.2797151, 0.2498715, 0.1623686, 0.1465617, -4.715317e-05, 
    0.04446096, 0.2062292, 0.2018831, 0.1244197, 0.1708727,
  8.670743e-05, 0.0004127407, 0.01722501, 0.007196205, 0.0461513, 0.09232894, 
    0.1491853, 0.06699505, 0.1615923, 9.4387e-05, 2.029134e-07, 1.071744e-05, 
    0.04478271, 0.07019481, 0.1197466, 0.08595002, 0.08750366, 0.1385753, 
    0.06294281, 0.05954615, 0.3101519, 0.2238784, 0.07201798, 1.612477e-06, 
    0.00129584, 0.009885923, 0.05152031, 0.08924013, 0.03227369,
  1.702194e-05, -3.751926e-05, 0.000189055, 0.02790756, 0.01863524, 
    0.03961988, 0.07816272, 0.09431256, 0.02017561, 0.01601163, 0.01497773, 
    0.01642009, 0.1173011, 0.08204351, 0.0442396, 0.0349786, 0.02696722, 
    0.02827291, 0.01769206, 0.03435958, 0.1162038, 0.009685579, 1.943447e-05, 
    0.04584625, 0.01776779, 2.009694e-05, 0.06548297, 0.03051655, 0.001405758,
  0.02576568, 0.1965558, 0.01761763, 0.01059883, 0.02202982, 0.02371144, 
    0.04712041, 0.03486039, 0.09186225, 0.1978179, 0.04206828, 0.01840756, 
    0.02377873, 0.02237326, 0.01824185, 0.01534889, 0.02373962, 0.01445814, 
    0.02064179, 0.02650354, 0.002653519, 0.001656523, 0.009103539, 
    0.04454344, 0.02826722, 0.007999764, 0.0221495, 0.02063324, 0.0005889567,
  0.01266261, 0.003418153, 0.001586425, 0.02045499, 0.0002339821, 0.01829815, 
    0.06315036, 0.02863159, 0.02088031, 0.03642228, 0.06353477, 0.02213084, 
    0.03739423, 0.02641035, 0.04275184, 0.07251145, 0.07644781, 0.09312078, 
    0.07008618, 0.2056711, 0.183753, 0.1235752, 0.2069106, 0.03905967, 
    0.02611516, 0.02858629, 0.05680696, 0.0411203, 0.03335042,
  1.041696e-07, 2.968386e-07, 1.295938e-07, 6.151045e-10, 5.402406e-09, 
    -2.612995e-06, 0.07660361, 0.02753731, 0.1832884, 0.06211316, 0.1038714, 
    0.03543806, 0.03483189, 0.03942769, 0.02875839, 0.03115383, 0.04933734, 
    0.08336743, 0.04240033, 0.08005788, 0.05210986, 0.1174758, 0.02163786, 
    0.01533535, 0.02028516, 0.059118, 0.03039539, 1.60686e-05, 2.403154e-07,
  7.631235e-07, 7.775297e-06, 0.0009529373, 3.514803e-11, 5.145498e-07, 
    2.693782e-08, 3.454099e-05, 0.1828419, 0.2911284, 0.2005561, 0.1167057, 
    0.1032863, 0.07941151, 0.04721371, 0.05914898, 0.05475065, 0.06108089, 
    0.1219199, 0.01292907, 0.002518994, 0.03528833, 0.0234605, 0.06734651, 
    0.03704035, 0.03909936, 0.05032966, 0.05099263, 0.06820121, 0.0001060107,
  0.009216929, 0.0003697681, 0.009162788, 0.09528202, 0.0006607551, 
    -7.46986e-05, 0.04569716, 2.155145e-06, 0.003020292, 0.06328394, 
    0.08378661, 0.0726187, 0.08980304, 0.2397034, 0.2671193, 0.2477374, 
    0.2624855, 0.1741941, 0.159159, -0.000179652, -3.364317e-05, 0.02983191, 
    0.1160085, 0.1047131, 0.07904858, 0.1022464, 0.1583029, 0.1356272, 
    0.04834496,
  0.08869094, 0.2023275, 0.250641, 0.2497747, 0.06175708, 0.02763431, 
    0.06091851, 0.2384017, 0.1969602, 0.1242742, 0.170284, 0.2443006, 
    0.300171, 0.3347974, 0.3069654, 0.3664362, 0.3163739, 0.1973024, 
    0.1544943, 0.08471894, 0.07770175, 0.03133981, 0.1520887, 0.3164123, 
    0.1815752, 0.1926577, 0.209445, 0.2648799, 0.1514714,
  0.2444248, 0.2264953, 0.2176727, 0.2346978, 0.2005261, 0.2117752, 
    0.1889502, 0.2793017, 0.2502663, 0.2576169, 0.2269501, 0.3547694, 
    0.2690751, 0.2289221, 0.1597472, 0.3832139, 0.376735, 0.575581, 
    0.3334387, 0.1608603, 0.1684757, 0.3358919, 0.2295504, 0.6499085, 
    0.4149858, 0.2739548, 0.3441159, 0.3454405, 0.1803521,
  0.5043468, 0.389745, 0.39897, 0.2976933, 0.2784125, 0.3048976, 0.4735112, 
    0.4755219, 0.3607318, 0.2682201, 0.4378114, 0.3956654, 0.3283758, 
    0.3981073, 0.3538418, 0.2957608, 0.487612, 0.3706796, 0.2486717, 
    0.2837475, 0.2326561, 0.2984814, 0.2878584, 0.2472215, 0.1878243, 
    0.2671496, 0.1955283, 0.1027283, 0.4112554,
  0.1666558, 0.2520927, 0.1865018, 0.236167, 0.34039, 0.2513413, 0.3042689, 
    0.3531586, 0.5310314, 0.4070089, 0.3690237, 0.3917794, 0.420328, 
    0.3183241, 0.3747247, 0.3766647, 0.4180177, 0.3073205, 0.3571335, 
    0.3006168, 0.1791984, 0.2389672, 0.310941, 0.3533893, 0.2746581, 
    0.3332202, 0.2564327, 0.1959237, 0.2065823,
  0.286597, 0.2815888, 0.2765807, 0.2715725, 0.2665644, 0.2615562, 0.256548, 
    0.2494678, 0.2556319, 0.261796, 0.2679601, 0.2741242, 0.2802883, 
    0.2864524, 0.2893362, 0.2875132, 0.2856902, 0.2838672, 0.2820441, 
    0.2802211, 0.2783981, 0.2563358, 0.2570029, 0.25767, 0.2583371, 
    0.2590042, 0.2596713, 0.2603384, 0.2906035,
  0.1986619, 0.09331097, 0.1118456, 0.04670848, 0.02364247, -0.0006968578, 0, 
    0, 0, 0.005163176, 0.04171941, 0.2179785, 0.3253735, 0.1693243, 
    0.1600355, 0.183837, 0.2404745, 0.1649902, 0.1544997, 0.1619826, 
    0.3151487, 0.2939481, 0.2259762, 0.1644027, 0.2011361, 0.1633788, 
    0.2027403, 0.1823552, 0.1970029,
  0.2485283, 0.2989091, 0.227232, 0.1573128, 0.1101831, 0.02856841, 
    0.1425408, 0.3223748, 0.253975, 0.2088952, 0.1878763, 0.1639931, 
    0.2738549, 0.232113, 0.2630911, 0.3006701, 0.29063, 0.2830798, 0.4030829, 
    0.449815, 0.3487695, 0.4210643, 0.3505993, 0.5156354, 0.422733, 
    0.3422414, 0.3191683, 0.300047, 0.2386524,
  0.3128454, 0.4005204, 0.4966882, 0.486454, 0.5153636, 0.4196726, 0.3341326, 
    0.4091051, 0.5412025, 0.2951792, 0.2800488, 0.3662501, 0.3993287, 
    0.3893469, 0.3064011, 0.3667209, 0.389646, 0.4707678, 0.345899, 
    0.2476321, 0.3148177, 0.314314, 0.4180075, 0.3435736, 0.321411, 
    0.3303759, 0.274871, 0.2710045, 0.3022003,
  0.2844145, 0.3123337, 0.3130752, 0.2565167, 0.304167, 0.2746278, 0.2876338, 
    0.268588, 0.2946979, 0.2836677, 0.2652255, 0.2862679, 0.1891212, 
    0.2655587, 0.1791341, 0.222738, 0.2266901, 0.2928766, 0.2862906, 
    0.3171296, 0.3321454, 0.2937146, 0.3091088, 0.2431459, 0.08158484, 
    0.2899283, 0.4173689, 0.4715911, 0.3281311,
  0.3056507, 0.2450837, 0.2142111, 0.285653, 0.2593153, 0.2495791, 0.2298049, 
    0.2838859, 0.2031751, 0.1427286, 0.1117525, 0.1048734, 0.0376224, 
    0.2359221, 0.1266528, 0.2058145, 0.1686417, 0.2465103, 0.2339809, 
    0.1490015, 0.1716107, 0.1775699, 0.2457042, 0.2585181, 0.06532826, 
    0.1776676, 0.2192134, 0.2971569, 0.3030227,
  0.1406692, 0.03796906, 0.02948132, 0.1014139, 0.08451113, 0.2134331, 
    0.1612069, 0.2444552, 0.2536285, 0.07526427, 0.01141729, 0.007067616, 
    0.05353574, 0.09119117, 0.2045957, 0.2887059, 0.1532123, 0.09771959, 
    0.2599969, 0.26592, 0.200035, 0.2981894, 0.2181576, 2.290693e-05, 
    0.06703585, 0.2054622, 0.2958505, 0.2207734, 0.2250346,
  0.03921085, 0.0001454246, 0.01688976, 0.01840744, 0.06257342, 0.09594147, 
    0.1796386, 0.1020219, 0.1568587, 0.007810248, 4.736279e-08, 3.015996e-06, 
    0.08606521, 0.08771734, 0.1307806, 0.09987826, 0.1028269, 0.162494, 
    0.06857974, 0.1109036, 0.3467929, 0.5617676, 0.334067, -5.833771e-06, 
    0.01215475, 0.02978206, 0.05905769, 0.1137239, 0.2665698,
  0.002680098, 0.002414498, 6.706479e-05, 0.01691344, 0.0362254, 0.08668865, 
    0.08561113, 0.08947279, 0.03302896, 0.0330889, 0.02149019, 0.0449292, 
    0.1179284, 0.09217767, 0.03988917, 0.04942753, 0.03653128, 0.04737538, 
    0.04111299, 0.05310842, 0.2290999, 0.1376853, 0.001860849, 0.03617586, 
    0.01252192, 8.032015e-06, 0.09851056, 0.2054474, 0.02931823,
  0.1187385, 0.1867892, 0.01216975, 0.01359704, 0.03497053, 0.03177006, 
    0.04752242, 0.03549436, 0.09338236, 0.183069, 0.04697959, 0.02508069, 
    0.02918598, 0.05601645, 0.03176508, 0.07017832, 0.04042305, 0.01423408, 
    0.03084357, 0.04866917, 0.03352863, 0.005089432, 0.002950165, 0.0299516, 
    0.01303578, 0.02891584, 0.05858452, 0.04673996, 0.01589236,
  0.009785493, 0.001770837, 0.0009771845, 0.007862726, 9.785386e-05, 
    0.02882595, 0.05848643, 0.0369122, 0.01639627, 0.03280538, 0.0374454, 
    0.02854818, 0.05097434, 0.03242182, 0.04205944, 0.06306273, 0.08310117, 
    0.0824755, 0.08801842, 0.1711758, 0.1450877, 0.1152738, 0.1787068, 
    0.03270809, 0.0607397, 0.04050774, 0.0558232, 0.04347908, 0.02388541,
  8.919248e-08, 1.679467e-07, 4.122267e-08, 1.597899e-10, 5.0405e-09, 
    -0.0001232343, 0.05607014, 0.02375166, 0.1512674, 0.05533104, 0.09806286, 
    0.03556792, 0.04067441, 0.04715648, 0.03789807, 0.04062301, 0.06690764, 
    0.1066544, 0.2012383, 0.1164545, 0.06027089, 0.1278899, 0.03281023, 
    0.02244342, 0.03204956, 0.06842459, 0.05470948, 0.0001395607, 2.252796e-07,
  5.986172e-07, -9.518346e-05, 0.002481705, 6.663428e-12, 3.901818e-07, 
    1.651856e-08, 1.975794e-05, 0.1857036, 0.313799, 0.2037502, 0.1594985, 
    0.06552906, 0.0866584, 0.05713813, 0.06614368, 0.08313935, 0.1053353, 
    0.1609611, 0.1196895, 0.001977263, 0.02427771, 0.02420915, 0.06678801, 
    0.04423803, 0.05164596, 0.04886905, 0.05216893, 0.1121317, 0.0009581975,
  0.00956688, 0.0007775179, 0.002852946, 0.1047612, 0.0005655963, 
    -6.049342e-05, 0.041813, -9.78765e-06, 0.006636779, 0.04598662, 
    0.07463266, 0.07122434, 0.09584463, 0.2872189, 0.2975698, 0.2847842, 
    0.2061763, 0.1749573, 0.2896655, -0.0001037209, -4.365303e-05, 
    0.03045999, 0.1718322, 0.1075018, 0.1258211, 0.158461, 0.2328437, 
    0.2632036, 0.06317811,
  0.09005564, 0.2304213, 0.2919995, 0.2916425, 0.07267098, 0.01254701, 
    0.05658199, 0.2370423, 0.1777349, 0.1209846, 0.1520509, 0.2291587, 
    0.3846611, 0.3369495, 0.3277416, 0.3739433, 0.2939951, 0.2466866, 
    0.1671372, 0.07656375, 0.06221329, 0.01440933, 0.1309931, 0.2642365, 
    0.175694, 0.227427, 0.3009599, 0.2933224, 0.1898236,
  0.2325395, 0.2340498, 0.2592915, 0.2396379, 0.1935737, 0.1647158, 
    0.1831938, 0.1852642, 0.3008234, 0.2544026, 0.1849832, 0.3515022, 
    0.2050143, 0.2592905, 0.1903276, 0.4305704, 0.4151414, 0.5534891, 
    0.3560304, 0.1637359, 0.2359135, 0.3180177, 0.3350702, 0.7062925, 
    0.4046113, 0.2924178, 0.3801385, 0.4578388, 0.2078469,
  0.6114392, 0.3388812, 0.4438388, 0.3148809, 0.3747179, 0.3670458, 
    0.4580024, 0.5967436, 0.4005775, 0.2875178, 0.477195, 0.3466103, 
    0.4206564, 0.3951228, 0.3948108, 0.3969529, 0.5269533, 0.3998089, 
    0.3275949, 0.3424075, 0.2927654, 0.3798759, 0.2633879, 0.2627037, 
    0.2225295, 0.2964592, 0.2098569, 0.09299441, 0.4789909,
  0.2418648, 0.3420234, 0.3670823, 0.3850687, 0.4336777, 0.3588603, 
    0.3626347, 0.4049642, 0.5750643, 0.4799433, 0.4108965, 0.3795226, 
    0.3698671, 0.3447286, 0.409811, 0.4412932, 0.4613446, 0.3969493, 0.35677, 
    0.312418, 0.2347423, 0.2695208, 0.2909912, 0.3641625, 0.2780662, 
    0.3789611, 0.2705198, 0.2133652, 0.2242533,
  0.3021533, 0.2996509, 0.2971484, 0.294646, 0.2921436, 0.2896411, 0.2871387, 
    0.2712997, 0.2778864, 0.2844731, 0.2910598, 0.2976465, 0.3042332, 
    0.31082, 0.3497819, 0.3454779, 0.3411739, 0.3368699, 0.3325658, 
    0.3282618, 0.3239578, 0.276049, 0.2762687, 0.2764885, 0.2767082, 
    0.2769279, 0.2771477, 0.2773675, 0.3041553,
  0.2091256, 0.106077, 0.1253612, 0.05670077, 0.02559028, -0.0009822197, 0, 
    0, 0, 0.003044943, 0.08402709, 0.2370608, 0.3015567, 0.1272074, 
    0.1577504, 0.1913215, 0.2108411, 0.2024416, 0.1588838, 0.1451054, 
    0.3408817, 0.2822221, 0.2206954, 0.1469794, 0.1890288, 0.1674945, 
    0.2028368, 0.1854436, 0.2186564,
  0.2338426, 0.271326, 0.2234055, 0.1399172, 0.09408676, 0.03009475, 
    0.1231386, 0.3294009, 0.2461533, 0.2180738, 0.1800737, 0.1318161, 
    0.2509412, 0.2013265, 0.276323, 0.4167909, 0.3234861, 0.322437, 
    0.4137667, 0.4276369, 0.3802723, 0.4433229, 0.3656972, 0.5285414, 
    0.4316757, 0.374323, 0.3557947, 0.2915448, 0.2378741,
  0.3766471, 0.4380992, 0.5396127, 0.3997581, 0.5043485, 0.4386164, 
    0.3227977, 0.4895763, 0.4701507, 0.2035983, 0.2127537, 0.3735371, 
    0.3714527, 0.3685337, 0.2941345, 0.3543871, 0.3799374, 0.4275263, 
    0.2748894, 0.1966397, 0.2697889, 0.2916779, 0.3532958, 0.3439319, 
    0.3579172, 0.3573249, 0.2871619, 0.3153216, 0.2978357,
  0.2957299, 0.3243884, 0.3246271, 0.2905907, 0.3391399, 0.3154443, 
    0.3164715, 0.2676447, 0.2868536, 0.2811396, 0.2736566, 0.3058837, 
    0.2565529, 0.2814801, 0.1887322, 0.2055397, 0.2361754, 0.2627112, 
    0.2765079, 0.3372115, 0.3695852, 0.3349179, 0.3177211, 0.2330917, 
    0.07265328, 0.217257, 0.3705339, 0.5197024, 0.3589158,
  0.2973046, 0.2582014, 0.1526486, 0.2423393, 0.2769847, 0.275144, 0.2870574, 
    0.2720461, 0.2543966, 0.1129029, 0.1390837, 0.09412436, 0.03278606, 
    0.1610086, 0.1238305, 0.246282, 0.1974359, 0.1692386, 0.117349, 
    0.09171996, 0.1246361, 0.1329864, 0.1803544, 0.2961836, 0.04106047, 
    0.1833819, 0.2534239, 0.2421088, 0.3148446,
  0.2825251, 0.09138247, 0.0204892, 0.1247579, 0.1348232, 0.2316979, 
    0.2091264, 0.2264621, 0.2632231, 0.08192088, 0.01679049, 0.001973658, 
    0.05114297, 0.1070237, 0.1940896, 0.1970576, 0.1102446, 0.06164581, 
    0.175223, 0.2175114, 0.1253261, 0.2603781, 0.2623994, 0.0007004038, 
    0.06958182, 0.2048707, 0.2019166, 0.2226985, 0.1797172,
  0.3419575, -8.061135e-05, 0.01259748, 0.04474577, 0.07370404, 0.06757731, 
    0.1120879, 0.08582056, 0.08659478, 0.0005476461, 2.651476e-08, 
    1.960744e-06, 0.1024012, 0.1244815, 0.1671571, 0.1316956, 0.1027835, 
    0.1495061, 0.1077034, 0.1063924, 0.197107, 0.386672, 0.5020232, 
    -0.0002831694, 0.01863494, 0.03749907, 0.1475144, 0.1506543, 0.390163,
  0.08001942, 0.02390597, 2.838552e-05, 0.01400664, 0.05496775, 0.06234304, 
    0.1035425, 0.08205901, 0.06011396, 0.06278103, 0.02615195, 0.03204416, 
    0.1341639, 0.1058312, 0.04003663, 0.04471767, 0.04336291, 0.03659658, 
    0.03199545, 0.02703825, 0.1570991, 0.5008516, 0.05097109, 0.0153641, 
    0.004715177, 9.052036e-07, 0.1418704, 0.25916, 0.4524308,
  0.1723838, 0.1535524, 0.006571724, 0.02072724, 0.08354048, 0.08027244, 
    0.07842952, 0.03877845, 0.05623326, 0.1455579, 0.07228439, 0.04261705, 
    0.05364948, 0.06926465, 0.1116114, 0.03202962, 0.03925749, 0.05045994, 
    0.06198746, 0.08097723, 0.1223802, 0.0368457, 0.01444682, 0.01585066, 
    0.004486362, 0.1257002, 0.1298652, 0.09663403, 0.08371299,
  0.005452437, 0.0007699057, 0.0007196376, 0.002072172, -3.003986e-05, 
    0.07346058, 0.05641239, 0.04724937, 0.01345529, 0.03743432, 0.01417506, 
    0.1867899, 0.0738287, 0.07015487, 0.0428405, 0.08808771, 0.1003735, 
    0.1421306, 0.1335103, 0.1405082, 0.1342929, 0.1256517, 0.1567369, 
    0.03334209, 0.08521734, 0.1401351, 0.08131064, 0.05462951, 0.01405736,
  8.16096e-08, 1.209478e-07, 2.029885e-08, -2.41249e-12, 4.698771e-09, 
    -0.0003644534, 0.03837041, 0.02538895, 0.1023748, 0.07314805, 0.1112691, 
    0.04382828, 0.04931553, 0.0884855, 0.06940627, 0.04192451, 0.06767673, 
    0.1309362, 0.1945893, 0.2878836, 0.1344413, 0.1365096, 0.07400551, 
    0.02363654, 0.0913387, 0.1021228, 0.1459888, 0.02453829, 2.09559e-07,
  4.69357e-07, 0.0009756983, 0.0005247428, -1.583685e-09, 3.199834e-07, 
    1.159465e-08, -7.234528e-06, 0.203055, 0.3435401, 0.2414392, 0.1539499, 
    0.05993271, 0.08873272, 0.08423778, 0.08044938, 0.1675164, 0.1568658, 
    0.158537, 0.2392838, 0.0008986662, 0.02163544, 0.03489999, 0.04977712, 
    0.092025, 0.07111254, 0.08030985, 0.1075154, 0.1104084, 0.003341786,
  0.008892289, 0.005023358, 0.0003112958, 0.1221375, 0.0009433471, 
    -4.207753e-05, 0.04414415, 1.765044e-06, 0.003601221, 0.03176636, 
    0.06954663, 0.06641153, 0.1872833, 0.3200313, 0.3085718, 0.2576618, 
    0.1703285, 0.1602568, 0.3101096, 7.671166e-05, -0.0001037892, 0.02045033, 
    0.1513181, 0.1056528, 0.1059395, 0.129927, 0.2078105, 0.1574509, 
    0.07349245,
  0.06606434, 0.2626545, 0.2666631, 0.2782043, 0.05014844, 0.01256852, 
    0.04419621, 0.2184445, 0.1544907, 0.1210007, 0.1167347, 0.199813, 
    0.4471944, 0.3852613, 0.3616823, 0.3354875, 0.3087692, 0.2151643, 
    0.2058731, 0.07145103, 0.06484491, 0.008783178, 0.1230127, 0.2367551, 
    0.1678472, 0.4105136, 0.4193517, 0.3066488, 0.1878164,
  0.2313891, 0.2422375, 0.2473144, 0.1723413, 0.1774964, 0.1308087, 
    0.1203149, 0.1179261, 0.2886647, 0.2102069, 0.13758, 0.3370459, 
    0.2224537, 0.2715678, 0.2050999, 0.3721437, 0.4295381, 0.5410582, 
    0.3537722, 0.1491567, 0.1599946, 0.3038663, 0.5389161, 0.6709157, 
    0.4388897, 0.3145052, 0.4335121, 0.3560439, 0.2655162,
  0.5437791, 0.2681171, 0.416783, 0.297128, 0.3743924, 0.2767494, 0.4506584, 
    0.5732248, 0.3874847, 0.199385, 0.4708021, 0.3370332, 0.4234512, 
    0.4009832, 0.4170308, 0.4727645, 0.5737188, 0.38209, 0.4802509, 
    0.3510247, 0.4348477, 0.430087, 0.318093, 0.3138956, 0.3471171, 
    0.3458538, 0.1909007, 0.09885813, 0.5312696,
  0.4536183, 0.5994479, 0.4883493, 0.5312944, 0.5463031, 0.4317085, 
    0.4848868, 0.540543, 0.5050901, 0.4702333, 0.4106425, 0.3534606, 
    0.3916809, 0.3959857, 0.4191639, 0.450449, 0.5039952, 0.5455378, 
    0.436241, 0.3692553, 0.3851768, 0.2728712, 0.2926426, 0.4030856, 
    0.3661707, 0.4125169, 0.2580427, 0.2360451, 0.2896987,
  0.2722183, 0.2704413, 0.2686642, 0.2668871, 0.2651101, 0.263333, 0.2615559, 
    0.2432086, 0.2517309, 0.2602533, 0.2687756, 0.277298, 0.2858203, 
    0.2943427, 0.3568153, 0.3524265, 0.3480378, 0.343649, 0.3392603, 
    0.3348715, 0.3304828, 0.2885908, 0.2862343, 0.2838777, 0.2815212, 
    0.2791646, 0.2768081, 0.2744516, 0.27364,
  0.2283738, 0.1207343, 0.1266762, 0.07056126, 0.02605448, -0.0007817562, 
    5.779286e-06, 0, -8.781737e-09, 0.0004696399, 0.08274925, 0.2381753, 
    0.3152635, 0.09007886, 0.1551563, 0.2345293, 0.2369658, 0.2074074, 
    0.1591351, 0.1401686, 0.3549742, 0.2970614, 0.2097296, 0.1283768, 
    0.1660274, 0.1846946, 0.1702056, 0.1949353, 0.2350907,
  0.2205511, 0.2326217, 0.2170639, 0.08386702, 0.07234467, 0.03436491, 
    0.09206314, 0.3435152, 0.227445, 0.2260297, 0.1716343, 0.1190159, 
    0.1946231, 0.1716051, 0.3115197, 0.4334027, 0.3628326, 0.3984558, 
    0.4317912, 0.4490986, 0.3696558, 0.4582448, 0.4322362, 0.5527667, 
    0.4010831, 0.4415228, 0.4100542, 0.3389498, 0.2362783,
  0.4273534, 0.430819, 0.4769071, 0.3213904, 0.4192783, 0.3946901, 0.3042628, 
    0.5436543, 0.317682, 0.1342992, 0.1437733, 0.3065042, 0.3171678, 
    0.3402837, 0.3060657, 0.3176464, 0.3474623, 0.384661, 0.2143494, 
    0.172711, 0.2513435, 0.2779568, 0.370371, 0.327774, 0.3832931, 0.3933656, 
    0.3409542, 0.3808755, 0.3417106,
  0.2888878, 0.3036665, 0.3339966, 0.3238346, 0.3482847, 0.32384, 0.346597, 
    0.2456392, 0.2699465, 0.2642761, 0.2454877, 0.2845882, 0.2618607, 
    0.3049406, 0.1502235, 0.2109328, 0.2371511, 0.2415287, 0.2506503, 
    0.2993828, 0.3374841, 0.3282679, 0.3145261, 0.2162484, 0.0630753, 
    0.2596247, 0.406451, 0.4590414, 0.3645417,
  0.2406025, 0.1973784, 0.1232961, 0.2158139, 0.282295, 0.2577349, 0.2665441, 
    0.2331456, 0.222035, 0.05511177, 0.09311755, 0.04655432, 0.02818423, 
    0.1080841, 0.1222158, 0.1959309, 0.1520416, 0.1060099, 0.07423888, 
    0.06504843, 0.09764815, 0.1244298, 0.1530335, 0.3280554, 0.02670031, 
    0.1190425, 0.1745971, 0.167731, 0.254458,
  0.149812, 0.08772342, 0.01574774, 0.1528175, 0.1336531, 0.1308502, 
    0.0761208, 0.08640252, 0.1103872, 0.03124454, 0.02353626, 0.0006702708, 
    0.05339738, 0.04496325, 0.1325999, 0.139899, 0.080151, 0.03113665, 
    0.1244533, 0.1785201, 0.1307582, 0.127301, 0.1820797, 0.005246527, 
    0.06481491, 0.1488179, 0.11851, 0.1249662, 0.09124216,
  0.3427145, -0.0004551834, 0.01220225, 0.07007825, 0.0128999, 0.04081592, 
    0.06065712, 0.02961248, 0.04539057, 0.0004776512, 2.47798e-08, 
    -2.082215e-06, 0.0268866, 0.09366877, 0.1588943, 0.1168857, 0.06220628, 
    0.08285017, 0.04505938, 0.03999062, 0.06589215, 0.1224797, 0.2424098, 
    0.009507299, 0.005116802, 0.048843, 0.04722243, 0.06196677, 0.2183318,
  0.6118023, 0.1198198, 1.115079e-05, 0.01380883, 0.020632, 0.02930299, 
    0.05821529, 0.06126239, 0.01226576, 0.01981822, 0.02065834, 0.009625087, 
    0.1129579, 0.09840684, 0.03146484, 0.01392727, 0.01132733, 0.006680143, 
    0.006989383, 0.004054029, 0.04660524, 0.2831826, 0.3173898, 0.006582351, 
    0.001297817, 2.856505e-07, 0.04075849, 0.07661627, 0.3668169,
  0.1266638, 0.111556, 0.003727085, 0.02386934, 0.04765401, 0.04086427, 
    0.03794365, 0.0400924, 0.06362543, 0.09588365, 0.07108305, 0.04963067, 
    0.0303052, 0.02173245, 0.01578504, 0.004655037, 0.01693002, 0.02736059, 
    0.0432201, 0.06773682, 0.2012063, 0.3256969, 0.1052432, 0.006665295, 
    0.001586979, 0.0374185, 0.0362538, 0.1147733, 0.3824677,
  0.002640424, 0.0004478453, 0.0006648942, 0.0003274077, -0.0001398206, 
    0.03314953, 0.05941723, 0.03016001, 0.006545355, 0.02891015, 0.005090386, 
    0.1103568, 0.03399369, 0.04259998, 0.04921857, 0.05222432, 0.0539928, 
    0.1089187, 0.07068474, 0.136677, 0.0938298, 0.1201744, 0.1787957, 
    0.02126698, 0.0183215, 0.02986364, 0.05855305, 0.1677275, 0.007436402,
  7.512541e-08, 1.010742e-07, 1.439442e-08, -6.286843e-12, 4.664636e-09, 
    0.0787598, 0.02363465, 0.02510599, 0.06097357, 0.07681699, 0.1353167, 
    0.03558542, 0.0148939, 0.02160832, 0.01957703, 0.01922214, 0.02956708, 
    0.1000729, 0.1802922, 0.2269211, 0.06357877, 0.1293215, 0.009486137, 
    0.004476542, 0.06923542, 0.1131109, 0.1723325, 0.1645591, 1.996688e-07,
  4.251416e-07, 0.005577004, 2.158578e-05, -3.745006e-08, 2.736197e-07, 
    1.03478e-08, -5.10113e-05, 0.2250089, 0.3288314, 0.2421152, 0.1313864, 
    0.08204317, 0.1110525, 0.08842909, 0.1249637, 0.1194988, 0.1028165, 
    0.1275593, 0.2677415, 0.01216671, 0.02403606, 0.02876568, 0.0305006, 
    0.0462782, 0.05579853, 0.04838473, 0.07725877, 0.04178244, 0.004628694,
  0.004022879, 0.003453556, -3.040691e-05, 0.1401355, 0.0004987065, 
    -2.507689e-05, 0.0505982, 2.400272e-06, 3.185815e-05, 0.0234739, 
    0.07612914, 0.069689, 0.1488235, 0.2900067, 0.3020353, 0.2270624, 
    0.1320468, 0.1500344, 0.2807284, 0.0006393986, -0.0001196223, 0.02440555, 
    0.1396424, 0.0969697, 0.09854482, 0.1270149, 0.1705123, 0.1031401, 
    0.09240793,
  0.04501893, 0.2903248, 0.2555318, 0.2993861, 0.04487794, 0.01553915, 
    0.0340309, 0.2240705, 0.1314626, 0.1113372, 0.1007414, 0.1742107, 
    0.4153061, 0.4111994, 0.295513, 0.375962, 0.3269416, 0.1975061, 
    0.1631316, 0.07108761, 0.0712232, 0.006429002, 0.1044341, 0.2346792, 
    0.1766711, 0.4228125, 0.3868152, 0.2593278, 0.1332784,
  0.2034117, 0.2714032, 0.1908621, 0.1448647, 0.1689654, 0.1212593, 
    0.1152073, 0.09693924, 0.2640258, 0.1881097, 0.1640765, 0.3144485, 
    0.2499868, 0.2639468, 0.2083076, 0.3331262, 0.4289562, 0.5129816, 
    0.3415132, 0.1377266, 0.1032379, 0.2876444, 0.6557902, 0.6255856, 
    0.4258002, 0.2830102, 0.4384818, 0.2518609, 0.1765598,
  0.4550851, 0.2472594, 0.3957287, 0.2178057, 0.2849363, 0.2499971, 
    0.4358658, 0.5571984, 0.3713231, 0.1575357, 0.4407182, 0.3212338, 
    0.4452125, 0.3819176, 0.4423864, 0.4112904, 0.5621498, 0.3482407, 
    0.4036153, 0.4191917, 0.5557567, 0.6235093, 0.4612139, 0.3466875, 
    0.3758234, 0.3481214, 0.1688211, 0.07449381, 0.4811113,
  0.5697713, 0.5003242, 0.6188172, 0.6148013, 0.6947517, 0.5261086, 
    0.5454149, 0.5397887, 0.5024055, 0.4274836, 0.3971541, 0.3666646, 
    0.3817346, 0.3381329, 0.3607816, 0.4926276, 0.5659893, 0.5928276, 
    0.5435431, 0.539812, 0.4666801, 0.3360796, 0.3388861, 0.4845597, 
    0.395373, 0.3930336, 0.2653456, 0.2822988, 0.3836386,
  0.2331161, 0.2317068, 0.2302975, 0.2288882, 0.2274789, 0.2260696, 
    0.2246603, 0.170131, 0.1797427, 0.1893543, 0.198966, 0.2085776, 
    0.2181892, 0.2278009, 0.2847356, 0.2806785, 0.2766213, 0.2725642, 
    0.2685071, 0.26445, 0.2603928, 0.2554762, 0.251331, 0.2471858, 0.2430406, 
    0.2388954, 0.2347502, 0.230605, 0.2342435,
  0.2175328, 0.1341003, 0.1193551, 0.0824532, 0.02669074, -0.0005833688, 
    5.779286e-06, 0, 0, 0.0001095919, 0.04144735, 0.2135155, 0.3495826, 
    0.05896301, 0.1752537, 0.2583403, 0.2847057, 0.2205217, 0.1482717, 
    0.1471714, 0.3539863, 0.3124297, 0.1779679, 0.1236207, 0.1375913, 
    0.1758099, 0.1762838, 0.2080416, 0.2474241,
  0.2079976, 0.1987581, 0.204268, 0.04879147, 0.04692022, 0.03529528, 
    0.0674115, 0.3404263, 0.2276049, 0.2097075, 0.1538576, 0.1257554, 
    0.1481382, 0.1387736, 0.3254914, 0.4584023, 0.4117232, 0.45185, 
    0.4365574, 0.4741432, 0.3386904, 0.4413792, 0.4332137, 0.5782526, 
    0.3583088, 0.5068956, 0.484877, 0.3858202, 0.2366923,
  0.4617933, 0.472595, 0.4053025, 0.2528011, 0.3314127, 0.3364784, 0.3067758, 
    0.4439486, 0.2072951, 0.09007139, 0.110268, 0.2388499, 0.2818691, 
    0.2954136, 0.2840191, 0.2915204, 0.307741, 0.3315433, 0.1848038, 
    0.1497076, 0.2373449, 0.2512046, 0.3945585, 0.2899914, 0.4036729, 
    0.4503402, 0.4032436, 0.457999, 0.394655,
  0.293165, 0.3163023, 0.3003802, 0.2822985, 0.2940736, 0.299523, 0.326451, 
    0.2268701, 0.234497, 0.2345751, 0.1916061, 0.2486378, 0.2001854, 
    0.274018, 0.1110262, 0.2022886, 0.2215898, 0.2131057, 0.2098155, 
    0.2338325, 0.2473428, 0.2799486, 0.2671314, 0.1914316, 0.05282916, 
    0.2745194, 0.4286216, 0.4452424, 0.3310201,
  0.1756968, 0.1221352, 0.102867, 0.1842738, 0.255397, 0.1822998, 0.19242, 
    0.1765546, 0.1419856, 0.02432411, 0.04223747, 0.02702397, 0.01256841, 
    0.0999928, 0.1288574, 0.1258443, 0.1098762, 0.06034584, 0.06413361, 
    0.04728395, 0.08517604, 0.1167661, 0.1463308, 0.330236, 0.01605301, 
    0.1063756, 0.1095429, 0.1544266, 0.2079628,
  0.05334385, 0.0388452, 0.01763066, 0.1192744, 0.07472476, 0.05308109, 
    0.03479035, 0.03297651, 0.04208569, 0.01141693, 0.01921642, 0.000686136, 
    0.0470358, 0.01773681, 0.08736682, 0.1211831, 0.07009123, 0.01587727, 
    0.09258905, 0.1734697, 0.0988069, 0.07540559, 0.0814336, 0.004879731, 
    0.04463756, 0.1355868, 0.08956452, 0.07402328, 0.05146815,
  0.1428, 0.001696871, 0.01217723, 0.03522374, -0.001232125, 0.02924427, 
    0.03228822, 0.004901444, 0.01284996, 0.001937839, 1.672712e-08, 
    -7.486098e-07, 0.006982978, 0.07095726, 0.136844, 0.03825433, 0.0238143, 
    0.03340496, 0.02180076, 0.008969189, 0.01829822, 0.03954535, 0.09115378, 
    0.03691348, 0.001442982, 0.06066317, 0.01644904, 0.02006472, 0.0817062,
  0.392598, 0.2745741, 1.505035e-06, 0.02797888, 0.006475885, 0.009270454, 
    0.0304762, 0.03748259, 0.000733432, -0.001079887, 0.01299257, 
    0.001948113, 0.0854083, 0.05111187, 0.01225082, 0.001941532, 
    0.0003516233, 0.0001498966, 0.0002949947, 0.0002674037, 0.01290618, 
    0.1017784, 0.3366604, 0.001858459, 0.0004735206, 3.229712e-07, 
    0.00509299, 0.02082616, 0.1437862,
  0.1211962, 0.09007622, 0.002209158, 0.01917884, 0.006895413, 0.005856398, 
    0.01778493, 0.01682032, 0.05160123, 0.05725561, 0.03384688, 0.01235213, 
    0.003944421, 0.005591675, 0.002723133, 0.0005236429, 0.004811661, 
    0.006367658, 0.01898396, 0.02921342, 0.0831176, 0.4488709, 0.3277746, 
    0.002641782, 0.0006212848, 0.00669442, 0.007262026, 0.02208559, 0.2701219,
  0.001899221, 0.0003080674, 0.0004434186, -7.519844e-05, -0.0001298094, 
    0.008125938, 0.07286189, 0.00399615, -0.0003613094, 0.01505477, 
    0.002070315, 0.01839062, 0.01108336, 0.0126621, 0.01751537, 0.03538363, 
    0.02623838, 0.04752945, 0.02420188, 0.1100325, 0.0493817, 0.07258854, 
    0.2097525, 0.01380556, 0.005820883, 0.00863213, 0.01611662, 0.08239365, 
    0.005828836,
  7.186703e-08, 8.652435e-08, 1.273238e-08, -1.727353e-12, 4.601119e-09, 
    0.2872516, 0.02803442, 0.01202498, 0.03928249, 0.04689045, 0.05445674, 
    0.00925476, 0.003607697, 0.008248649, 0.005256862, 0.002573493, 
    0.004309211, 0.03215871, 0.1105159, 0.16084, 0.08332705, 0.1003626, 
    0.001345555, -0.0006446482, 0.008481762, 0.03024661, 0.09614116, 
    0.167421, 1.921503e-07,
  3.962379e-07, 0.01036972, 3.071172e-06, -1.497414e-07, 2.431242e-07, 
    9.736697e-09, -4.856932e-05, 0.2376901, 0.2912503, 0.2170885, 0.08107911, 
    0.03019592, 0.05422031, 0.05184257, 0.08473322, 0.04514674, 0.05235559, 
    0.08389703, 0.2157191, 0.1146919, 0.02902574, 0.01311023, 0.01741546, 
    0.01149645, 0.01828058, 0.009513012, 0.01231686, 0.0175954, 0.008320858,
  0.003520631, 0.01415285, 8.523507e-05, 0.1558894, 1.191941e-05, 
    -3.047748e-05, 0.04316711, 2.646342e-06, 1.392244e-05, 0.02081135, 
    0.08511449, 0.02965493, 0.1222165, 0.2466798, 0.3013204, 0.1893945, 
    0.1086967, 0.1265938, 0.2655562, 0.0006041771, -0.000113373, 0.03958765, 
    0.116368, 0.08746938, 0.069423, 0.09627265, 0.122889, 0.06470902, 
    0.1126329,
  0.02087484, 0.2662472, 0.2470847, 0.281273, 0.04289469, 0.01996865, 
    0.03007656, 0.2270209, 0.1117958, 0.1060742, 0.08763231, 0.1868305, 
    0.39234, 0.3646099, 0.2589129, 0.3631787, 0.2676038, 0.1495384, 
    0.1669196, 0.06957586, 0.06707133, 0.002298675, 0.08241267, 0.2256944, 
    0.1679305, 0.3766783, 0.2996589, 0.2295119, 0.1291536,
  0.1874483, 0.2939143, 0.1543386, 0.1493379, 0.1833731, 0.1074264, 
    0.09381588, 0.08177249, 0.2408097, 0.1750528, 0.1642301, 0.2982916, 
    0.2740904, 0.267356, 0.1909378, 0.290102, 0.4409715, 0.471556, 0.3678509, 
    0.1344245, 0.08273655, 0.2371661, 0.5010355, 0.5903817, 0.4592176, 
    0.2140185, 0.4510967, 0.2583337, 0.1293003,
  0.3875576, 0.1700891, 0.3727023, 0.2064065, 0.2610815, 0.256134, 0.4206541, 
    0.5055029, 0.3542787, 0.1489045, 0.4536906, 0.3436493, 0.3764129, 
    0.4081264, 0.3807519, 0.3121068, 0.5236123, 0.3156892, 0.3167904, 
    0.3709114, 0.582696, 0.647425, 0.5670797, 0.4604884, 0.3935309, 
    0.3483121, 0.1432302, 0.06003398, 0.4365262,
  0.5119187, 0.4262098, 0.5256578, 0.5389243, 0.5749464, 0.5779215, 
    0.5457871, 0.5648583, 0.573751, 0.4608735, 0.4572514, 0.3454516, 
    0.3721916, 0.3514423, 0.3304008, 0.4848837, 0.59494, 0.6080446, 
    0.5774073, 0.5208172, 0.4431643, 0.2619045, 0.4154167, 0.629439, 
    0.385128, 0.3776433, 0.2615724, 0.3121069, 0.4075638,
  0.1082781, 0.1056106, 0.1029431, 0.1002756, 0.09760806, 0.09494056, 
    0.09227305, 0.06620404, 0.07868116, 0.09115829, 0.1036354, 0.1161125, 
    0.1285897, 0.1410668, 0.1682706, 0.1652074, 0.1621442, 0.159081, 
    0.1560178, 0.1529545, 0.1498913, 0.1637587, 0.1570123, 0.1502659, 
    0.1435195, 0.1367731, 0.1300267, 0.1232802, 0.1104121,
  0.2153779, 0.1122836, 0.1034772, 0.07834904, 0.02934959, -0.0005549125, 
    7.224949e-06, 0, 0, 0, 0.01828771, 0.1296811, 0.3809857, 0.03298771, 
    0.2109581, 0.2905722, 0.3088336, 0.1962766, 0.1320474, 0.1705271, 
    0.3498008, 0.316385, 0.149767, 0.114674, 0.09565201, 0.1961107, 
    0.1768716, 0.1923214, 0.263023,
  0.1872846, 0.1599191, 0.1833199, 0.02942714, 0.02148956, 0.02986574, 
    0.04273355, 0.3077582, 0.1994367, 0.183464, 0.1537077, 0.1386982, 
    0.1168936, 0.1099595, 0.3289121, 0.4431152, 0.4389183, 0.4881921, 
    0.4570227, 0.5109228, 0.3387643, 0.43231, 0.4376268, 0.5684224, 
    0.3170367, 0.6133707, 0.5118124, 0.39485, 0.2230299,
  0.458528, 0.464104, 0.3133407, 0.1916322, 0.266275, 0.2548478, 0.2888185, 
    0.3467046, 0.1301071, 0.06120241, 0.0859964, 0.1865782, 0.2520482, 
    0.2626664, 0.251515, 0.2533866, 0.2737163, 0.2709928, 0.1549645, 
    0.1327161, 0.2004174, 0.2114717, 0.343269, 0.255175, 0.4025648, 
    0.4613551, 0.4135569, 0.4971587, 0.3998625,
  0.2559677, 0.2824706, 0.2581661, 0.2295899, 0.2581014, 0.2578283, 
    0.2804811, 0.189445, 0.1984783, 0.19947, 0.1384894, 0.1913955, 0.1293852, 
    0.2101112, 0.07492321, 0.1566906, 0.1518056, 0.1523687, 0.1525777, 
    0.1684697, 0.1721515, 0.2121432, 0.1918034, 0.1630388, 0.03630499, 
    0.2672901, 0.3824596, 0.4394809, 0.2991711,
  0.1456617, 0.078398, 0.07095893, 0.140317, 0.2139946, 0.124671, 0.1348438, 
    0.132886, 0.08557887, 0.008821216, 0.02646595, 0.01672404, 0.007941167, 
    0.07642587, 0.115448, 0.09110524, 0.08592331, 0.03919695, 0.05280768, 
    0.03970476, 0.07153778, 0.1053116, 0.1235372, 0.3115343, 0.009897748, 
    0.08333343, 0.06685375, 0.1266694, 0.178303,
  0.02445857, 0.01324353, 0.01624355, 0.06151822, 0.04076589, 0.02605677, 
    0.01428234, 0.01554345, 0.02096692, 0.005984153, 0.01246157, 
    0.0003588212, 0.03688429, 0.009751544, 0.06079383, 0.09664869, 
    0.06335613, 0.005614739, 0.0687393, 0.1342408, 0.0534131, 0.05083828, 
    0.03547056, 0.0021273, 0.02910095, 0.1326779, 0.05876372, 0.04663579, 
    0.03067877,
  0.06860134, 0.00516711, 0.007271152, 0.008073453, -0.003574102, 0.01691684, 
    0.01364707, 0.001317098, 0.005038848, 0.003650798, 1.21806e-08, 
    1.005254e-07, 0.002411193, 0.03470933, 0.0969446, 0.01393802, 
    0.006718895, 0.008577799, 0.006930158, 0.002758695, 0.007167753, 
    0.01609447, 0.04142546, 0.0347659, 0.0006663602, 0.06782607, 0.002805868, 
    0.004611941, 0.03299761,
  0.1716441, 0.1672698, 1.343496e-06, 0.05981057, 0.001025656, 0.001389062, 
    0.006976007, 0.01513712, 0.0001477488, -0.001857138, 0.005416208, 
    0.0001852802, 0.0534697, 0.009337076, 0.001363602, 0.0003332726, 
    2.162233e-05, 4.504888e-05, 9.615149e-05, 0.0001211286, 0.004736677, 
    0.04246061, 0.1560533, 0.0006854523, 0.0003659504, 1.734628e-07, 
    0.001777205, 0.008089771, 0.05928462,
  0.02018733, 0.08988095, 0.00273649, 0.007358226, 0.0006455775, 0.000689025, 
    0.008744556, 0.004942021, 0.03992855, 0.03746727, 0.006971258, 
    0.001930108, 0.0002626288, 0.001046555, 0.001096511, 0.0002078713, 
    0.0003848056, 0.001062766, 0.002085771, 0.004295348, 0.01976913, 
    0.1966112, 0.1433713, 0.00219214, 0.0002858963, 0.002375733, 0.002131576, 
    0.005582682, 0.08095153,
  0.003635249, 0.0001963819, 0.0002037744, -0.0001183381, -5.236002e-07, 
    0.001568172, 0.06775068, 0.0003009051, -0.001575151, 0.003696334, 
    0.0002937173, 0.006261212, 0.004346268, 0.004084212, 0.008853146, 
    0.01269807, 0.007326457, 0.02506074, 0.01261846, 0.05848836, 0.01524877, 
    0.03626627, 0.2117914, 0.010698, 0.002056711, 0.003831628, 0.002798781, 
    0.01969958, 0.004476807,
  7.1934e-08, 7.408357e-08, 1.241035e-08, 1.231779e-11, 4.582766e-09, 
    0.2808451, 0.02078591, 0.00180995, 0.02780047, 0.009903987, 0.02929426, 
    0.001303311, 0.00075141, 0.003958303, 0.000966704, 0.0005281318, 
    0.001584056, 0.01161307, 0.05068864, 0.1244844, 0.01463759, 0.07497366, 
    0.0003697612, -0.001292384, 0.002749475, 0.01075811, 0.03424098, 
    0.04882457, 1.870435e-07,
  3.834626e-07, 0.008621518, 3.997216e-07, 5.362093e-06, 2.224412e-07, 
    9.598113e-09, -3.619767e-05, 0.2373961, 0.2552154, 0.1787576, 0.02795397, 
    0.008505716, 0.01893806, 0.02154831, 0.01910586, 0.01249863, 0.01066044, 
    0.05096185, 0.08177611, 0.2551178, 0.02652921, 0.006549686, 0.01154915, 
    0.005057621, 0.003197555, 0.002161109, 0.004051843, 0.01304835, 0.0171683,
  0.004243196, 0.004034404, 0.002415152, 0.1647619, -0.000301657, 
    -2.409606e-05, 0.03900139, 2.03881e-06, -9.954305e-05, 0.01799049, 
    0.08313083, 0.01399233, 0.0912246, 0.2140971, 0.2790096, 0.1396521, 
    0.07358085, 0.07837974, 0.2367596, 0.0008069737, -0.0001602271, 
    0.05385616, 0.09002046, 0.06813513, 0.04927495, 0.1099544, 0.08652171, 
    0.0437765, 0.0964381,
  0.009088858, 0.2389605, 0.2415754, 0.2467164, 0.03458456, 0.01465759, 
    0.01943201, 0.2136676, 0.09929964, 0.1015206, 0.07940912, 0.1902458, 
    0.3690644, 0.3281237, 0.235452, 0.3146925, 0.198391, 0.1162809, 
    0.1607996, 0.06603064, 0.05519603, 0.0009712562, 0.06865226, 0.2125556, 
    0.1509939, 0.3236392, 0.2549527, 0.19539, 0.1310737,
  0.1370505, 0.2788025, 0.1411404, 0.1389831, 0.1918411, 0.09118044, 
    0.07888132, 0.07269368, 0.2459827, 0.1559112, 0.1470285, 0.3357145, 
    0.263758, 0.2567901, 0.1675366, 0.2768179, 0.4254366, 0.426274, 
    0.3614433, 0.1338577, 0.06972615, 0.208952, 0.4143146, 0.5858844, 
    0.4694799, 0.192486, 0.4193915, 0.2146175, 0.1040472,
  0.3245775, 0.1190151, 0.3375463, 0.1608681, 0.2533034, 0.197917, 0.3918066, 
    0.4671451, 0.3355168, 0.1318291, 0.4633098, 0.3507857, 0.3249266, 
    0.3736222, 0.2909906, 0.2516353, 0.4812653, 0.2645753, 0.264377, 
    0.3185575, 0.6291285, 0.5847206, 0.5081657, 0.5495021, 0.3584663, 
    0.301066, 0.1339085, 0.05507572, 0.3814642,
  0.466543, 0.3209724, 0.4552566, 0.4587021, 0.4670796, 0.5079949, 0.5447581, 
    0.527018, 0.5355284, 0.5289613, 0.4240224, 0.3250575, 0.3775335, 
    0.3840547, 0.3533408, 0.4448286, 0.5328769, 0.5639296, 0.5554136, 
    0.4547088, 0.3748607, 0.2056605, 0.4055362, 0.6272358, 0.3355275, 
    0.3432306, 0.2514969, 0.2877444, 0.369495,
  0.005673736, 0.005389275, 0.005104815, 0.004820355, 0.004535894, 
    0.004251434, 0.003966974, -0.01514331, -0.00964655, -0.004149793, 
    0.001346964, 0.006843721, 0.01234048, 0.01783724, 0.02740064, 0.02620409, 
    0.02500754, 0.02381099, 0.02261444, 0.02141789, 0.02022134, 0.03300041, 
    0.02898466, 0.02496891, 0.02095317, 0.01693742, 0.01292167, 0.008905928, 
    0.005901304,
  0.2400678, 0.08253906, 0.08628913, 0.05479774, 0.01456643, -0.0002774977, 
    4.843556e-06, 0, 0, 0, -0.0006253705, 0.06288233, 0.2951778, 0.02032216, 
    0.2510845, 0.3533152, 0.365559, 0.2014536, 0.1011215, 0.2733449, 
    0.3741385, 0.3169712, 0.1134735, 0.08349164, 0.07570026, 0.2258028, 
    0.225662, 0.1691047, 0.2532063,
  0.1880099, 0.1293122, 0.1597586, 0.01814481, 0.007735169, 0.02306903, 
    0.02856677, 0.2411512, 0.1485697, 0.1262053, 0.1498034, 0.1238509, 
    0.09348864, 0.09441622, 0.3224474, 0.4673636, 0.4107219, 0.4201389, 
    0.4119561, 0.4753694, 0.3419431, 0.3862776, 0.4187096, 0.5164266, 
    0.3233514, 0.6438594, 0.4787873, 0.415145, 0.2215269,
  0.4046406, 0.4074171, 0.2544265, 0.1413182, 0.1960718, 0.1961722, 
    0.2550676, 0.2588718, 0.08808314, 0.04338166, 0.06265062, 0.1382016, 
    0.1967009, 0.2259798, 0.1975306, 0.2066879, 0.2211215, 0.2115481, 
    0.1227384, 0.1100479, 0.1623283, 0.1589882, 0.2602378, 0.2000035, 
    0.3536589, 0.4150496, 0.3953871, 0.4659918, 0.3801057,
  0.2080818, 0.2287293, 0.2044431, 0.1850693, 0.207953, 0.206923, 0.224225, 
    0.141292, 0.1552669, 0.1487949, 0.08929148, 0.1277282, 0.08074152, 
    0.1453068, 0.04366209, 0.09949768, 0.09273709, 0.09335252, 0.09614787, 
    0.1129592, 0.1182984, 0.1279693, 0.1253073, 0.1314148, 0.02881799, 
    0.2182417, 0.2919471, 0.3736872, 0.2457296,
  0.1236019, 0.04744535, 0.04223032, 0.1031951, 0.1529725, 0.07578491, 
    0.09298489, 0.09350534, 0.04859818, 0.003998047, 0.01364373, 0.01014798, 
    0.003874221, 0.04898361, 0.1061786, 0.06355479, 0.05510341, 0.02766388, 
    0.04019735, 0.02956174, 0.05687297, 0.0837256, 0.08731418, 0.2797308, 
    0.004749209, 0.07027216, 0.04445921, 0.08886959, 0.1412229,
  0.01328475, 0.007550475, 0.01252541, 0.02801678, 0.02384509, 0.01989017, 
    0.007407937, 0.009482144, 0.01327536, 0.003830627, 0.007707015, 
    0.0001465285, 0.02523961, 0.005309138, 0.04621356, 0.07148808, 
    0.04495832, 0.002002834, 0.04637365, 0.08063262, 0.02875476, 0.03257278, 
    0.0205579, 0.001184156, 0.02047693, 0.09826929, 0.03972008, 0.02901748, 
    0.01768118,
  0.04116895, 0.004048298, 0.002696583, 0.00302506, -0.003564939, 0.00799107, 
    0.00553366, 0.0005943929, 0.002532499, 0.00113508, 9.91069e-09, 
    1.320208e-07, 0.001455338, 0.01734056, 0.0643609, 0.005171305, 
    0.001773192, 0.002718138, 0.001940777, 0.001209591, 0.003785773, 
    0.008767031, 0.02344799, 0.03229386, 0.0003005371, 0.06977779, 
    0.001246541, 0.002121897, 0.01737548,
  0.0858064, 0.07231794, 6.917241e-07, 0.07451002, 0.000397977, 0.0002864288, 
    0.00152623, 0.004777759, 6.548275e-05, -0.0008835343, 0.001794329, 
    8.4356e-05, 0.02874112, 0.001531995, 0.000208793, 0.0001385914, 
    6.461721e-06, 2.413195e-05, 4.567029e-05, 7.046314e-05, 0.002429019, 
    0.02269986, 0.08625775, 0.0005020347, 0.0002744552, 1.609555e-07, 
    0.001241615, 0.004288551, 0.03105217,
  0.007074707, 0.09544115, 0.001069424, 0.002607687, 0.0002344015, 
    0.0002497509, 0.00387085, 0.00167239, 0.03312426, 0.03270562, 
    0.001551054, 0.0004357329, 3.638827e-06, 0.00041546, 0.0006159536, 
    0.0001101557, 0.0001636936, 0.0005043172, 0.0006150827, 0.001407067, 
    0.007232776, 0.08886445, 0.07626237, 0.001373732, 0.0001297615, 
    0.001313712, 0.001138149, 0.002682127, 0.03561316,
  0.004092318, 8.05889e-05, 6.328096e-05, -0.0001497068, 1.335273e-05, 
    0.0006083819, 0.04205233, 8.121351e-05, -0.001134915, 0.001111177, 
    4.775633e-05, 0.003261755, 0.001415699, 0.001477924, 0.005594941, 
    0.005170768, 0.005864922, 0.01374128, 0.008336802, 0.02611784, 
    0.005679713, 0.01796474, 0.1834009, 0.009853803, 0.0008487384, 
    0.001955266, 0.0006428378, 0.006432819, 0.008949221,
  6.66092e-08, 6.643064e-08, 1.237085e-08, 1.421186e-11, 4.56239e-09, 
    0.1562216, 0.01303229, 9.088459e-05, 0.02560625, 0.004626386, 0.01573009, 
    0.0003827613, 0.0001208093, 0.001267809, 0.0003563359, 8.013155e-05, 
    0.0008634904, 0.005813648, 0.01866574, 0.08883634, 0.004376656, 
    0.06311992, 0.0001838191, -0.001437866, 0.001453664, 0.004468181, 
    0.01565156, 0.02304463, 1.8449e-07,
  3.793298e-07, 0.007906542, -3.081284e-06, 4.09841e-06, 2.075974e-07, 
    9.588356e-09, -3.00938e-05, 0.2189753, 0.2187916, 0.1196412, 0.009719874, 
    0.003011208, 0.007211708, 0.008410488, 0.006566036, 0.005387905, 
    0.004145166, 0.01362898, 0.04189188, 0.2545891, 0.02093232, 0.003817764, 
    0.005216388, 0.002636505, 0.001385171, 0.001065783, 0.001986916, 
    0.009332247, 0.01639071,
  0.002848588, 0.0009167224, 0.003062909, 0.1561017, -0.000342294, 
    -7.064937e-06, 0.03497487, 3.53501e-07, -0.0002244941, 0.01453812, 
    0.07968309, 0.01594534, 0.06904715, 0.1754926, 0.2309891, 0.09765453, 
    0.04540166, 0.04055525, 0.2074998, 0.0007189718, -0.0001939304, 
    0.05502296, 0.06258494, 0.04877639, 0.03114175, 0.08060055, 0.05906108, 
    0.02767674, 0.06835273,
  0.003607857, 0.2203325, 0.2266886, 0.2040381, 0.02261825, 0.01002964, 
    0.01506086, 0.1852198, 0.08205113, 0.08987368, 0.07043271, 0.1803726, 
    0.3116488, 0.2932382, 0.2127284, 0.2625132, 0.1626357, 0.09494252, 
    0.1534311, 0.06159899, 0.04368746, 0.0005939944, 0.05143163, 0.1929932, 
    0.1287932, 0.3058376, 0.212529, 0.1686648, 0.08669984,
  0.09182182, 0.2522063, 0.1228984, 0.1187314, 0.1673851, 0.08141185, 
    0.06548523, 0.06531845, 0.2298604, 0.1359312, 0.1246019, 0.3154198, 
    0.2460853, 0.2089985, 0.1293561, 0.23196, 0.3950008, 0.3812632, 
    0.3111293, 0.1278079, 0.06443936, 0.1881086, 0.3074669, 0.5582963, 
    0.4157515, 0.1652327, 0.3883953, 0.1732387, 0.09154374,
  0.273086, 0.08074342, 0.2950916, 0.13081, 0.2018133, 0.1525814, 0.3520355, 
    0.4193008, 0.2961873, 0.1178155, 0.45052, 0.3156737, 0.2992901, 
    0.3180746, 0.2319159, 0.2135126, 0.4204035, 0.2109052, 0.2264095, 
    0.2477298, 0.5764744, 0.4976269, 0.4265311, 0.6151943, 0.305246, 
    0.2634064, 0.1374194, 0.03965976, 0.3056547,
  0.4538364, 0.2677064, 0.4081584, 0.3992878, 0.3977148, 0.4519249, 
    0.4812399, 0.4484982, 0.434006, 0.4925445, 0.3816081, 0.3019026, 
    0.3834999, 0.3884018, 0.3218572, 0.3898501, 0.4282162, 0.4648729, 
    0.4472339, 0.3997755, 0.3228263, 0.1643065, 0.3847093, 0.5909386, 
    0.2956661, 0.3051703, 0.2189629, 0.2451935, 0.3513692,
  0.003098136, 0.003332698, 0.003567261, 0.003801823, 0.004036385, 
    0.004270947, 0.00450551, 0.005081718, 0.007306512, 0.009531305, 
    0.0117561, 0.01398089, 0.01620569, 0.01843048, 0.01464553, 0.01304482, 
    0.01144412, 0.009843417, 0.008242714, 0.006642011, 0.005041308, 
    0.008097312, 0.00723866, 0.006380007, 0.005521354, 0.004662701, 
    0.003804049, 0.002945396, 0.002910486,
  0.2325847, 0.07793682, 0.06723715, 0.01670292, -0.002125592, 2.691675e-06, 
    4.129401e-06, 0, 0, 0, 0.0006252663, 0.01606436, 0.1767025, 0.01143961, 
    0.3257943, 0.3835696, 0.39098, 0.2144599, 0.08158051, 0.3397739, 
    0.4342893, 0.391324, 0.08140967, 0.05226725, 0.09771146, 0.2661154, 
    0.2199147, 0.1709024, 0.2721772,
  0.1708081, 0.1008336, 0.1484257, 0.01155957, 0.005614329, 0.01680674, 
    0.01848816, 0.1516695, 0.07290488, 0.08055893, 0.1186331, 0.08541128, 
    0.07698215, 0.07664729, 0.2927169, 0.430014, 0.3742065, 0.3147666, 
    0.3490531, 0.4079446, 0.3008645, 0.3378564, 0.3738586, 0.4493468, 
    0.3170657, 0.5661417, 0.4212284, 0.3840298, 0.2004236,
  0.333467, 0.3155752, 0.2035329, 0.1101989, 0.1539746, 0.1525213, 0.2283057, 
    0.2052596, 0.06523542, 0.02921292, 0.04608432, 0.1073966, 0.1466828, 
    0.1851248, 0.1501689, 0.1645273, 0.1714973, 0.1590638, 0.09553239, 
    0.08252643, 0.1233006, 0.1149751, 0.2030018, 0.1379237, 0.291634, 
    0.352627, 0.3600407, 0.3829226, 0.3191868,
  0.1665851, 0.1816141, 0.1600777, 0.1503322, 0.1712134, 0.1674002, 
    0.1815848, 0.1052845, 0.1212813, 0.1030589, 0.0560603, 0.07931548, 
    0.05058023, 0.09536387, 0.02362917, 0.06362235, 0.05597557, 0.05575106, 
    0.06145129, 0.0760915, 0.07965671, 0.08245529, 0.08133705, 0.1055006, 
    0.02668707, 0.1601088, 0.2167245, 0.2845479, 0.2000201,
  0.08448499, 0.02699369, 0.02859893, 0.06926896, 0.09380879, 0.04280237, 
    0.06068727, 0.05687104, 0.02812969, 0.002351649, 0.006673679, 
    0.005937885, 0.002043638, 0.030514, 0.09183052, 0.04382556, 0.03211554, 
    0.01738721, 0.0268226, 0.02034787, 0.03620638, 0.05438252, 0.05103186, 
    0.2449448, 0.00219369, 0.05782716, 0.03060969, 0.05702035, 0.09578131,
  0.008636649, 0.005778204, 0.008959865, 0.01321668, 0.01359424, 0.01203405, 
    0.005140889, 0.006850332, 0.009651323, 0.00276345, 0.004550022, 
    8.938659e-05, 0.0160101, 0.002868912, 0.03395752, 0.05191043, 0.02066461, 
    0.001026273, 0.02698332, 0.04478843, 0.01477876, 0.01936749, 0.01445909, 
    0.0008242474, 0.01981594, 0.0574453, 0.02338449, 0.01545391, 0.009953148,
  0.02779085, 0.003341603, 0.001200847, 0.001844941, -0.00273019, 0.00360614, 
    0.002547225, 0.0003436535, 0.001610254, 0.0001880951, 8.512664e-09, 
    1.078272e-07, 0.001007941, 0.008452485, 0.02622507, 0.00211737, 
    0.0009016513, 0.001016029, 0.0008093555, 0.0006714444, 0.00239926, 
    0.005632883, 0.01567029, 0.02608801, 0.0001441682, 0.06487861, 
    0.001061295, 0.001307155, 0.0112408,
  0.05293139, 0.03804607, 4.988699e-07, 0.06242516, 0.0002556692, 
    0.0001566118, 0.0007425692, 0.001447564, 3.853283e-05, -0.0003209834, 
    0.0007081294, 5.317607e-05, 0.01343203, 0.0004936426, 0.0001069094, 
    7.441509e-05, 3.601529e-06, 1.64196e-05, 2.760101e-05, 4.837118e-05, 
    0.001522781, 0.01464528, 0.05563291, 0.0003841636, 0.0002002516, 
    1.118219e-07, 0.001065484, 0.002750124, 0.01992439,
  0.003736685, 0.0778868, 0.0005171046, 0.001108346, 0.0001364806, 
    0.000153696, 0.001503893, 0.0008067749, 0.02685865, 0.03309951, 
    0.0006345396, 0.0001649162, -6.370551e-06, 0.0002806536, 0.0004078943, 
    7.02836e-05, 9.771193e-05, 0.0003121413, 0.0003550453, 0.0008137039, 
    0.004012286, 0.0500805, 0.04842336, 0.00172961, 0.0001544251, 
    0.0008608075, 0.0007048382, 0.0016533, 0.02119655,
  0.002917554, 3.430255e-05, 4.249039e-05, -0.0001620027, -3.537469e-06, 
    0.0003464415, 0.02253145, 4.318756e-05, -0.0005839205, 0.0003020974, 
    2.516963e-05, 0.002061612, 0.0004804555, 0.000751009, 0.002693279, 
    0.002248499, 0.004700466, 0.006516811, 0.003763399, 0.01009677, 
    0.002442601, 0.008191853, 0.1416662, 0.01037321, 0.0004264043, 
    0.00108236, 0.0003039832, 0.003197692, 0.01143848,
  6.513375e-08, 6.327869e-08, 1.243422e-08, -1.694406e-12, 4.58169e-09, 
    0.08540247, 0.006890937, 3.867096e-05, 0.0235401, 0.002400644, 
    0.00465671, 0.0001892319, 4.854975e-05, 0.0005400877, 0.0002277563, 
    1.598162e-05, 0.0005636231, 0.003659519, 0.01034447, 0.05740273, 
    0.0024345, 0.05382085, 0.000111185, -0.001288024, 0.0009119375, 
    0.002570719, 0.009111092, 0.01386779, 1.826592e-07,
  3.78579e-07, 0.006166301, -7.998461e-06, -2.110747e-06, 1.958953e-07, 
    9.858926e-09, -2.319607e-05, 0.2007707, 0.1861017, 0.06142737, 
    0.004063995, 0.001717243, 0.003015477, 0.002294353, 0.0034318, 
    0.003101912, 0.002601903, 0.004116811, 0.02601524, 0.2144973, 0.01570964, 
    0.004076947, 0.00305025, 0.001274108, 0.0008650112, 0.0007030642, 
    0.001173422, 0.001554125, 0.01278659,
  0.002469245, 0.0001399767, 0.002353275, 0.1435783, -0.0003024861, 
    -3.619185e-06, 0.03302277, -1.006865e-06, -0.0002590857, 0.01075193, 
    0.0673487, 0.01019476, 0.05361999, 0.1243534, 0.1775854, 0.06149134, 
    0.02697256, 0.01682333, 0.1940173, 0.0005818138, -0.0001900039, 
    0.04828355, 0.04001307, 0.02929366, 0.01718936, 0.04455026, 0.03117577, 
    0.009853485, 0.04767411,
  0.00133583, 0.2005623, 0.2015738, 0.1560836, 0.01570192, 0.007452243, 
    0.01135602, 0.1580832, 0.07070962, 0.08048333, 0.0611791, 0.1578663, 
    0.2439831, 0.2601768, 0.1689019, 0.2120084, 0.118957, 0.06829698, 
    0.1151721, 0.05701523, 0.0338931, 0.0004085637, 0.03646404, 0.1718272, 
    0.1086222, 0.2895514, 0.1670377, 0.1321801, 0.05469358,
  0.05663706, 0.2182536, 0.1028375, 0.09699813, 0.1450017, 0.06679033, 
    0.05216107, 0.05966807, 0.2032715, 0.1173961, 0.1008943, 0.2795554, 
    0.2235635, 0.1670713, 0.09654827, 0.1742177, 0.36213, 0.3270997, 
    0.2497706, 0.1194378, 0.05362252, 0.1653352, 0.2114234, 0.5042271, 
    0.3152558, 0.1209852, 0.3260721, 0.1171578, 0.0730817,
  0.2157108, 0.0494095, 0.2343008, 0.1118843, 0.1660544, 0.1276182, 
    0.2944169, 0.3506922, 0.2574283, 0.09961351, 0.4005834, 0.2717062, 
    0.2649727, 0.2571569, 0.1857262, 0.1830027, 0.3576083, 0.177489, 
    0.2028134, 0.1970424, 0.5041322, 0.4313707, 0.3612722, 0.5854584, 
    0.2724823, 0.2219324, 0.1729461, 0.03210131, 0.2290001,
  0.3922127, 0.2479551, 0.3563235, 0.3477, 0.3332677, 0.4022034, 0.4032859, 
    0.3572071, 0.3334168, 0.3842836, 0.3053526, 0.2476884, 0.3354602, 
    0.3563077, 0.2656391, 0.3067338, 0.3237973, 0.3654827, 0.3532422, 
    0.3373717, 0.3028815, 0.1300492, 0.3468288, 0.5629663, 0.2580109, 
    0.24949, 0.1845849, 0.2137215, 0.346188,
  0.002048941, 0.002089897, 0.002130852, 0.002171807, 0.002212763, 
    0.002253718, 0.002294673, -0.002103767, -0.0008625709, 0.0003786251, 
    0.001619821, 0.002861017, 0.004102213, 0.005343409, 0.007209148, 
    0.006448855, 0.005688562, 0.004928269, 0.004167976, 0.003407683, 
    0.00264739, 0.002208186, 0.001686327, 0.001164469, 0.0006426107, 
    0.0001207525, -0.0004011058, -0.0009229641, 0.002016177,
  0.1668127, 0.07191476, 0.03618788, 0.002909273, 4.15563e-05, 0, 0, 0, 0, 0, 
    7.261468e-05, 0.01042767, 0.1167623, 0.007659262, 0.3128671, 0.3190521, 
    0.3842901, 0.2480711, 0.07325004, 0.4150492, 0.4978317, 0.4867355, 
    0.07210984, 0.04112202, 0.09586191, 0.2791609, 0.2093614, 0.169221, 
    0.2945835,
  0.1354641, 0.07823978, 0.1088311, 0.007219588, 0.003040053, 0.008967485, 
    0.01100144, 0.09924928, 0.02222312, 0.0394401, 0.07411205, 0.07224645, 
    0.06754299, 0.06798375, 0.270004, 0.3674767, 0.3328843, 0.2663046, 
    0.3026157, 0.3412549, 0.2650981, 0.295289, 0.3351167, 0.3940102, 
    0.3137333, 0.4785451, 0.348217, 0.3110193, 0.1987804,
  0.2883577, 0.2551634, 0.1736756, 0.09209005, 0.1304095, 0.1278076, 
    0.2128263, 0.1757012, 0.05332543, 0.02278354, 0.03672796, 0.08486729, 
    0.1197542, 0.1560252, 0.1179121, 0.1352434, 0.1418574, 0.1302701, 
    0.07959481, 0.06640455, 0.1010593, 0.08853965, 0.1691964, 0.1035178, 
    0.2465057, 0.3056427, 0.3261562, 0.3324151, 0.2622934,
  0.1435431, 0.1543484, 0.1312267, 0.1311137, 0.1460942, 0.1418503, 
    0.1538809, 0.08383796, 0.09833345, 0.07448303, 0.03820185, 0.05270391, 
    0.03626306, 0.06577854, 0.01391993, 0.04247219, 0.0386026, 0.03685636, 
    0.04403111, 0.05504057, 0.05018401, 0.05786385, 0.05970426, 0.09267464, 
    0.02159373, 0.1242148, 0.1675533, 0.2197714, 0.1652052,
  0.05659565, 0.01558541, 0.02039588, 0.05022601, 0.06251966, 0.02601785, 
    0.04067106, 0.03544245, 0.01822031, 0.00162974, 0.00436373, 0.003898286, 
    0.001416837, 0.0179704, 0.07690388, 0.03046959, 0.02062086, 0.01068188, 
    0.01876756, 0.01353768, 0.02465894, 0.03456349, 0.03213352, 0.211655, 
    0.001301526, 0.04518316, 0.02115211, 0.04082358, 0.06708027,
  0.006640392, 0.004156902, 0.006207072, 0.007311557, 0.008025038, 
    0.006685687, 0.004039407, 0.005521068, 0.00770538, 0.002202437, 
    0.003163418, 7.252047e-05, 0.01049463, 0.001717294, 0.0209811, 
    0.03002588, 0.01029308, 0.0007521379, 0.01470012, 0.02710779, 
    0.007760079, 0.01165435, 0.01135886, 0.0006343086, 0.01850578, 
    0.03795193, 0.01210375, 0.008645924, 0.005761873,
  0.02095607, 0.002436677, 0.0006641538, 0.001309042, -0.002017975, 
    0.001680802, 0.00150749, 0.0002359757, 0.001179788, 8.960557e-05, 
    7.685691e-09, 9.082208e-08, 0.000775308, 0.004321961, 0.01540518, 
    0.001283253, 0.0006112042, 0.0006637769, 0.0005018756, 0.0004439246, 
    0.001740877, 0.004136628, 0.01185184, 0.02154533, 9.057867e-05, 
    0.06072976, 0.0008791382, 0.0009495633, 0.008314402,
  0.0378048, 0.02483303, 2.216167e-07, 0.04706315, 0.0001900617, 
    0.0001102456, 0.0005147143, 0.0006574602, 2.706681e-05, -0.0001079084, 
    0.0004428513, 4.043408e-05, 0.006821484, 0.0003009588, 6.113962e-05, 
    5.435368e-05, 2.535243e-06, 1.27696e-05, 1.96027e-05, 3.706866e-05, 
    0.001102803, 0.01078631, 0.04083057, 0.002937697, 6.278756e-05, 
    7.339484e-08, 0.0008645981, 0.002018092, 0.01458103,
  0.00247412, 0.05335152, 5.220557e-05, 0.0006552648, 9.734113e-05, 
    0.0001264742, 0.0007447915, 0.0004325009, 0.02343955, 0.03733567, 
    0.0003831829, 0.0001079553, 1.038569e-05, 0.000172184, 0.0003022056, 
    5.115021e-05, 6.96293e-05, 0.0002254303, 0.000252944, 0.0005702674, 
    0.002695482, 0.03438274, 0.03517513, 0.002226369, 0.000514957, 
    0.0006415352, 0.0005087584, 0.001186774, 0.01495601,
  0.001869146, 8.173682e-06, 9.978804e-06, -0.0001707002, -3.361971e-06, 
    0.0002378875, 0.01000306, 2.961215e-05, -0.0003941171, 0.0001396608, 
    2.020796e-05, 0.001469046, 0.0002979526, 0.000502278, 0.001413198, 
    0.001179217, 0.002203718, 0.003477825, 0.001960513, 0.004452922, 
    0.001142741, 0.003734634, 0.1160787, 0.0236746, 0.0002936217, 
    0.0006633727, 0.0002263776, 0.00203689, 0.01119715,
  6.395855e-08, 6.198723e-08, 1.254917e-08, -3.738431e-12, 4.036208e-09, 
    0.05665855, 0.0053011, 1.648993e-05, 0.02778525, 0.001195725, 
    0.001978736, 0.0001190074, 4.285201e-05, 0.0002715315, 0.0001696348, 
    6.767404e-06, 0.0004183661, 0.002635782, 0.006911304, 0.03867659, 
    0.001693666, 0.04821859, 7.752398e-05, -0.001222524, 0.0006597601, 
    0.001778458, 0.00617654, 0.009714143, 1.809678e-07,
  3.768662e-07, 0.003790359, -4.102562e-05, -1.393758e-06, 1.871569e-07, 
    1.010089e-08, -2.292494e-05, 0.1935878, 0.1638867, 0.03092145, 
    0.002258661, 0.001008788, 0.001778802, 0.001309529, 0.002110321, 
    0.002296045, 0.001904423, 0.002123066, 0.01893387, 0.1738502, 0.01268933, 
    0.01299667, 0.00595349, 0.0007443228, 0.0006294069, 0.0005350754, 
    0.0008251849, 0.0007214127, 0.009076392,
  0.001690614, 0.0001138228, 0.001758628, 0.1332438, -0.0002594212, 
    -2.240962e-06, 0.03057083, 2.684272e-07, -0.0002313259, 0.008912144, 
    0.05961461, 0.007081971, 0.03819165, 0.08640407, 0.1221749, 0.03557768, 
    0.01474794, 0.008181338, 0.1559345, 0.0004374216, -0.0001990389, 
    0.03979824, 0.0257848, 0.01526291, 0.009892656, 0.01927269, 0.01898725, 
    0.005662637, 0.03562159,
  0.0007238813, 0.180359, 0.1694858, 0.1219564, 0.01208993, 0.005884731, 
    0.009036304, 0.1411213, 0.0673495, 0.0734156, 0.05312865, 0.1433179, 
    0.1769908, 0.1970586, 0.1210142, 0.1583585, 0.08833638, 0.05158704, 
    0.08245102, 0.05660728, 0.02820579, 0.0003350335, 0.02630577, 0.1516313, 
    0.09276422, 0.2378871, 0.1214363, 0.0877914, 0.02854041,
  0.03732428, 0.185962, 0.08538645, 0.09259715, 0.130693, 0.05611186, 
    0.03984082, 0.05493622, 0.1835693, 0.1055897, 0.09085497, 0.2469922, 
    0.2018951, 0.1328255, 0.07253437, 0.1360579, 0.3313372, 0.2826585, 
    0.2128705, 0.1075648, 0.05037348, 0.1478411, 0.1411266, 0.4404898, 
    0.2370367, 0.09107482, 0.2454448, 0.07885107, 0.05685191,
  0.1595405, 0.02646834, 0.1940735, 0.09624843, 0.1331239, 0.1023641, 
    0.2511247, 0.297884, 0.2210609, 0.08124826, 0.3546289, 0.2382233, 
    0.2397371, 0.2177648, 0.1633962, 0.1568667, 0.3157844, 0.1524107, 
    0.1844739, 0.1540396, 0.4477173, 0.3800526, 0.3087641, 0.5456927, 
    0.2270896, 0.1890994, 0.2657747, 0.02631168, 0.179205,
  0.3442481, 0.2166435, 0.3308872, 0.283711, 0.2865043, 0.364023, 0.3432418, 
    0.2894428, 0.2695129, 0.2930908, 0.2444079, 0.2062417, 0.2875557, 
    0.3062106, 0.2269878, 0.2405367, 0.2552183, 0.293668, 0.2764024, 
    0.2962394, 0.260017, 0.1077615, 0.3025665, 0.5369272, 0.2285324, 
    0.2039462, 0.1578124, 0.1923948, 0.330694,
  0.001871879, 0.001887264, 0.001902649, 0.001918034, 0.001933419, 
    0.001948804, 0.00196419, -0.0002098269, 0.0002728744, 0.0007555758, 
    0.001238277, 0.001720979, 0.00220368, 0.002686381, 0.0008262972, 
    0.0005995916, 0.0003728861, 0.0001461806, -8.05249e-05, -0.0003072304, 
    -0.0005339359, 0.001227866, 0.0009564845, 0.0006851035, 0.0004137225, 
    0.0001423415, -0.0001290395, -0.0004004205, 0.001859571,
  0.1019444, 0.04080886, 0.002605122, 0.0015511, 6.19978e-05, 0, 0, 0, 0, 0, 
    9.359483e-05, 0.009637594, 0.06427655, 0.007427601, 0.3020667, 0.2513164, 
    0.3423837, 0.2825433, 0.1092383, 0.4635399, 0.5343727, 0.5315215, 
    0.07876337, 0.03534696, 0.08289553, 0.2137496, 0.1799161, 0.1842979, 
    0.2484508,
  0.1224404, 0.07310323, 0.09270545, 0.005778538, 0.002676624, 0.007131597, 
    0.0115037, 0.08975045, 0.02050478, 0.03513893, 0.03270141, 0.043563, 
    0.0614982, 0.06196385, 0.2666392, 0.3364654, 0.3053706, 0.233729, 
    0.2685132, 0.3074242, 0.2332729, 0.2785338, 0.3117864, 0.3683767, 
    0.2966637, 0.4187712, 0.3133215, 0.2679231, 0.1780968,
  0.2593272, 0.2274133, 0.1620655, 0.08369321, 0.120246, 0.1173014, 
    0.2044074, 0.16558, 0.04868031, 0.01954782, 0.03172097, 0.07515039, 
    0.1084044, 0.1378371, 0.101463, 0.1208348, 0.1282937, 0.1194222, 
    0.0709095, 0.05860677, 0.08622524, 0.07274286, 0.1445022, 0.086848, 
    0.2269094, 0.2783084, 0.3136421, 0.305007, 0.235408,
  0.1229191, 0.1292145, 0.1105384, 0.1079612, 0.1291578, 0.1235417, 
    0.1365571, 0.07269628, 0.0860233, 0.06158945, 0.03014187, 0.04037958, 
    0.03028461, 0.05146721, 0.01057367, 0.03374505, 0.03064408, 0.02801972, 
    0.03568411, 0.0452252, 0.03796631, 0.0445155, 0.04962943, 0.1060193, 
    0.01658977, 0.1028872, 0.1371341, 0.1831767, 0.1443216,
  0.04487869, 0.01077477, 0.01656314, 0.04036287, 0.04626632, 0.01815702, 
    0.02986537, 0.02490289, 0.01332924, 0.001345241, 0.003472853, 
    0.002996899, 0.001102904, 0.01168715, 0.0665618, 0.02296982, 0.0155485, 
    0.00779003, 0.01452103, 0.01074985, 0.01895058, 0.02502341, 0.02201446, 
    0.2011117, 0.0009536049, 0.03604842, 0.01612199, 0.03347026, 0.04910985,
  0.00567149, 0.003441765, 0.01149446, 0.004990493, 0.00569467, 0.004846751, 
    0.003469432, 0.004815679, 0.006662245, 0.001893523, 0.002473538, 
    6.051187e-05, 0.008039201, 0.001288082, 0.01333655, 0.0186925, 
    0.006277923, 0.0006317742, 0.009984461, 0.01588767, 0.004943313, 
    0.008386923, 0.00968103, 0.0005422775, 0.02765446, 0.02757524, 
    0.007417451, 0.005895686, 0.003835322,
  0.01758247, 0.002204967, 0.0004330941, 0.001064276, -0.001905596, 
    0.001070115, 0.001134302, 0.0001925986, 0.000982702, 8.610418e-05, 
    7.347013e-09, 9.181096e-08, 0.0006597358, 0.002937445, 0.008780468, 
    0.0009826025, 0.0004843656, 0.000540964, 0.0003860107, 0.0003449439, 
    0.001437031, 0.003438858, 0.01003041, 0.01885665, 5.843294e-05, 
    0.08059342, 0.0007603366, 0.000777143, 0.006890839,
  0.03054776, 0.01929393, -6.677239e-08, 0.03664213, 0.0001593519, 
    9.238803e-05, 0.0004169061, 0.0004546242, 2.248327e-05, -0.0001423944, 
    0.0003530083, 3.432264e-05, 0.00451915, 0.0002328145, 4.898935e-05, 
    4.53967e-05, 2.119191e-06, 1.106337e-05, 1.652633e-05, 3.19992e-05, 
    0.000917858, 0.008981816, 0.03343009, 0.04450237, -0.0002081984, 
    1.531047e-07, 0.0007291919, 0.001674352, 0.01201783,
  0.001919925, 0.08082091, -5.854422e-05, 0.0004739848, 8.063585e-05, 
    0.0001076603, 0.0005097614, 0.0002988664, 0.03550098, 0.05342144, 
    0.0002989986, 8.471881e-05, 1.547704e-05, 0.000117675, 0.0002479112, 
    4.270887e-05, 5.758435e-05, 0.0001859143, 0.0002143293, 0.0004634281, 
    0.002137246, 0.02709979, 0.02858912, 0.00218143, 0.007793718, 
    0.0005376305, 0.0004100538, 0.0009656023, 0.01196796,
  0.003776803, -2.510261e-05, 4.967153e-06, -0.000147432, -2.720114e-06, 
    0.000194807, 0.009243973, 3.457465e-05, -0.002354343, 9.816274e-05, 
    1.806256e-05, 0.001170028, 0.0002185033, 0.0003968746, 0.0009597163, 
    0.0008097512, 0.00125724, 0.002390559, 0.001335734, 0.00278672, 
    0.0007340428, 0.002263554, 0.1552316, 0.03395924, 0.0002329688, 
    0.000513882, 0.0001865667, 0.001569375, 0.02684904,
  6.325149e-08, 6.121041e-08, 1.263623e-08, -3.600239e-12, -1.028369e-10, 
    0.04259692, 0.01053272, 1.57365e-05, 0.08821762, 5.168904e-05, 
    0.001252856, 8.830024e-05, 3.65436e-05, 0.0001845383, 0.0001402864, 
    5.048528e-06, 0.0003462681, 0.002142081, 0.005365079, 0.0275058, 
    0.001362574, 0.04589727, 6.163484e-05, -0.0020463, 0.0005364807, 
    0.001426216, 0.004801734, 0.007776477, 1.8118e-07,
  3.770725e-07, 0.002328441, -2.782991e-05, -6.812381e-07, 1.810734e-07, 
    1.026339e-08, -2.205783e-05, 0.2234803, 0.1682616, 0.0240498, 
    0.001563411, 0.0007229968, 0.001321664, 0.001102755, 0.001569788, 
    0.00190011, 0.00157679, 0.001562596, 0.01548035, 0.1495646, 0.01107623, 
    0.06774966, 0.03638523, 0.0005535757, 0.0005140252, 0.0004499339, 
    0.0006672136, 0.0005572251, 0.006475154,
  0.001366194, -0.0002378919, 0.001467276, 0.1321545, -0.000233997, 
    -1.575361e-06, 0.02698346, 6.564435e-07, -0.0002104091, 0.008459916, 
    0.0735774, 0.005587034, 0.02704406, 0.05697019, 0.09153861, 0.02318505, 
    0.009111668, 0.004945473, 0.1124224, 0.0002508201, -0.0002095789, 
    0.03884326, 0.02513544, 0.01045398, 0.007039376, 0.01250307, 0.01248725, 
    0.004322289, 0.02927959,
  0.0002518889, 0.1826622, 0.1624695, 0.1187145, 0.01020759, 0.004957352, 
    0.007796608, 0.1392134, 0.07511007, 0.08053517, 0.0609015, 0.1531136, 
    0.1332279, 0.1417874, 0.08465639, 0.1152586, 0.06882501, 0.04024014, 
    0.05780025, 0.06564488, 0.02715567, 0.001010793, 0.03316272, 0.166935, 
    0.08558206, 0.1812653, 0.08721341, 0.06169659, 0.01852482,
  0.02757332, 0.1931094, 0.0763039, 0.09964956, 0.1481299, 0.07290925, 
    0.05625196, 0.07821296, 0.2119662, 0.1342775, 0.105212, 0.2432123, 
    0.2074164, 0.1374072, 0.06046097, 0.1110381, 0.3355535, 0.2845004, 
    0.2249245, 0.1100815, 0.05824334, 0.1597012, 0.09830219, 0.4283188, 
    0.1846023, 0.07434774, 0.2036158, 0.06066, 0.04366459,
  0.1157222, 0.01727033, 0.1816732, 0.06866991, 0.1045323, 0.08549143, 
    0.2586278, 0.2883531, 0.2141492, 0.0917144, 0.3729547, 0.2467353, 
    0.2419053, 0.185973, 0.1552883, 0.1378447, 0.2968895, 0.1478737, 
    0.1675147, 0.1254081, 0.4068687, 0.3441477, 0.2966262, 0.511888, 
    0.1851609, 0.1685374, 0.3556955, 0.02153417, 0.1459498,
  0.3330589, 0.1927848, 0.3036271, 0.2442645, 0.2552659, 0.3414078, 
    0.3109087, 0.2503702, 0.2331537, 0.2496339, 0.2021393, 0.1769851, 
    0.2417011, 0.2593901, 0.1957289, 0.1998286, 0.2191452, 0.2549241, 
    0.2394413, 0.2570831, 0.2177191, 0.1010723, 0.276957, 0.5133287, 
    0.2046205, 0.1798583, 0.1372022, 0.1806233, 0.3021172,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.5757e-05, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3.595335e-10, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -6.505753e-06, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -7.327763e-05, -7.306319e-05, 0.002092247, 
    0, 0, -2.791655e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.297688e-06, 0.000614674, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, -4.082224e-06, 0, 0, 0, 0, 0, 0, 0, 0, -1.861105e-05, 0, 0, 
    0, 0, 0, 0, 0, 0, -2.47581e-05, 0, 0, 0, 0, 0,
  0, 8.053495e-05, 0.0003058382, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3.978134e-06, 
    -2.06794e-05, 0, 0, 0, 0, 0, 0, 0, 0, -9.775374e-06, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.0001478657, 0, 0, 0, -0.0002158521, -2.315168e-05, 
    0.004823857, 0, 0, 0.001665237, -2.29145e-05, 0, -2.371262e-05, 
    0.002546354, 0, 0, -2.269591e-05, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0.006712401, 0, 0, -9.501627e-05, -4.15447e-06, 
    0.0008465446, -3.084527e-05, 0.0001612802, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.204892e-05, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -2.630863e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.068622e-05, 0, 0, 0, 0, 
    0, 0, 0, -2.968707e-05, 0, 0, 0, 0,
  0, -8.055252e-06, 0, 0, 0, -6.340804e-05, -2.185235e-05, -2.910272e-05, 0, 
    0, 0, 0, 0, 0, -5.336392e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0.000715794, 0, 0, 
    0, 0, 0,
  0, 0.0003985132, 0.002113849, 0, 0, 9.433163e-05, 0, 5.222554e-05, 
    -6.320902e-06, -1.525033e-05, 0, 0, 0, 3.443036e-05, -9.305731e-05, 0, 0, 
    0, 0, 0, 0, 0, 0, 1.823394e-05, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -2.912538e-05, 0.00607908, -7.959956e-05, 0, 
    -1.835361e-05, 0.0003924075, 0.007715731, 0.01002597, 0, -8.703235e-05, 
    0.007849777, 0.001236176, -3.703789e-05, -0.0001610277, 0.00552292, 0, 
    -2.492219e-05, -1.535315e-05, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0.01029937, -4.617849e-07, 0, 0.0005479078, 0.0009246533, 
    0.001363896, -0.0001759661, 0.004312099, 0, 0, 0, 0, 0, 0, 0, 
    -8.888091e-05, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -4.912105e-05, 0.0004954412, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8.539172e-05, 3.707005e-05, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -7.439907e-05, -6.844195e-06, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0005116745, 0, 0, 0, 0, 
    0, 0, 0, -7.320221e-05, 0, 0, 0, 0,
  0, -3.246401e-05, 0, 0, -5.274641e-06, 8.782687e-05, -9.621735e-05, 
    0.0002189372, -1.660844e-05, 0, 0, 0, 0, 0, -0.0001829216, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.001508245, 0, 0, 0, 0, 0,
  0, 0.003234383, 0.003458254, 0, 0, 0.00408125, 0, 4.432279e-05, 
    -1.079164e-05, -4.098113e-05, 0, 0, 0, 0.0007068119, -0.0001497589, 0, 0, 
    0, 0, 0, 0, 0, 0, -1.40289e-05, 0, 0, 0.002087062, 0, 0,
  0, 0, 0, 0, 0, 0, 0.0009646955, 0.0081461, 0.002586214, -2.679266e-05, 
    0.0007008958, 0.003880844, 0.0269563, 0.0221167, -6.180635e-05, 
    0.004264117, 0.01724878, 0.006208977, 0.0001005564, 0.001275908, 
    0.01140116, 0.001628636, -0.0001312811, -7.237257e-05, -5.615747e-06, 0, 
    -1.597527e-05, 0, 0,
  0, 0, 0, 0, 0, 0, 0.0141993, -1.852609e-05, -6.08069e-06, 0.002908076, 
    0.005576957, 0.00330531, 0.003936287, 0.01681675, 0, -3.491811e-05, 0, 0, 
    0, 0, 0, 0.001063495, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 6.602271e-08, 0, 0, -8.15917e-05, 0.007043483, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0007681621, 0.001649573, 0, 
    0.0004397913, 0, 0, 0, 0, 0, 0, 0.0001786412, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7.79916e-05, 0, 0, 0, 0,
  0, 0, 0, 0.0003762679, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7.980918e-05, 0, 0, 0, 0, -0.0001029004, 0.00445903, -1.958373e-06, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.003142962, -1.653967e-05, 
    0, 0, 0, 0, 0, 0, 0.0002961442, 7.938496e-05, 0, 0, 0,
  0, -8.322149e-05, 0, 0, -1.501865e-05, 0.003302388, -4.042602e-05, 
    0.003589004, -4.982531e-05, 0, 0, 0, 0, 0, 7.752012e-05, -7.705691e-05, 
    -2.351224e-05, 0, 0, 0, 0, 0, 0, 0.004091916, -3.717223e-06, 0, 0, 0, 0,
  0, 0.005448278, 0.003966914, 0, 0, 0.009031678, 0, -7.02497e-06, 
    -2.672846e-05, -8.172462e-05, 0, 0, -1.17898e-06, 0.00195517, 
    0.0001373047, 0, 0, 0, 0, 0, 0, 0, 0, 0.0006224645, 0, -2.207251e-05, 
    0.005104896, 0, 0,
  0, 0, 0, 0, 0, 0, 0.002199977, 0.0126109, 0.0116702, -9.582568e-05, 
    0.001404359, 0.007466739, 0.04986932, 0.04227483, 0.0004967997, 
    0.008665108, 0.02857848, 0.01320206, 0.0007153497, 0.003835952, 
    0.01793315, 0.003957897, -0.0004524785, -3.113511e-05, -8.41408e-06, 
    0.0002422788, -3.993819e-05, -1.032384e-05, 0,
  0, 0, 0, 0, 0, 0, 0.01804549, 0.0003053079, -1.621517e-05, 0.005562137, 
    0.01465124, 0.008742746, 0.009409713, 0.02889866, 0, -7.298033e-05, 0, 0, 
    0, 0, 0, 0.002164118, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, -8.581587e-05, 0.003247149, 0, 0, -0.0001252106, 
    0.01352302, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -7.024717e-07, 
    -1.231658e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.004604574, 0.01020418, 0.003177779, 
    0.0005646132, 0, 0, 0, 0, 0, 0, 0.002841443, -8.349783e-06, 0, 
    -3.605636e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.804752e-05, 8.420373e-05, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2.552287e-05, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, -1.762389e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, -6.160865e-06, 0, 
    0.0009669603, 0, 0, 0, 0, 0, 0, 0, 0.002743187, -3.338615e-07, 
    -5.143549e-06, 0.000139609, 0,
  0, 0, 0, 0.007207765, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -7.981697e-07, 0, 0, 
    -7.811577e-05, 0.005023363, 0, 0, 0, 0, 0.0003254596, 0.006776284, 
    0.002560077, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.000396154, 0, 0, 0, 0, 0, 0, 0, 0, 0.005043859, 
    -0.0002456061, 0, 0, 0, 0, 0, 0, 0.001332081, 0.004245009, 0, 0, 0,
  0, -0.0002217041, 1.190447e-06, 0, -4.380783e-05, 0.0111532, 0.001612421, 
    0.01518704, -0.0001391747, 0, -1.795399e-06, 0, -2.70162e-05, 0, 
    0.000472085, -0.0001375361, 0.0008575217, 0, 0, 0, 0, 0, 0, 0.005711919, 
    4.674345e-05, 3.282354e-05, 0, 0, 0,
  0, 0.009155165, 0.004073877, 0, 0, 0.01237821, -1.560382e-05, 0.0002065862, 
    0.0003515723, -0.0001353321, 0, -6.058557e-06, 1.155491e-05, 0.002874162, 
    0.00126492, 0, 0, 0, 0, 0, 0, 0, 0, 0.003673846, -2.030123e-06, 
    -1.995698e-05, 0.009018335, 0, 0,
  0, 0, 0, 0, 0, 0, 0.004388765, 0.01983671, 0.02186377, -0.0002054507, 
    0.005204733, 0.02683449, 0.07591664, 0.08781605, 0.002482781, 
    0.009576365, 0.03834214, 0.02373434, 0.003080422, 0.00881198, 0.03014395, 
    0.008727594, 0.002530989, 0.000235959, -1.19753e-05, 0.00300706, 
    0.00212685, 1.812907e-05, 0,
  0, 0, 0, 0, 0, 0, 0.02467625, 0.0006778813, -2.45155e-05, 0.01010572, 
    0.02923658, 0.01935921, 0.0176272, 0.04661537, 0, -9.994677e-05, 0, 0, 0, 
    0, 0, 0.003863615, 0, -1.550373e-05, 0, -4.585543e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, -0.0004334941, 0.006655087, 0, 0, -0.0001691499, 
    0.01730021, 6.540828e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002547177, 
    -6.349888e-05, 0.002118462, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.613767e-06, 0, 0.01180659, 0.02247871, 
    0.00471177, 0.0007576483, 0, 0, 0, 0, 0, 0, 0.0100655, 0.001687206, 
    -3.766122e-05, 0.0003892668, -8.137938e-05, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3.714454e-05, 0, 0.006385124, 
    0.00477918, -2.496352e-05, 0, 0, 0, 0, -1.98496e-05, -1.018157e-05, 0, 0, 
    0, 0.00285634, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, -1.722868e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 5.823814e-06, 0.00118971, -1.664088e-05, 0.002718301, 0, 0, 0, 0, 
    0, -4.837222e-05, 6.909292e-05, 5.897817e-05, 0, 0.002771224, 0, 
    0.0005979455, 0.0002294579, 0.001316621, 0, 0, 0, 0.00647005, 
    -1.789648e-05, -2.734916e-05, 0.001278892, 0,
  0, 0, 0, 0.01706615, -5.545014e-06, 0, 0, 0, 0, 0, -5.713741e-05, 0, 0, 0, 
    0.0001154932, 0.001497951, 0, -5.445324e-06, 0.0003136821, 0.01094965, 
    0.000310898, 0, 0, 0, 0.003018945, 0.01721737, 0.007844293, 0, 0,
  0, 0.0001842961, -1.694404e-05, 0, -1.011609e-05, 0, 0, 0.00171755, 
    -1.779602e-07, 0, 0, 0, 0, -1.811965e-05, 0, -2.275094e-05, 0.01047501, 
    0.002099475, 0, -4.54215e-06, 0, 0, 0, 0, 0.002343163, 0.006780314, 
    -0.0001727849, 0, 0,
  0, 0.001042848, 0.001502603, 0, -0.0002130008, 0.02627334, 0.005170421, 
    0.03571124, -0.0002434913, 0, 0.0009014718, -8.80161e-05, -6.846995e-05, 
    -5.628464e-05, 0.003838937, -0.0002817374, 0.002748804, -8.766468e-07, 0, 
    0, 0, 0, 0, 0.01351877, 0.001290335, 0.0003753252, 0, 0, 0,
  0, 0.01835497, 0.005136091, 0, 0, 0.01710329, 0.0001677459, 0.002786787, 
    0.00145159, 0.0001068114, -5.301022e-05, -4.188932e-05, 0.0003444616, 
    0.00849333, 0.003350518, -2.224517e-06, 0, 0, 0, 0, 0, 0, -1.310224e-08, 
    0.009416408, 4.604428e-05, 4.132638e-05, 0.01147576, 0, 0,
  0, 0, 0, 0, 0, 0, 0.007740802, 0.03350649, 0.02962637, 0.001811903, 
    0.01215061, 0.05554377, 0.108276, 0.1251203, 0.01076053, 0.01632304, 
    0.05493282, 0.03688768, 0.007873355, 0.01856072, 0.04497602, 0.0138753, 
    0.005992282, 0.0009892933, 0.0003401783, 0.005446436, 0.003721008, 
    0.0007712964, 0,
  0, 0, 0, 0, 0, 0, 0.03090236, 0.003944351, 0.0007118878, 0.0155223, 
    0.04420342, 0.04025308, 0.02739176, 0.07320998, -1.769607e-05, 
    -9.061832e-05, 0, 0.001627077, 0, 0, 0, 0.01024256, 5.270876e-05, 
    -6.139309e-05, -1.145109e-05, -9.304517e-05, 0, 0, 0,
  0, 0, 0, 0.000170665, 0, 0, 0, 0.0005525477, 0.01319996, 0.0001264846, 
    0.0006430128, 0.001850608, 0.01977463, 0.0002193723, -2.995366e-05, 
    -6.942363e-06, -2.968839e-05, 0, 0.0006914982, 0, 0, -5.657382e-06, 
    0.0008750228, 0, 0.00760686, -4.033394e-05, 0.004200633, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0008915237, -6.459123e-05, 0.02378921, 
    0.03014508, 0.006162292, 0.002572651, 0.0006690131, 0.0001408072, 0, 0, 
    0, -2.749921e-06, 0.01453832, 0.008505635, 0.002632805, 0.007225121, 
    0.000649571, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.585591e-06, 0.001586352, 6.778596e-05, 
    0.01087747, 0.007806179, 0.002811321, 0.001422498, 0, 0, 0, 0.0001112312, 
    -2.552761e-05, 0, -3.142655e-05, -5.565343e-05, 0.005665439, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -1.262015e-06, 0, 0, 0, 0, -4.619478e-05, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, -9.965818e-06, 0.00187881, -2.290154e-05, -6.025109e-05, 
    0.0002292252, 0, 0, 0, 0, 0, 0.0007191277, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.0002035073, 0, 0,
  1.434414e-05, 0, 7.595296e-05, 0.002090981, 0.004926182, 0.001716842, 
    0.005577337, 0, 0, 0, 0, 0, 0.0001604081, 0.001446906, 0.0009063195, 0, 
    0.00366245, -7.204808e-06, 0.001436302, 0.001694408, 0.00530939, 
    -3.02886e-06, 0, 0, 0.01171266, -0.000116133, 0.002098412, 0.002806163, 
    -7.885994e-05,
  0, 0, 0, 0.02538593, 0.001966019, -4.834277e-06, 0, 0, 0, -2.977451e-09, 
    2.21314e-05, 8.787743e-07, -7.037528e-08, -1.403273e-06, 0.009635787, 
    0.01081483, -2.615483e-05, 0.001890991, 0.004548864, 0.01804963, 
    0.005746732, -7.621395e-10, 0, 0, 0.007518934, 0.03646438, 0.01382599, 
    5.0888e-05, 0,
  0, 0.0005427723, 6.969472e-05, -6.523186e-06, 4.321312e-05, 0, 0, 
    0.003535704, 0.001936699, 0, 2.027846e-07, 0, 2.030249e-07, 0.0001109324, 
    -5.417005e-06, 0.001533094, 0.02603132, 0.01642044, 0.0002909398, 
    -4.601044e-05, 0, 0, 0, 1.354352e-05, 0.005407744, 0.0103325, 
    0.005341509, 0, 0,
  0, 0.004784428, 0.003146142, -1.321276e-06, 4.278334e-05, 0.048008, 
    0.01448743, 0.05561177, 0.002448826, 0, 0.005214177, -3.113463e-05, 
    -0.0002237843, 0.0003698502, 0.01824134, 0.00463788, 0.01022738, 
    -8.416787e-06, 0, 0, 0, 0, -3.259438e-06, 0.04645807, 0.01976282, 
    0.0007838448, 0, 0, 0,
  0, 0.04267279, 0.01645075, 0, 0, 0.03150966, 0.0002645736, 0.01305137, 
    0.0204755, 0.005757101, 7.763391e-05, 0.00142495, 0.00133072, 0.03906375, 
    0.007137132, 3.322931e-05, 0, -1.542979e-05, 0, -3.280595e-07, 0, 
    3.344873e-08, 8.107166e-05, 0.05336991, 0.001957208, 0.0002412709, 
    0.01392788, -1.705606e-09, 0,
  0, 0, -1.01427e-07, 0, -1.088171e-05, 0, 0.0129186, 0.05102414, 0.05435415, 
    0.01053344, 0.02906235, 0.09709375, 0.1688647, 0.1600747, 0.03625111, 
    0.03312204, 0.08866996, 0.04969439, 0.01799912, 0.03423792, 0.05708691, 
    0.03221171, 0.02402728, 0.01533548, 0.002042655, 0.0129079, 0.009671158, 
    0.00260744, -1.542879e-05,
  0, 0, 0, -1.497422e-06, 0, 3.723266e-07, 0.03355201, 0.01453738, 
    0.009480495, 0.02374541, 0.06123719, 0.06619289, 0.05375194, 0.09423221, 
    0.0001805554, 0.003496295, 0.001077578, 0.007819276, 1.043343e-06, 
    -1.074192e-08, 0.0001053518, 0.02099389, 0.0004876212, 0.0009762377, 
    8.829295e-05, 0.0003772511, 0, 0, 0,
  0, 0, 0, 0.001324227, -2.821936e-10, 0, 0, 0.001335929, 0.01901946, 
    0.003317839, 0.0116154, 0.008261469, 0.02881887, 0.0006140961, 
    0.00740969, -2.823368e-05, 0.003145647, 0.00134565, 0.005513784, 0, 
    0.0004806765, -0.0002748712, 0.003136804, 0.0006474458, 0.009997948, 
    0.0008842768, 0.005488784, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.008901076, 0.01816062, 0.04858025, 
    0.0459695, 0.01651801, 0.009706277, 0.009700969, 0.007260328, 
    -8.452928e-08, 0, 0, -1.1656e-05, 0.0232841, 0.02184234, 0.01101291, 
    0.0234177, 0.00878907, 0.005286867, 0,
  0.001217436, -2.964018e-05, -1.431379e-05, 0, 0, 0, 0, 0, 0, 0, 0, 
    -0.0001063622, 0.007784186, 0.002220511, 0.01432184, 0.01017827, 
    0.01325121, 0.0106373, 0.0007553011, -1.540933e-05, 0, 0.002005504, 
    -7.417486e-05, 0.0003664907, 0.0014583, 0.001736412, 0.01278886, 
    0.0004840862, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.204328e-09, 0, 0, 0, 
    -1.270335e-05, 0, -1.465711e-06, -2.481143e-05, 0.0001634056, 
    -0.0001284008, -2.486518e-05, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  -7.979602e-05, 0.0001162287, 8.720454e-05, 0.003213052, 0.002352996, 
    0.001381084, 0.003956632, 0.002159399, 0, 0, 0, 0, 0, 0.002733965, 0, 0, 
    -4.046361e-06, 0, 0, 0, 0, -1.896039e-06, 0, 0, -1.12314e-06, 0, 
    0.001803025, 0, -1.440416e-05,
  0.002483225, 0, 0.002941644, 0.005434999, 0.01518034, 0.004709146, 
    0.008634786, 0, 0, 0, -2.460492e-15, 0, 0.003189423, 0.005745725, 
    0.01171949, 0.0003780391, 0.006815245, 0.00088805, 0.006050147, 
    0.005175186, 0.007537525, 0.001002878, 0, 0, 0.01841905, -0.0001897656, 
    0.006737897, 0.007557603, 0.003959914,
  1.369783e-06, -8.612146e-06, -6.178677e-06, 0.03890126, 0.006379568, 
    0.0001092889, -1.82814e-10, -1.445818e-07, -2.042096e-06, 3.461005e-05, 
    0.001950174, 0.002146392, 0.0004672283, 0.0001112458, 0.02528897, 
    0.01668584, -0.0003007876, 0.01730811, 0.03490487, 0.03558692, 
    0.01662077, -5.319421e-07, 0, 4.553267e-07, 0.01427187, 0.05661352, 
    0.03530488, 0.005725941, 0.0001533268,
  -1.1276e-07, 0.001660354, 0.0003064132, 0.000366708, 0.0005119881, 
    0.000225199, -3.164955e-08, 0.00780958, 0.01031077, -2.446113e-06, 
    4.120563e-05, -3.251098e-08, 0.00251812, 3.772644e-05, -1.830063e-05, 
    0.01075582, 0.05245616, 0.06876934, 0.008758451, 0.0009277293, 
    -2.715187e-05, 3.537678e-05, 0, 0.000166874, 0.02535472, 0.01866102, 
    0.01180346, -4.696924e-06, -1.309037e-05,
  0, 0.02949271, 0.01229211, -4.213419e-05, 0.003243825, 0.07100136, 
    0.02413167, 0.09442416, 0.02156917, 9.931585e-06, 0.01355051, 0.07757837, 
    0.02670019, 0.04841874, 0.1320473, 0.04909096, 0.03023832, -2.185309e-05, 
    -7.217355e-07, 0, -1.567245e-10, -5.949779e-07, 3.957066e-05, 0.2052855, 
    0.1418049, 0.007211671, 1.547654e-05, 0, -1.278989e-07,
  -8.485094e-10, 0.09194311, 0.05999139, 0, -7.3064e-09, 0.04758409, 
    0.001153392, 0.04512209, 0.06528322, 0.05261386, 0.0009981802, 
    0.09322871, 0.1215027, 0.2014492, 0.04698726, 5.438025e-05, 3.336598e-05, 
    -0.0001051591, -2.997868e-06, 0.0001184666, 1.143992e-06, 6.225261e-05, 
    0.02550719, 0.2304257, 0.07347336, 0.009737259, 0.01814046, 1.691122e-07, 
    -6.724896e-07,
  0.0004905983, -9.686921e-05, -4.968012e-06, 0.000503319, 8.261847e-05, 
    2.651197e-09, 0.06964126, 0.1603224, 0.1686388, 0.1589069, 0.2186466, 
    0.2720225, 0.4236994, 0.3014146, 0.2376446, 0.1369395, 0.2127742, 
    0.06976223, 0.03681867, 0.09403976, 0.0851391, 0.1649306, 0.0702227, 
    0.05895206, 0.02318319, 0.02985364, 0.02535589, 0.007759154, -5.462295e-05,
  -4.383742e-07, -1.716865e-05, 0, -6.205171e-07, -3.719626e-11, 0.007399481, 
    0.05654343, 0.159736, 0.02609134, 0.02928416, 0.09005112, 0.1244955, 
    0.1107623, 0.1496668, 0.01714632, 0.01373855, 0.007022335, 0.03141202, 
    0.0003387951, 0.0008753044, 0.003285303, 0.07282893, 0.01536338, 
    0.03080897, 0.0007108612, 0.00349802, -9.937712e-05, 0.0003461035, 
    -7.563776e-06,
  0, 0, -1.81308e-07, 0.003709778, -4.609257e-07, -4.112353e-10, 
    -6.503374e-07, 0.003152585, 0.03440388, 0.008017479, 0.03994943, 
    0.05246557, 0.04466068, 0.0172014, 0.02721354, 0.002384073, 0.007390792, 
    0.008621718, 0.02187754, -1.742964e-05, 0.007096923, 0.006439754, 
    0.01684234, 0.005207628, 0.02234242, 0.006515031, 0.01200728, 
    8.505758e-05, 0,
  0.003911513, 0, 0.0004809198, 0, -6.741942e-08, -3.399953e-09, 
    -2.924531e-10, 0, 0, -5.900817e-06, 0.02025783, 0.04357406, 0.09701203, 
    0.1030939, 0.03489878, 0.02774544, 0.02878464, 0.02886847, 0.0007584855, 
    0, 0, 0.001872321, 0.03043539, 0.02958051, 0.02230191, 0.04933501, 
    0.02718132, 0.02058735, 0,
  0.003531431, 0.0005605638, 2.823264e-05, 0.004108857, -4.847128e-05, 0, 0, 
    0, 0, 0, 0, 0.005495994, 0.01259843, 0.01229167, 0.01933306, 0.01584677, 
    0.0275541, 0.03563698, 0.003253573, -5.119536e-05, 0, 0.003968893, 
    -0.0001942869, 0.001238638, 0.007444961, 0.007148067, 0.0358158, 
    0.005543408, -8.859659e-06,
  0, -1.096244e-05, 0, 0, 0, -5.014283e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -1.165118e-05, 0.002649982, -3.038479e-06, 0.01111107, -0.0003572826, 
    -2.553986e-05, 0, 0.001924011, -0.0001381656, 0.005800363, 0.000560764, 
    0.0005432118, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0004480206, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0.001799606, 0, 0, 0, 0, 0, 0, 0, 0.0002064422, 0, 0, 0, 
    0, 0, 0, 0.0007298733, 0, 0, 0, 0, 0, 0, 0,
  0.0001006163, 0.002174684, 0.004609591, 0.005165121, 0.004829434, 
    0.00516913, 0.007571718, 0.007775912, 0.0001921256, 0.0001471189, 0, 
    0.0001217374, 0.0003374785, 0.003364711, -6.740001e-06, 0, -1.794593e-05, 
    -5.643565e-06, 0.000254272, 0.0010399, 0.0009184208, -4.956464e-06, 
    -4.363437e-05, -3.431295e-09, -3.417363e-05, -9.094922e-06, 0.003759528, 
    -2.22003e-06, -7.117846e-06,
  0.02378346, 0.007918399, 0.005133996, 0.006803001, 0.03601332, 0.01148791, 
    0.01247817, 0.001678653, -3.56708e-10, -4.175118e-09, 0.0008696076, 0, 
    0.007620217, 0.01346507, 0.02673238, 0.006918254, 0.01746492, 
    0.005062591, 0.01038808, 0.01400033, 0.02279788, 0.002642798, 
    -1.155189e-05, 0, 0.03180861, 0.004534924, 0.02081948, 0.02642961, 
    0.02074911,
  0.0001824101, 0.0001463217, 5.589573e-05, 0.0970408, 0.04369834, 
    0.002942545, 0.0004109133, 0.001029137, 0.002421252, 4.100922e-05, 
    0.01621928, 0.01987606, 0.001905552, 0.003311486, 0.04978134, 0.03094292, 
    0.009393373, 0.0345809, 0.09256975, 0.06049248, 0.03600198, 0.001039319, 
    9.570043e-05, 0.007978201, 0.04261851, 0.1040095, 0.1161948, 0.06264427, 
    0.01829171,
  0.000191614, 0.0468904, 0.03221053, 0.04949001, 0.01816219, 0.03287987, 
    0.0001966943, 0.009479143, 0.026935, -1.659743e-05, 0.0001246899, 
    9.58772e-06, 0.002654936, 0.0002828739, 0.0006872463, 0.07514383, 
    0.1712139, 0.2192048, 0.1169984, 0.03374196, 0.01450357, 0.00711095, 
    3.912728e-06, 0.04010677, 0.1111662, 0.09444538, 0.0858488, 0.04372906, 
    0.001576255,
  9.416582e-08, 0.05056103, 0.2287162, 0.01301783, 0.03877547, 0.133305, 
    0.05597209, 0.1380875, 0.02514617, 0.0005156428, 0.00957287, 0.05537516, 
    0.01393646, 0.05436548, 0.1279082, 0.0630713, 0.1099703, 0.001603946, 
    1.40029e-07, 1.465646e-07, 1.966313e-06, 3.852537e-05, 0.007335315, 
    0.3943837, 0.218076, 0.05574618, 0.06573229, 0.0007614273, 3.278907e-05,
  1.591543e-05, 0.270867, 0.3885777, 0.000564927, 2.943838e-05, 0.06034099, 
    0.01798019, 0.07266454, 0.3358553, 0.325299, 0.01624019, 0.08005993, 
    0.1578462, 0.2075554, 0.03401268, 0.0001529609, 0.0006837865, 
    0.0006483903, -1.611361e-06, 0.00460792, 0.0001320267, 0.04748439, 
    0.112358, 0.3760286, 0.08634272, 0.01198652, 0.03854909, 0.00500226, 
    0.0008935269,
  0.1217204, 0.06051777, -0.0001748197, 0.00157382, 0.0001833302, 
    2.117318e-05, 0.1621259, 0.1750849, 0.2093053, 0.1232622, 0.2040216, 
    0.2150357, 0.3663673, 0.286806, 0.2262373, 0.1797275, 0.2746377, 
    0.1232161, 0.08005078, 0.1189445, 0.1006688, 0.1896784, 0.3279303, 
    0.1450806, 0.1086275, 0.2087191, 0.2479872, 0.165877, 0.01378896,
  0.006999836, 0.008758602, 0.0001819878, 0.0008632446, -9.311454e-08, 
    0.01395931, 0.04621286, 0.1721903, 0.04148937, 0.02846241, 0.07883271, 
    0.0942205, 0.09626538, 0.1501236, 0.0420569, 0.08045133, 0.1049638, 
    0.1243424, 0.04388051, 0.004961124, 0.09526689, 0.06929318, 0.04872877, 
    0.06051026, 0.0681686, 0.04469809, 0.05070636, 0.301007, 0.03747526,
  -4.283475e-06, 0.001115133, 4.461514e-05, 0.00500916, 0.0004700032, 
    2.872613e-05, 0.0001842282, 0.0098714, 0.04781799, 0.06732737, 
    0.06567113, 0.1125691, 0.0885085, 0.04950728, 0.0777214, 0.05523032, 
    0.06850837, 0.02154245, 0.04816797, 0.01848799, 0.008765541, 0.03045309, 
    0.04346182, 0.07386176, 0.1656725, 0.09281863, 0.05294923, 0.004539375, 
    0.0004697072,
  0.007054644, 0.0001143797, 0.001755969, -4.008443e-06, -1.081598e-05, 
    0.0006311886, -1.078321e-07, 0, -7.762861e-07, -3.260913e-05, 0.03759184, 
    0.07961337, 0.1480999, 0.2035287, 0.1101584, 0.07982409, 0.05905485, 
    0.05582519, 0.01508867, -6.213311e-06, 0, 0.004424356, 0.04102419, 
    0.05697466, 0.05897229, 0.1196948, 0.04893299, 0.03101421, -2.55017e-07,
  0.006235218, 0.003232808, 6.268118e-05, 0.007940108, 0.0003573805, 
    0.001729612, 0, 0, 0, 0, -4.819031e-06, 0.01204547, 0.02436775, 
    0.03613684, 0.02402789, 0.01999608, 0.04220076, 0.07703342, 0.0178889, 
    -0.000201001, 3.06095e-05, 0.01208411, 0.003687483, 0.009755986, 
    0.01525475, 0.01826997, 0.09044616, 0.01019572, 0.0109928,
  4.039525e-05, 0.0001280318, 0.0002450795, 0, 0, 0.000137539, 0.0001651777, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1.38094e-05, 0.01760036, 0.004265619, 
    0.01947739, 0.001187339, 5.662968e-05, 0, 0.007666306, 0.004346552, 
    0.02146255, 0.01090096, 0.006397672, 0.002897858,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7.204133e-06, 
    -1.164383e-05, 1.837079e-07, -1.134561e-05, 0.001421411, 0.0004321802, 
    -7.8131e-08, 0, 0, 0, -1.109948e-06, 0.001434061, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0007280041, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1.840192e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0, -1.788559e-11, 0.002451596, 0, 0, 0, 0, 0, -4.917691e-05, 
    1.411432e-05, 0.00297007, 0.0001485945, 0, 8.865131e-05, 0, 0, 0, 
    0.001478694, 0, 0, 0, 0, 0, 0, 0,
  0.00456104, 0.006506867, 0.0101271, 0.02211303, 0.01392127, 0.01604474, 
    0.01555339, 0.01498711, 0.006486205, 0.01305672, 0.003565936, 
    0.003797037, 0.0003789031, 0.006497168, 0.002246143, 2.368806e-05, 
    1.315313e-05, 0.006726052, 0.00301932, 0.007880202, 0.01201881, 
    0.003155533, 0.00313337, -4.589084e-05, 0.002330763, -7.372138e-05, 
    0.005921393, -0.0002750778, 0.002285475,
  0.05420724, 0.015779, 0.04866266, 0.03872624, 0.09401955, 0.08410624, 
    0.04372097, 0.02386211, 0.007065884, 0.001045606, 0.01076607, 
    -2.324025e-05, 0.01711946, 0.0211215, 0.05759694, 0.02168174, 0.03038542, 
    0.01226499, 0.01933756, 0.02854446, 0.04136532, 0.02086676, 0.002229738, 
    -4.973554e-05, 0.04306509, 0.03424243, 0.05530802, 0.03880515, 0.04445639,
  0.03668369, 0.007657594, 0.03070738, 0.1285632, 0.1059031, 0.09572364, 
    0.01757864, 0.0304342, 0.02271166, 0.02115564, 0.02144371, 0.04403098, 
    0.01318636, 0.01982475, 0.07596957, 0.1076996, 0.05661809, 0.1013327, 
    0.2609794, 0.1595916, 0.1192778, 0.04978166, 0.02902226, 0.0397865, 
    0.05657412, 0.1354745, 0.1623589, 0.175189, 0.1164905,
  0.0001138741, 0.04133168, 0.1291479, 0.03125275, 0.08079327, 0.01458532, 
    0.002880363, 0.001207554, 0.02987951, 2.255101e-05, 0.006572049, 
    0.001805091, 0.000269743, 0.000234968, 0.00843078, 0.08487747, 0.1761494, 
    0.2390752, 0.1506229, 0.04969823, 0.03114989, 0.01729594, 9.017844e-07, 
    0.03976839, 0.08293128, 0.08889783, 0.08406149, 0.02051243, -6.939028e-05,
  -1.402053e-11, 0.03149222, 0.1360828, 0.008498746, 0.02698983, 0.08997505, 
    0.04142607, 0.1204594, 0.02335807, 0.000373984, 0.0004129533, 0.03797372, 
    0.005691804, 0.02191983, 0.1058782, 0.04865083, 0.08284979, 0.003440732, 
    1.775166e-08, 3.768521e-07, 1.229938e-07, 1.050817e-06, 0.0001479427, 
    0.3412625, 0.1833276, 0.02858535, 0.06839985, 0.001620279, 1.756602e-07,
  2.59395e-05, 0.1956719, 0.320356, 0.0003140013, -1.498327e-06, 0.05510618, 
    0.009169782, 0.05230152, 0.2376821, 0.2165737, 0.02168904, 0.06870412, 
    0.08578407, 0.1524805, 0.02339917, 0.0009619007, 3.433223e-05, 
    -1.005981e-05, 5.896854e-07, 0.0002633302, 1.563902e-05, 0.006461319, 
    0.07410096, 0.3578814, 0.05210987, 0.001310284, 0.03456409, 0.001123284, 
    3.649081e-05,
  0.07737834, 0.03570789, 0.0001025928, 0.03977089, 0.0004763179, 
    1.737715e-05, 0.1133168, 0.1277247, 0.1765808, 0.0783428, 0.164719, 
    0.1782073, 0.3054982, 0.2767681, 0.1776739, 0.1324032, 0.2294589, 
    0.09767376, 0.04193247, 0.1086068, 0.08767188, 0.1108547, 0.2473835, 
    0.1179618, 0.06525653, 0.1706873, 0.1662602, 0.1254263, 0.006636765,
  0.009353552, 0.004413316, 7.684859e-05, 0.001015114, -8.826564e-09, 
    0.004919433, 0.03780653, 0.1399496, 0.04626734, 0.03142713, 0.07231192, 
    0.07911267, 0.07092191, 0.1241955, 0.0139996, 0.04276323, 0.1114955, 
    0.1064411, 0.04431351, 0.01345519, 0.09146737, 0.05978271, 0.02973335, 
    0.0367906, 0.04281035, 0.04448223, 0.04858358, 0.3742795, 0.1032777,
  0.05988692, 0.02167158, 0.01318723, 0.01396726, 0.006689719, 0.003720973, 
    0.003584133, 0.0185687, 0.06955095, 0.09406328, 0.07565979, 0.08390133, 
    0.07657494, 0.01684074, 0.04663849, 0.06287616, 0.06554078, 0.04960364, 
    0.08052508, 0.04943403, 0.01629552, 0.07644732, 0.09699454, 0.08135816, 
    0.1673217, 0.09910086, 0.1083184, 0.07619213, 0.0994793,
  0.05222688, 0.02142769, 0.005918496, -1.105118e-05, 0.006351036, 
    0.005263766, 3.254126e-06, 4.419328e-05, 0.0003133832, 1.858853e-05, 
    0.07992496, 0.1300806, 0.2125474, 0.2376753, 0.1605004, 0.1285681, 
    0.111351, 0.1653075, 0.1140399, 0.0003864789, -1.509418e-05, 0.008771398, 
    0.04696976, 0.07225399, 0.1278911, 0.2146133, 0.1396925, 0.04943858, 
    0.03456806,
  0.05006341, 0.01113201, 0.000420716, 0.0117567, 0.002246393, 0.003186058, 
    0, 0, 0, 0, -0.0001010609, 0.03105075, 0.04218477, 0.0432853, 0.06535995, 
    0.05166406, 0.1061014, 0.1953017, 0.208912, 0.008807913, 0.00104898, 
    0.01806752, 0.02980373, 0.0307788, 0.04586345, 0.09036951, 0.1820305, 
    0.1152386, 0.07444257,
  0.01842404, 0.003619334, 0.004310453, 9.422679e-05, 0, 0.0001901686, 
    0.002054604, 0, 0, 0, 0, 0, 0, -6.115663e-08, 6.98116e-06, 2.321374e-05, 
    0.001199174, 0.06667395, 0.01518004, 0.04656151, 0.01545703, 0.009368429, 
    -4.240868e-05, 0.01405187, 0.02482606, 0.06328735, 0.06297109, 
    0.06541657, 0.04857432,
  -2.837016e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0003888744, 
    -0.0002483814, 0.01084617, 0.007559247, 0.01051029, 0.006737224, 
    0.0002739481, 0.001699827, -1.292951e-05, -4.307643e-06, 1.029141e-06, 
    0.006176839, 0.0009700849,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002003158, 0, 0, 0, 0, 0, 
    -1.363565e-05, 0, 0, 0, 0.000359139, 0, 0, 0, 0,
  0, 0, -1.383309e-06, 0, 0, 0.0001769311, 0.006083008, -3.968853e-05, 0, 0, 
    0, 0, 0.001178102, 0.0009402864, 0.00769352, 0.003546271, -2.78211e-06, 
    0.0003477959, 0, 0, 0, 0.003298854, 0, 2.913001e-05, -4.12987e-06, 0, 
    2.898972e-08, -1.312023e-05, 0,
  0.02636077, 0.0399631, 0.04113157, 0.06232073, 0.07337388, 0.07179458, 
    0.06754769, 0.1058377, 0.1017433, 0.07240292, 0.02801601, 0.03770777, 
    0.03111943, 0.05360368, 0.04077698, 0.02256809, 0.02891196, 0.05688754, 
    0.03499597, 0.03082472, 0.0363907, 0.00940329, 0.01666983, 0.008094239, 
    0.002431492, 0.003208708, 0.01248728, 0.01524141, 0.02763294,
  0.1119758, 0.0826208, 0.07584816, 0.08270685, 0.1241414, 0.1047863, 
    0.1045556, 0.1106146, 0.0748262, 0.06764974, 0.06642236, 0.02938421, 
    0.04427749, 0.07707357, 0.09504514, 0.1401345, 0.1811807, 0.0974528, 
    0.1223684, 0.1022979, 0.10706, 0.06448281, 0.01772566, 0.004997071, 
    0.07938882, 0.05452925, 0.1200578, 0.1047407, 0.09923367,
  0.03152845, 0.01064323, 0.09015114, 0.1248937, 0.1049205, 0.08323646, 
    0.004901241, 0.01568327, 0.01774183, 0.01908243, 0.03148856, 0.07703623, 
    0.06298903, 0.08378953, 0.1195622, 0.1424035, 0.0750154, 0.09397385, 
    0.2651681, 0.1807373, 0.1262393, 0.07851078, 0.02268328, 0.05144204, 
    0.04894688, 0.1177004, 0.1660677, 0.1747421, 0.1210613,
  3.180906e-05, 0.02795715, 0.1047279, 0.009445644, 0.05407502, 0.01695797, 
    0.0004483018, 0.0001230688, 0.03991782, 0.001991361, 0.008969606, 
    0.004137937, 7.65042e-06, 0.003559092, 0.01733039, 0.08053179, 0.1905098, 
    0.2160279, 0.06515928, 0.0244472, 0.006361158, 0.005724774, -9.62243e-08, 
    0.0354871, 0.06358757, 0.08383017, 0.07926795, 0.007412255, 3.186281e-06,
  0, 0.02777018, 0.08295961, 0.002057907, 0.01936167, 0.06545676, 0.03639493, 
    0.1099594, 0.03159796, 0.00138166, 1.837093e-05, 0.02803795, 0.005232876, 
    0.02201635, 0.08683727, 0.0507137, 0.07414206, 0.003466093, 3.603886e-09, 
    1.554868e-07, 2.623312e-08, 4.370926e-07, 1.710446e-05, 0.2969496, 
    0.1852311, 0.02803, 0.03281394, 0.0004677578, 3.046938e-08,
  0.0001348183, 0.1679572, 0.2768768, 0.0001216459, 7.714977e-06, 0.05637883, 
    0.008215227, 0.04593811, 0.1644865, 0.161783, 0.0156535, 0.04435404, 
    0.05841282, 0.1433464, 0.02288333, 0.0003945172, -1.600735e-06, 
    1.821717e-06, 3.486602e-07, -2.604348e-05, 2.617883e-06, 9.764433e-05, 
    0.03381383, 0.3154731, 0.0373809, -3.580935e-05, 0.02756697, 
    2.411175e-05, 7.852236e-06,
  0.05917333, 0.02560893, 0.000510433, 0.02743059, 0.0003038295, 
    8.809056e-06, 0.0922317, 0.1127433, 0.1520141, 0.0611038, 0.113005, 
    0.156233, 0.2570269, 0.2880999, 0.144912, 0.105742, 0.215132, 0.09465175, 
    0.03130077, 0.1040718, 0.08290295, 0.08492255, 0.2023715, 0.09555857, 
    0.03881434, 0.1381332, 0.1297565, 0.08212386, 0.005012155,
  0.003525082, 0.007244152, 2.777124e-05, 0.001131625, -3.705429e-09, 
    0.0009266157, 0.03454635, 0.1274025, 0.04136983, 0.03099966, 0.07467797, 
    0.06634156, 0.06916463, 0.1062475, 0.01205337, 0.03644722, 0.08876726, 
    0.06749274, 0.02750438, 0.01967335, 0.08235446, 0.05221664, 0.01763396, 
    0.02724961, 0.02967966, 0.04379766, 0.03508896, 0.2978373, 0.06749696,
  0.09821109, 0.03533429, 0.01115517, 0.0253502, 0.01131523, 0.0005778802, 
    0.003586996, 0.02883002, 0.1152491, 0.1083273, 0.07535738, 0.05733858, 
    0.06312337, 0.002231787, 0.04240247, 0.05241847, 0.06622689, 0.05907992, 
    0.08765762, 0.04995822, 0.04263274, 0.05351738, 0.07642497, 0.06585027, 
    0.1363288, 0.08049347, 0.09256428, 0.06621034, 0.1247204,
  0.1377696, 0.06489813, 0.05353562, 0.006270223, 0.02824133, 0.04519469, 
    4.02378e-05, 0.001144849, 0.01175172, 0.002185457, 0.1341538, 0.1617611, 
    0.2354272, 0.1973108, 0.1539357, 0.1725631, 0.1473586, 0.2545773, 
    0.115422, 0.01972727, 0.0008479956, 0.055148, 0.08764505, 0.08994181, 
    0.1418945, 0.2245536, 0.1298423, 0.07828658, 0.07387062,
  0.1192362, 0.08052746, 0.01975577, 0.04623108, 0.06615718, 0.03765043, 
    0.0006979383, -6.113022e-06, 4.843637e-06, -2.858872e-05, 0.0004611191, 
    0.05528908, 0.0726651, 0.05899953, 0.09440129, 0.09450885, 0.1157663, 
    0.266361, 0.3268695, 0.05604974, 0.02495958, 0.08278386, 0.08682646, 
    0.06697933, 0.0895616, 0.148595, 0.2422019, 0.1646211, 0.1069801,
  0.09341859, 0.01918575, 0.01139759, 0.01372221, 0.001434501, 0.01502263, 
    0.01565724, 0.002633665, -9.335099e-06, -3.925658e-05, -4.212481e-05, 0, 
    -2.043851e-05, -0.0001181517, 0.009187536, 0.007026934, 0.01465808, 
    0.1349395, 0.04756612, 0.06594206, 0.03078557, 0.06040969, 0.02074583, 
    0.03489178, 0.05790488, 0.09796197, 0.1237684, 0.08156776, 0.1333738,
  0.001092972, 0.007080099, -1.397999e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.0008508965, 0.01114834, 0.05075917, 0.09289874, 0.06522723, 
    0.03598085, 0.01338488, 0.006185225, 7.258009e-05, -4.416251e-05, 
    -7.056793e-07, 0.03120861, 0.01445699,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -6.170274e-07, 
    9.137936e-05, -7.066476e-07, 0, 2.569558e-07, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0007374954, 0.004163043, 0, 
    -2.174443e-05, -0.0002082272, 8.540343e-06, 0, 0.001907988, 3.660139e-05, 
    2.495401e-06, 0.0007887751, 0.009519418, -4.528335e-06, -3.876038e-06, 0, 0,
  0.009191852, 0.003813892, 6.066777e-06, 0, -9.308899e-06, 0.007669826, 
    0.01104866, 0.001340175, 0.001129857, -2.162168e-05, 2.386376e-05, 
    0.009557187, 0.005864715, 0.01538667, 0.03631802, 0.03826871, 0.04447769, 
    0.06205594, 0.03826012, 0.01859015, 0.003784706, 0.02304724, 0.03352293, 
    0.02034697, 0.005713972, 0.005286315, 0.00769091, 0.003662601, 0.01252992,
  0.109147, 0.1132733, 0.1165149, 0.1699093, 0.1269038, 0.1440784, 0.1147228, 
    0.1646939, 0.1603664, 0.1486019, 0.1271298, 0.109558, 0.08583091, 
    0.1046688, 0.1009153, 0.1872873, 0.1231621, 0.1219083, 0.1054089, 
    0.1251944, 0.1370929, 0.1168362, 0.06828523, 0.02076479, 0.05634325, 
    0.05823798, 0.08744957, 0.1621506, 0.1198356,
  0.1610761, 0.1140161, 0.08572471, 0.08680924, 0.1141266, 0.1004143, 
    0.1097257, 0.1333929, 0.1125794, 0.142265, 0.0963162, 0.03625049, 
    0.09785084, 0.1206974, 0.1691868, 0.1617333, 0.1994384, 0.1425924, 
    0.1185695, 0.1019954, 0.1278094, 0.0889893, 0.05131204, 0.01904463, 
    0.08699054, 0.1056462, 0.1576847, 0.1261962, 0.130651,
  0.02368961, 0.003778354, 0.07731564, 0.1182681, 0.09472418, 0.05321961, 
    0.00565067, 0.001659525, 0.01550028, 0.02922658, 0.03903881, 0.05674636, 
    0.07855166, 0.07265516, 0.1288083, 0.0737718, 0.03982197, 0.05446181, 
    0.2585607, 0.1796973, 0.1279771, 0.05660626, 0.03182374, 0.01933216, 
    0.03833137, 0.09795014, 0.1463808, 0.143, 0.1183963,
  1.81169e-05, 0.01599306, 0.07580455, 0.001979512, 0.01519225, 0.0173516, 
    -7.024324e-06, -0.001382195, 0.03831091, 0.01359162, 0.005429343, 
    0.0008962614, 6.396307e-07, 0.008058355, 0.03127582, 0.08357079, 
    0.1900922, 0.1738909, 0.04162433, 0.007839141, 0.0002799986, 0.001618396, 
    -1.573888e-09, 0.01536798, 0.05646125, 0.09119466, 0.08366503, 
    0.005385475, 1.220154e-05,
  -1.194641e-09, 0.03008184, 0.06565629, 0.001101444, 0.01157471, 0.0423816, 
    0.03530375, 0.1015103, 0.04132578, 0.001357582, 0.0001120932, 0.02096532, 
    0.005828436, 0.01716692, 0.06221381, 0.06493554, 0.06837269, 
    0.0001279524, 1.012842e-08, 1.229568e-08, 3.737938e-09, 1.823782e-07, 
    3.325999e-06, 0.2380975, 0.1490977, 0.02687437, 0.002259425, 
    0.0002511466, -1.139493e-10,
  1.086145e-05, 0.1419664, 0.1922184, 0.0001015173, 1.056511e-05, 0.05347596, 
    0.009914698, 0.04157034, 0.1000251, 0.09546708, 0.01296161, 0.030693, 
    0.05408096, 0.1160457, 0.02942438, 0.0001062854, -7.242531e-05, 
    9.07086e-07, -5.488692e-07, -4.2425e-06, 2.092541e-06, 1.519714e-05, 
    0.01304746, 0.2397299, 0.02319663, -2.865278e-06, 0.02443896, 
    9.602829e-05, 1.135299e-06,
  0.04140751, 0.02386522, 0.002407335, 0.009457403, 0.0005392884, 
    2.893547e-06, 0.07084575, 0.1094701, 0.143505, 0.04566309, 0.08016676, 
    0.1423544, 0.2227779, 0.2887893, 0.1221512, 0.07964513, 0.2268404, 
    0.08575817, 0.02861294, 0.09437264, 0.07774147, 0.05732238, 0.1621745, 
    0.06731769, 0.02838698, 0.1397597, 0.114241, 0.05337858, 0.005462027,
  0.002799104, 0.004193853, 1.080684e-05, 0.002081752, 1.047666e-07, 
    0.0001708939, 0.03321635, 0.1143544, 0.06477325, 0.03233381, 0.07283462, 
    0.06007617, 0.05953358, 0.08850269, 0.009432484, 0.02733902, 0.05785656, 
    0.04941895, 0.01326466, 0.01784129, 0.06669364, 0.04315266, 0.01703511, 
    0.02376492, 0.02084296, 0.04094203, 0.05328591, 0.2428978, 0.04347613,
  0.09725615, 0.0515143, 0.00524577, 0.01499595, 0.007273806, 7.359453e-05, 
    0.007926916, 0.03406873, 0.1629174, 0.1241597, 0.08043792, 0.0538503, 
    0.05431313, 0.001787277, 0.02344701, 0.05254095, 0.06760824, 0.06098782, 
    0.05816324, 0.04683817, 0.03952165, 0.03526329, 0.05559137, 0.03998876, 
    0.1108148, 0.05786216, 0.08316531, 0.05414543, 0.08827936,
  0.1681683, 0.06215193, 0.04824383, 0.02359211, 0.0373701, 0.05873078, 
    0.003574949, 0.06316578, 0.05469215, 0.04236923, 0.1393711, 0.1662404, 
    0.2480533, 0.1761964, 0.1377547, 0.1747608, 0.1733217, 0.2525104, 
    0.1052513, 0.01924508, 0.03834609, 0.09544644, 0.09682921, 0.08405805, 
    0.1358598, 0.1836534, 0.1295057, 0.0815279, 0.09073637,
  0.1311083, 0.1107258, 0.07659382, 0.1194823, 0.1349735, 0.09314818, 
    0.06060586, -6.072355e-05, -8.915771e-06, 0.001686278, 0.01579093, 
    0.09572782, 0.1195493, 0.05754588, 0.1017681, 0.1500691, 0.126465, 
    0.3042509, 0.3568417, 0.1218099, 0.06999616, 0.1165986, 0.09936894, 
    0.1459189, 0.1137134, 0.1734775, 0.2543968, 0.148811, 0.1043887,
  0.1885464, 0.08807359, 0.04702957, 0.0601485, 0.08594857, 0.09874081, 
    0.1035402, 0.05835646, 0.01461914, 0.007007981, -4.624878e-05, 0, 
    0.001321798, 0.0246448, 0.01473085, 0.04546076, 0.05344594, 0.155879, 
    0.06978329, 0.120837, 0.1101839, 0.1262269, 0.04288626, 0.08943376, 
    0.1486786, 0.1648779, 0.1808269, 0.1358691, 0.1833685,
  0.05393478, 0.01986108, -4.025161e-05, -7.352057e-06, -0.0001147387, 
    0.003229977, 0.002783997, -3.21912e-05, -1.635282e-07, 5.353124e-05, 
    1.061193e-07, 0, 0, 0, 1.407003e-07, 1.109193e-05, 0.0187369, 0.09093107, 
    0.116962, 0.1530554, 0.09873177, 0.1015703, 0.0596629, 0.01699885, 
    0.03707927, 0.0002242646, -0.0003355829, 0.1187676, 0.06706848,
  0, 0, 0, 0.0002682486, 0.0004605373, 0, 0, 0, -1.47016e-06, 9.260197e-07, 
    0, 0, 0, 0, -1.422386e-05, 0.00319756, 0.02695601, 0.03416907, 
    0.01008954, 0.001309248, 0.0004204881, 0.001748217, 0.0001484745, 
    -2.212997e-05, -7.851731e-09, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -4.40426e-05, 
    0.0002364608, 0, 0, 0, 0, 0.0001908041, 0.003737278, -0.0001675464, 0, 0, 0,
  4.323616e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.134533e-05, 0.001962798, 
    0.006419137, -3.644883e-05, 0.003100642, 0.004850817, 0.0002028553, 
    0.0003728259, 0.01353971, 0.02370333, 0.02503404, 0.02423561, 0.04526296, 
    0.01236641, 0.00572418, 0.0001748696, 0,
  0.07025171, 0.0792797, 0.08600365, 0.04443674, 0.01111893, 0.02803704, 
    0.05889175, 0.04210806, 0.04148051, 0.02362179, 0.03606487, 0.04897042, 
    0.05970653, 0.09151775, 0.1022933, 0.1123134, 0.07059253, 0.1032352, 
    0.1103148, 0.1059111, 0.09724496, 0.1089272, 0.09174255, 0.07824635, 
    0.05153935, 0.06334563, 0.06570484, 0.05264135, 0.06380538,
  0.1685397, 0.148687, 0.1656748, 0.209044, 0.1493178, 0.1620185, 0.1451097, 
    0.185466, 0.2018102, 0.2073667, 0.1603939, 0.1165212, 0.1267302, 
    0.1390857, 0.1472628, 0.2002224, 0.1493673, 0.1273721, 0.1339278, 
    0.1750347, 0.1784069, 0.1668993, 0.1454532, 0.08554778, 0.108282, 
    0.1617208, 0.2037816, 0.2542513, 0.1739873,
  0.1524419, 0.1040673, 0.07548694, 0.08298076, 0.1045547, 0.1007117, 
    0.1126923, 0.1086134, 0.1183976, 0.137396, 0.06625151, 0.03232882, 
    0.09140154, 0.1055854, 0.1731662, 0.1475125, 0.1812402, 0.1214694, 
    0.1170175, 0.09265626, 0.1101878, 0.08731406, 0.06023121, 0.04313483, 
    0.0912283, 0.1103643, 0.1673645, 0.1256627, 0.1332467,
  0.02671978, 0.002082209, 0.0629841, 0.1056792, 0.08386146, 0.03925899, 
    0.004227637, 0.001001996, 0.01737743, 0.009356146, 0.04225087, 
    0.04484102, 0.09741741, 0.07023068, 0.1264544, 0.05151694, 0.02805541, 
    0.04206452, 0.2643664, 0.17793, 0.1055229, 0.03553263, 0.02681185, 
    0.01012941, 0.03444608, 0.08585427, 0.1260104, 0.123487, 0.1317689,
  1.032501e-05, 0.01027627, 0.04755046, 0.0009374661, 0.006419282, 
    0.01265289, 0.001370093, -0.001113149, 0.05464387, 0.009601051, 
    0.007568517, 2.186718e-05, -2.826385e-07, 0.01442486, 0.05071782, 
    0.09805264, 0.1970697, 0.1657642, 0.03240441, 0.005414291, 2.268344e-05, 
    -1.770502e-05, -7.625165e-12, 0.007085792, 0.04719579, 0.1032447, 
    0.06239678, 0.00228559, 3.484003e-05,
  -1.573317e-07, 0.03545354, 0.04503253, 0.0009994518, 0.007074064, 
    0.03506682, 0.02936515, 0.09317954, 0.03587704, 0.0006469859, 
    0.0002207369, 0.01276511, 0.01929282, 0.01546714, 0.04307097, 0.09491481, 
    0.05984536, 6.829338e-05, 8.586283e-10, 8.102935e-09, -7.105652e-11, 
    1.236166e-07, 7.703012e-06, 0.1836838, 0.1122276, 0.01469071, 
    0.0006759361, 1.593363e-05, -9.238762e-11,
  0.0004239857, 0.1551874, 0.1325272, 0.001460988, 0.0003834021, 0.04963975, 
    0.01917851, 0.04308546, 0.06353828, 0.05640431, 0.007134062, 0.0174362, 
    0.04413659, 0.0805103, 0.01915153, 0.0003190857, 0.001230674, 
    3.899077e-07, 1.852483e-05, 2.188304e-06, 5.967121e-07, 5.798036e-06, 
    0.000618586, 0.1718034, 0.01725346, 0.0002360628, 0.02100574, 
    1.261732e-05, 4.575808e-07,
  0.03053917, 0.0228578, 0.00359082, 0.005533997, 0.0006722239, 7.179335e-06, 
    0.05056909, 0.08908961, 0.1251952, 0.03393914, 0.06283872, 0.1244304, 
    0.1800894, 0.2912635, 0.1002831, 0.0657207, 0.217613, 0.07601248, 
    0.03389423, 0.08435285, 0.08256785, 0.03908092, 0.1273495, 0.04845152, 
    0.03263722, 0.1399032, 0.1058732, 0.02921699, 0.008310432,
  0.003114675, 0.002849681, 3.217728e-06, 0.002453998, 4.713134e-08, 
    0.002331275, 0.03937598, 0.09392971, 0.06298028, 0.03196417, 0.06514934, 
    0.04593544, 0.05570226, 0.07376719, 0.005408589, 0.01603776, 0.02763561, 
    0.04345753, 0.01374502, 0.009873634, 0.04386188, 0.03501653, 0.01527588, 
    0.01654881, 0.01467938, 0.03178031, 0.0642827, 0.1995992, 0.02738532,
  0.1028544, 0.05087148, 0.002026669, 0.006420698, 0.003879592, 5.014105e-06, 
    0.005726291, 0.04283076, 0.2249688, 0.1153423, 0.08707838, 0.05160018, 
    0.05129988, 0.006849215, 0.009139509, 0.0370372, 0.07247189, 0.05100446, 
    0.0487283, 0.02951722, 0.03294006, 0.0300854, 0.04800259, 0.02774703, 
    0.09374207, 0.05410463, 0.08095702, 0.04286627, 0.06591823,
  0.1543924, 0.0521959, 0.03760688, 0.03249266, 0.03117449, 0.06064998, 
    0.009002999, 0.07884559, 0.06128749, 0.0678171, 0.125259, 0.1596137, 
    0.239626, 0.1711506, 0.1441478, 0.17163, 0.1729559, 0.2273857, 
    0.08938782, 0.01258556, 0.05755953, 0.09455113, 0.1012952, 0.0830813, 
    0.1238511, 0.1511893, 0.1355034, 0.07842749, 0.05758994,
  0.09973048, 0.1439876, 0.1860291, 0.1470838, 0.1391947, 0.1287838, 
    0.09116706, 0.02165937, 0.01154286, 0.03351659, 0.07749375, 0.1240745, 
    0.1611636, 0.0990519, 0.1616317, 0.2029696, 0.131155, 0.3083847, 
    0.3279614, 0.1178241, 0.1241893, 0.1074735, 0.09498799, 0.1636751, 
    0.1270781, 0.1587237, 0.2707202, 0.1360878, 0.09530034,
  0.2324043, 0.1418145, 0.1467254, 0.2321426, 0.1990589, 0.1810331, 
    0.2142221, 0.1944932, 0.1550468, 0.06735674, 0.0193692, 0.0005744787, 
    0.0108476, 0.04828754, 0.0206224, 0.07672221, 0.08073087, 0.1869344, 
    0.1475188, 0.1236971, 0.1454172, 0.1120859, 0.08132814, 0.1326432, 
    0.1568458, 0.1791843, 0.1758495, 0.1213611, 0.2339285,
  0.1435767, 0.1059352, 0.005565563, 0.01243917, 0.06068595, 0.1182322, 
    0.08419818, 0.06505315, 0.02611739, 0.009927811, 0.002326112, 
    -0.0002046666, -0.0004840897, 0.005228693, 0.04101017, 0.09099745, 
    0.1162948, 0.1876812, 0.1704915, 0.1677904, 0.1138592, 0.1378042, 
    0.1553768, 0.0876309, 0.1224895, 0.006523944, -0.001325798, 0.1959009, 
    0.1571634,
  0, -2.600708e-08, -0.0003312327, 0.02323729, 0.02477165, 0.03171593, 
    0.02885967, 0.0218159, 0.01930808, 0.04514899, -0.001368429, 
    0.0002060452, 0.004134642, -3.843086e-05, 0.00279104, 0.06716017, 
    0.1254548, 0.1129983, 0.07751599, 0.03003928, 0.02774446, 0.02814116, 
    0.009494253, -0.0008796001, 0.0001845951, 0, 0, -7.41226e-05, 2.584717e-06,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0003799961, 
    -0.0001404984, 0.002882567, -1.270157e-05, 0, 0, 0.0001055114, 
    0.001731475, 0.006969345, 0.004769879, 0.0009510076, -1.96135e-05, 0,
  0.006767104, 0.001099061, 1.796181e-06, -1.145576e-07, -7.94693e-06, 0, 
    -5.945516e-06, 0, 0, 0, 3.851092e-05, -4.022215e-06, 0.0001262012, 
    0.01213834, 0.01634032, 0.007614913, 0.0345685, 0.04201121, 0.02474432, 
    0.01256488, 0.0326786, 0.04830197, 0.06642262, 0.0813666, 0.06763247, 
    0.09292974, 0.1210766, 0.09597701, 0.04459343,
  0.2091318, 0.1630311, 0.2057506, 0.177501, 0.1116704, 0.1376709, 
    0.09922049, 0.07386151, 0.09933459, 0.08928189, 0.1106577, 0.1295205, 
    0.1040917, 0.1693854, 0.1661849, 0.1778386, 0.1548111, 0.1580889, 
    0.1508418, 0.1653116, 0.1549643, 0.1672806, 0.1466565, 0.1699765, 
    0.1614411, 0.131013, 0.1324462, 0.1685837, 0.1802049,
  0.1680109, 0.1358802, 0.1814598, 0.2219559, 0.1508144, 0.1451229, 
    0.1535451, 0.1862167, 0.2042782, 0.2117299, 0.1883332, 0.117082, 
    0.129348, 0.1606468, 0.1543417, 0.1775588, 0.141276, 0.1138831, 
    0.1261116, 0.176098, 0.1801392, 0.1664401, 0.1647684, 0.1383233, 
    0.1509434, 0.1625309, 0.2058087, 0.2648037, 0.2225419,
  0.154825, 0.1120265, 0.07407145, 0.08176647, 0.1037709, 0.1050718, 
    0.1086842, 0.101912, 0.0981961, 0.1155876, 0.0386858, 0.03006005, 
    0.08570933, 0.08827061, 0.1566156, 0.1313419, 0.1750393, 0.1094376, 
    0.1114191, 0.08532368, 0.08852911, 0.06982524, 0.06018075, 0.05280593, 
    0.0876492, 0.1050839, 0.161657, 0.1392898, 0.130094,
  0.03059154, 0.002191795, 0.05486417, 0.1021301, 0.07467675, 0.03554248, 
    0.006497335, 0.01166726, 0.01567762, 0.0001079022, 0.02607153, 
    0.05012934, 0.1048641, 0.06647434, 0.1356562, 0.03726664, 0.0333987, 
    0.04020135, 0.2789735, 0.1642234, 0.07962906, 0.02389592, 0.009164692, 
    0.007590056, 0.03569932, 0.07302007, 0.1195589, 0.1131953, 0.1266739,
  8.088756e-06, 0.009110575, 0.04530831, 0.0008908263, 0.01003723, 
    0.009727589, 0.0002689164, -0.0008461151, 0.03069137, 0.001162873, 
    0.004150509, 6.780703e-05, 1.901115e-06, 0.02790019, 0.05461546, 
    0.1021286, 0.2152727, 0.1414694, 0.03169272, 0.007364917, 0.001176541, 
    2.176355e-07, 0, 0.005892499, 0.04470744, 0.1076328, 0.05525537, 
    9.859526e-05, 4.142073e-05,
  -2.54951e-05, 0.04298412, 0.03725173, 0.0008706962, 0.007111775, 
    0.03450951, 0.026087, 0.08848736, 0.02307287, 0.0005642771, 0.0005766329, 
    0.007511775, 0.02467985, 0.01225361, 0.03257921, 0.1161535, 0.05823816, 
    7.203914e-05, -8.01919e-11, 1.090536e-08, 0, 6.488182e-08, 5.910764e-06, 
    0.1717463, 0.08490125, 0.007856808, -6.562538e-05, 4.828369e-06, 
    -7.526641e-09,
  0.006648147, 0.1669678, 0.09558362, 0.001832014, 0.0004239325, 0.06103892, 
    0.0428598, 0.04274362, 0.0562567, 0.04825178, 0.004971792, 0.01094856, 
    0.04508075, 0.05566184, 0.01287501, 0.002050867, 0.01020063, 
    1.911954e-07, 0.0005126034, 1.17046e-06, 3.973578e-07, 2.078856e-06, 
    -1.505493e-05, 0.1170479, 0.01279994, 0.000260555, 0.01371574, 
    3.000778e-05, 1.749499e-06,
  0.0218584, 0.02036753, 0.002309307, 0.001706974, 0.0005891136, 
    8.106953e-05, 0.03638677, 0.09317661, 0.1170461, 0.0356301, 0.05072482, 
    0.1127482, 0.1525863, 0.2811805, 0.09546412, 0.07762011, 0.2005313, 
    0.0728692, 0.03595055, 0.08412872, 0.09297635, 0.03274691, 0.1013036, 
    0.032859, 0.04175772, 0.1447779, 0.08847124, 0.01884743, 0.005325858,
  0.006188496, 0.00171388, 2.18406e-06, 0.001557526, 2.274896e-08, 
    0.0002040244, 0.04256551, 0.08621868, 0.06323264, 0.0466771, 0.06337675, 
    0.0403159, 0.05736193, 0.06228227, 0.003005419, 0.007325942, 0.01768804, 
    0.04222774, 0.004814198, 0.01003703, 0.02865883, 0.03721961, 0.0108648, 
    0.01369904, 0.009748084, 0.02466268, 0.05714548, 0.162981, 0.02138337,
  0.07168262, 0.04957339, -2.934715e-05, 0.005256431, 0.001869612, 
    1.265351e-07, 0.003498129, 0.06515267, 0.2725461, 0.113134, 0.07393956, 
    0.04650957, 0.05370884, 0.00244092, 0.01135226, 0.02568023, 0.0658769, 
    0.0439016, 0.03826628, 0.02107017, 0.02782275, 0.02364047, 0.05378209, 
    0.01679105, 0.07383805, 0.04956911, 0.06412559, 0.03876168, 0.07920791,
  0.1356852, 0.04079954, 0.03473365, 0.03142009, 0.02110282, 0.05592984, 
    0.02322349, 0.06157066, 0.06629883, 0.08792129, 0.1082326, 0.1543346, 
    0.2316424, 0.1672364, 0.1326724, 0.1592599, 0.1828648, 0.2192509, 
    0.0867748, 0.009698083, 0.06326969, 0.09641504, 0.1040263, 0.07729591, 
    0.1252643, 0.1308041, 0.1309122, 0.06875198, 0.04725636,
  0.111728, 0.1542412, 0.1928132, 0.1869438, 0.1424847, 0.1461614, 
    0.08595574, 0.06146124, 0.05237527, 0.08683457, 0.1456474, 0.1264914, 
    0.1676964, 0.1107164, 0.1803169, 0.2204489, 0.155979, 0.3122884, 
    0.3080142, 0.1043416, 0.120164, 0.117442, 0.1136746, 0.1777726, 
    0.1379709, 0.142333, 0.2630866, 0.1169364, 0.09915358,
  0.2278993, 0.1825146, 0.1876619, 0.2919635, 0.2437007, 0.2446845, 
    0.2292612, 0.2160325, 0.2401483, 0.1616109, 0.04302205, 0.00710119, 
    0.04640858, 0.1389936, 0.1079213, 0.1338308, 0.1244216, 0.2452555, 
    0.140843, 0.155475, 0.148353, 0.1250257, 0.113937, 0.1600259, 0.1775529, 
    0.2022477, 0.1795849, 0.1210461, 0.2205163,
  0.2461976, 0.2136698, 0.08964579, 0.1994785, 0.1781137, 0.1717423, 
    0.1714938, 0.1537462, 0.05628392, 0.03300627, 0.0738344, 0.1462625, 
    0.06088086, 0.107072, 0.1265275, 0.2280747, 0.2091525, 0.2792913, 
    0.3017732, 0.214866, 0.1184795, 0.157588, 0.1728226, 0.1621386, 
    0.1474728, 0.04829356, 0.008727804, 0.278092, 0.2450971,
  -0.003306906, 0.00127133, 0.008632963, 0.03647813, 0.03441543, 0.04324969, 
    0.04982443, 0.07388406, 0.07231295, 0.0479245, 0.01785852, 0.01189797, 
    0.03794214, 0.06813376, 0.1252907, 0.2256534, 0.1697181, 0.1341333, 
    0.07659252, 0.09116012, 0.1417599, 0.1160251, 0.0818693, 0.03454117, 
    0.01625843, -0.0005208951, -1.232506e-05, -0.01062402, 0.02105161,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0003455048, 0.00812649, 
    0.02097092, -0.001007993, 0.004475736, -1.940244e-05, 0, 0, 0.001784306, 
    0.02028886, 0.01781312, 0.01570035, 0.02955951, 0.001558341, 0,
  0.1448293, 0.05203951, 0.01156024, 0.0003832117, -0.000187073, 0, 
    0.01612039, -0.0001095355, 0, 0, 0.0001351588, -5.784473e-05, 
    0.004146298, 0.03935774, 0.0730162, 0.0787636, 0.08826166, 0.1279693, 
    0.1481422, 0.1016108, 0.1064214, 0.08409669, 0.1048034, 0.1535527, 
    0.2113935, 0.1960533, 0.2082603, 0.1872517, 0.193191,
  0.2263189, 0.1912794, 0.2833934, 0.2694972, 0.1831419, 0.1810907, 
    0.1096837, 0.09965711, 0.1370726, 0.1470028, 0.1486326, 0.2077024, 
    0.205768, 0.2218889, 0.2094631, 0.2229352, 0.2088742, 0.2224724, 
    0.2039825, 0.2131872, 0.1956921, 0.2203736, 0.1673764, 0.2304603, 
    0.1955873, 0.1603711, 0.1659843, 0.1664917, 0.1783733,
  0.1634408, 0.1331139, 0.1416092, 0.2170319, 0.1579865, 0.125291, 0.1496254, 
    0.1924071, 0.2054378, 0.2148354, 0.1907246, 0.1319619, 0.1337319, 
    0.1594526, 0.1608961, 0.1696718, 0.1296747, 0.1133689, 0.1339801, 
    0.1711898, 0.1715856, 0.1775694, 0.1816872, 0.1460902, 0.1393297, 
    0.1572606, 0.1792569, 0.2568907, 0.2241855,
  0.1505598, 0.1024131, 0.07818179, 0.08195499, 0.1024781, 0.1002633, 
    0.1233549, 0.07484784, 0.1108615, 0.06606332, 0.0277852, 0.02702694, 
    0.08145566, 0.08591174, 0.1576735, 0.1192418, 0.1828799, 0.09452102, 
    0.09785328, 0.07841836, 0.08962887, 0.05929033, 0.04497848, 0.05882721, 
    0.08971725, 0.09896858, 0.1551279, 0.1157354, 0.1267755,
  0.01820184, 0.004286622, 0.05106082, 0.1052967, 0.05501069, 0.02596671, 
    0.007143129, 0.001983738, 0.00228674, 5.954873e-05, 0.02462263, 
    0.05720134, 0.1077562, 0.06469985, 0.1262434, 0.02963493, 0.03067818, 
    0.03190864, 0.2649254, 0.1811815, 0.06802449, 0.01355274, 0.001705411, 
    0.001125447, 0.04120879, 0.06223276, 0.1117552, 0.0987627, 0.0766003,
  3.392667e-06, 0.009323303, 0.037496, 0.001221059, 0.01183502, 0.002145073, 
    0.0002272753, -0.000677076, 0.01114379, 0.002084696, 0.004795955, 
    1.235699e-05, 0.002743743, 0.04558584, 0.05637807, 0.1084059, 0.2015647, 
    0.1223424, 0.02353617, 0.01761103, 9.751636e-05, -9.251258e-07, 0, 
    0.0022521, 0.04522373, 0.1022873, 0.05558451, 2.286954e-05, 2.015172e-05,
  0.006183011, 0.05596527, 0.03273872, 0.0008487933, 0.00764354, 0.03839429, 
    0.0269239, 0.08101838, 0.01182188, 0.0008133902, 0.0007544757, 
    0.003570488, 0.04391638, 0.008871951, 0.02725673, 0.1330225, 0.05246793, 
    0.000112007, 8.880993e-09, 2.34571e-10, 0, 1.118889e-09, 1.546677e-05, 
    0.1656133, 0.06748796, 0.007620402, -3.163928e-05, 1.098269e-06, 
    -8.155855e-05,
  0.02202134, 0.1883351, 0.07668247, 0.002324498, 0.00703225, 0.0800468, 
    0.05383992, 0.04153749, 0.04268778, 0.03393067, 0.002996362, 0.01091837, 
    0.03758319, 0.04141379, 0.01051084, 0.002271723, 0.006783925, 
    1.409022e-07, 0.0001587896, 1.823346e-05, 1.208025e-07, 1.106927e-06, 
    0.00178688, 0.08859572, 0.01121614, 0.001205367, 0.005240251, 
    0.0006414658, 1.379187e-06,
  0.01980178, 0.01986683, 0.005359351, 0.002227985, 0.0005324309, 
    0.0001911208, 0.03882691, 0.08603562, 0.1220479, 0.03234169, 0.04315707, 
    0.1116043, 0.1393114, 0.2786219, 0.08359208, 0.07979123, 0.1807586, 
    0.07724733, 0.03820297, 0.07776416, 0.1011303, 0.03047406, 0.09964865, 
    0.02620473, 0.04172672, 0.1274759, 0.07329016, 0.01321556, 0.01414992,
  0.00377332, 1.450328e-05, 1.664043e-06, 0.00110898, 4.064139e-08, 
    0.0001523958, 0.04509854, 0.09321573, 0.06368638, 0.03730304, 0.06263278, 
    0.04443699, 0.05929301, 0.06037566, 0.002572293, 0.00610735, 0.01212508, 
    0.04139955, 0.00284221, 0.0118517, 0.01087714, 0.04440278, 0.008995244, 
    0.01436625, 0.007028027, 0.01363189, 0.03235562, 0.1358571, 0.0009581922,
  0.05379409, 0.04013309, -4.02187e-06, 0.003975905, 0.001830594, 
    -1.88644e-07, 0.003012406, 0.0831484, 0.2951705, 0.1126211, 0.06383707, 
    0.045282, 0.05673979, 0.002376933, 0.01729397, 0.02246425, 0.04473361, 
    0.03745587, 0.0312382, 0.01713335, 0.02816238, 0.02238461, 0.05245204, 
    0.01118502, 0.06099455, 0.03913554, 0.0505622, 0.02337135, 0.08506572,
  0.1097344, 0.03547716, 0.03987565, 0.03497021, 0.01596486, 0.05394802, 
    0.02136988, 0.05246399, 0.06096049, 0.09640786, 0.09420168, 0.1559008, 
    0.2142723, 0.1886241, 0.1321033, 0.1430852, 0.1791125, 0.1745807, 
    0.05883157, 0.009987986, 0.07043856, 0.1057504, 0.1129517, 0.07580877, 
    0.1064147, 0.1070176, 0.1152429, 0.09392773, 0.04048919,
  0.09870572, 0.1626552, 0.2011595, 0.2215994, 0.1470578, 0.1514741, 
    0.06885141, 0.09912439, 0.1205628, 0.147897, 0.1681601, 0.1592898, 
    0.1782669, 0.1086293, 0.1814848, 0.2032517, 0.1565708, 0.295985, 
    0.2925661, 0.09504766, 0.1317403, 0.1355784, 0.1489662, 0.1789387, 
    0.1429691, 0.1606949, 0.2308768, 0.1029366, 0.07435994,
  0.2468713, 0.2204097, 0.2224407, 0.3820914, 0.2620544, 0.2423972, 0.206831, 
    0.2035925, 0.2846148, 0.24693, 0.09083489, 0.07246472, 0.1715393, 
    0.1908062, 0.2041538, 0.2422768, 0.1544973, 0.2798663, 0.1670064, 
    0.1599444, 0.1523433, 0.1833783, 0.1971297, 0.1966028, 0.2338676, 
    0.2371774, 0.1946602, 0.139202, 0.2324446,
  0.3290045, 0.2630506, 0.2100424, 0.2741103, 0.3098651, 0.2206287, 
    0.2784896, 0.3022039, 0.1673643, 0.1937727, 0.1538624, 0.262409, 
    0.1499967, 0.1706828, 0.2166949, 0.2151089, 0.2304239, 0.3153532, 
    0.3452103, 0.3122654, 0.2034989, 0.1643725, 0.2024277, 0.2249483, 
    0.1462519, 0.09917566, 0.06264479, 0.3081155, 0.2942728,
  0.06831346, 0.02731924, 0.05402591, 0.128682, 0.1604912, 0.1101915, 
    0.1102028, 0.1534257, 0.1085277, 0.06794417, 0.08844761, 0.090882, 
    0.1125014, 0.1784323, 0.2416368, 0.3094158, 0.2133859, 0.1560882, 
    0.1061388, 0.1166962, 0.1681054, 0.1960111, 0.1488465, 0.1438439, 
    0.09192277, 0.005454755, -0.01250944, 0.1036967, 0.1115649,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.004604199, 0.03187829, 0.04065477, 
    0.06654239, 0.0507432, 0.02334858, 0.0001095047, -3.81354e-06, 0, 
    0.005244297, 0.3127878, 0.2832868, 0.113144, 0.1163361, 0.006417034, 
    1.842604e-06,
  0.1800574, 0.09663274, 0.02841494, 0.006349053, -0.0007186293, 
    -0.0004070476, 0.04782957, 0.002805777, -0.0001654798, -9.379951e-05, 
    0.0001024574, -0.0001663686, 0.01091065, 0.1537879, 0.1525786, 0.136731, 
    0.1799167, 0.1860989, 0.2073565, 0.1771332, 0.1760236, 0.1882208, 
    0.3085009, 0.3085421, 0.2942903, 0.2574613, 0.2377086, 0.2428629, 
    0.3088749,
  0.2336832, 0.2184183, 0.3138481, 0.297225, 0.2081025, 0.1860515, 0.1326188, 
    0.1184759, 0.1697802, 0.2093333, 0.1853485, 0.2679716, 0.2451651, 
    0.2946527, 0.257569, 0.235873, 0.2193493, 0.2461664, 0.2288929, 
    0.2524177, 0.2458593, 0.2387846, 0.2067777, 0.2644667, 0.2262894, 
    0.163894, 0.1810549, 0.1687179, 0.1660278,
  0.1657603, 0.1193652, 0.1306208, 0.2077188, 0.1468788, 0.11118, 0.1451661, 
    0.1889819, 0.2045381, 0.1960447, 0.1903806, 0.141363, 0.1451563, 
    0.159003, 0.163336, 0.1749531, 0.1158038, 0.1148201, 0.1320951, 0.165697, 
    0.1691153, 0.1813362, 0.1746889, 0.1298891, 0.133116, 0.1561451, 
    0.1557627, 0.2355135, 0.2148364,
  0.1379981, 0.09537945, 0.073645, 0.0610417, 0.09309593, 0.110158, 
    0.1050082, 0.09171196, 0.1026362, 0.05182667, 0.02331236, 0.03160127, 
    0.07929986, 0.09007116, 0.1627137, 0.1118397, 0.1772744, 0.08535021, 
    0.09269362, 0.06573483, 0.0838448, 0.05962716, 0.04081695, 0.04568601, 
    0.08634124, 0.08904153, 0.1397641, 0.106255, 0.1078171,
  0.01737166, 0.009479938, 0.04407587, 0.110897, 0.03343528, 0.0204039, 
    0.01512103, 0.00679413, 0.001072577, 0.004309429, 0.02418234, 0.06512666, 
    0.114286, 0.06552823, 0.1003601, 0.02445624, 0.03214717, 0.01914576, 
    0.2663899, 0.1905933, 0.05492986, 0.00729274, 0.0003399738, -7.4007e-05, 
    0.04494397, 0.05837075, 0.1044968, 0.0795573, 0.06525084,
  1.14934e-06, 0.01117462, 0.02591695, 0.0009495708, 0.01670282, 
    4.046862e-06, 0.0002621863, -0.0002193432, 0.002352988, 0.0002200651, 
    0.01394381, 0.001134867, 0.01098362, 0.06890584, 0.05827217, 0.105841, 
    0.1742753, 0.1136565, 0.01660188, 0.02927775, 4.736908e-06, 7.531406e-05, 
    -2.016852e-10, 0.0002534018, 0.04481016, 0.1012556, 0.06665833, 
    5.924752e-05, 3.735179e-06,
  8.619732e-05, 0.05697215, 0.02246637, 0.001345465, 0.02061571, 0.03597543, 
    0.03278128, 0.07444853, 0.01246732, 0.0005803299, 0.001038835, 
    0.003589903, 0.05536261, 0.006898013, 0.04268048, 0.1364531, 0.02997388, 
    0.0003330245, 9.449004e-08, -5.852466e-10, -6.277013e-11, 7.57015e-09, 
    1.813783e-05, 0.1553869, 0.05694294, 0.01715188, 1.157111e-05, 
    4.659978e-07, 0.009140271,
  0.03159138, 0.2153357, 0.07472859, 0.002855877, 0.0161081, 0.08331212, 
    0.05951058, 0.03981234, 0.03046163, 0.03073197, 0.002259159, 0.009284952, 
    0.01457574, 0.03424035, 0.009771033, 0.002988667, 0.000995845, 
    1.833908e-06, 4.118442e-05, 2.047317e-05, 1.892138e-07, 1.404499e-07, 
    0.009659551, 0.07561269, 0.01052478, 0.002102544, 0.001798538, 
    0.001512319, 0.003862758,
  0.01907305, 0.01069993, 0.006416152, 0.003740925, 0.00113436, 0.000381021, 
    0.03518549, 0.08257531, 0.1295309, 0.04067186, 0.04610845, 0.1086733, 
    0.1386872, 0.2780935, 0.07619443, 0.09153625, 0.1726251, 0.08464766, 
    0.04664615, 0.07360215, 0.1097301, 0.03795498, 0.1012742, 0.02276029, 
    0.04426867, 0.1160588, 0.05695901, 0.009362795, 0.0181547,
  0.001347118, 1.261524e-06, 1.014214e-06, 0.00121141, 3.636936e-08, 
    2.65732e-05, 0.05366915, 0.098683, 0.05055281, 0.03572131, 0.05811798, 
    0.04821209, 0.06270507, 0.05921932, 0.004315382, 0.005360935, 
    0.006785692, 0.02165284, 0.0007283918, 0.01386437, 0.008629568, 
    0.05478827, 0.009527382, 0.01878069, 0.006789233, 0.01092988, 0.01546114, 
    0.0885663, -1.985475e-06,
  0.05032486, 0.04113065, 0.0001220763, 0.00278727, 0.0007315259, 
    -5.571417e-08, 0.002143494, 0.116785, 0.3181266, 0.1370236, 0.05464175, 
    0.04328994, 0.06524304, 0.00370282, 0.02163555, 0.02699658, 0.03679545, 
    0.02865046, 0.020199, 0.00280963, 0.01847433, 0.02247952, 0.04954545, 
    0.01205823, 0.05593919, 0.03284566, 0.04632547, 0.01828358, 0.07314039,
  0.1008104, 0.03646767, 0.04995272, 0.03958099, 0.01870399, 0.05106325, 
    0.03125351, 0.0434424, 0.06217351, 0.09387955, 0.07164368, 0.133672, 
    0.2090844, 0.1996405, 0.128806, 0.1414773, 0.1763017, 0.1685893, 
    0.04413872, 0.009700932, 0.08620542, 0.113562, 0.1148526, 0.07885969, 
    0.09467465, 0.0950437, 0.1095738, 0.1110552, 0.03534743,
  0.09311623, 0.1759863, 0.1813603, 0.2224506, 0.1281333, 0.1354361, 
    0.05436596, 0.1443216, 0.1977905, 0.1477639, 0.1676755, 0.1980327, 
    0.1864084, 0.1140816, 0.1789172, 0.2137479, 0.1512581, 0.2947818, 
    0.2902493, 0.1203152, 0.1390809, 0.1564558, 0.1979437, 0.1930696, 
    0.1662348, 0.1670673, 0.2069371, 0.1009604, 0.08383296,
  0.2507225, 0.2469394, 0.2208036, 0.4077923, 0.3102886, 0.2334741, 
    0.1956995, 0.1876206, 0.2686437, 0.2559451, 0.1556499, 0.09377716, 
    0.2130299, 0.1800511, 0.2350612, 0.2463127, 0.173403, 0.3034991, 
    0.2460754, 0.1524071, 0.1727304, 0.1755833, 0.2227779, 0.223538, 
    0.2501062, 0.2467815, 0.1917034, 0.1293882, 0.2028077,
  0.3110588, 0.2734685, 0.2408053, 0.3429712, 0.3707492, 0.2632858, 
    0.3475904, 0.3902655, 0.2422012, 0.3000326, 0.2259096, 0.3899333, 
    0.1759389, 0.2251704, 0.2093386, 0.1981941, 0.2393663, 0.2966891, 
    0.3541795, 0.3359393, 0.2432714, 0.1889654, 0.224396, 0.2226368, 
    0.1657043, 0.1576521, 0.119354, 0.3261629, 0.3624221,
  0.1252659, 0.05486387, 0.1485679, 0.2274606, 0.2439612, 0.2244265, 
    0.2262244, 0.2225891, 0.1903815, 0.1261318, 0.09131318, 0.1575808, 
    0.1918933, 0.2402254, 0.2823555, 0.3177553, 0.1966314, 0.1364228, 
    0.1161802, 0.1399227, 0.1780882, 0.2070356, 0.153771, 0.1594185, 
    0.1522482, 0.03653026, 0.07551612, 0.1126181, 0.1778107,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  -1.821549e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0004390597, 0.06385583, 
    0.06884462, 0.08480014, 0.1546361, 0.1036378, 0.06637368, 0.002761332, 
    0.004234453, 0.002590545, 0.05886758, 0.4016886, 0.340447, 0.2447879, 
    0.2029829, 0.06668459, 0.0001879972,
  0.1794046, 0.1323269, 0.07187157, 0.05814554, 0.00207357, -0.003322045, 
    0.09777228, 0.002593562, -0.0001660156, -0.001839741, 0.001588834, 
    -0.000274484, 0.07636501, 0.2098149, 0.2101211, 0.1934935, 0.2419054, 
    0.2474372, 0.2322191, 0.2705544, 0.2964472, 0.2865539, 0.4287514, 
    0.4318733, 0.298364, 0.2537569, 0.2100734, 0.2583496, 0.3449163,
  0.2389796, 0.2269285, 0.3066268, 0.3110368, 0.2362092, 0.1978764, 
    0.1430477, 0.1435241, 0.2301701, 0.2680491, 0.2407652, 0.2826089, 
    0.2679937, 0.30439, 0.2751188, 0.2263803, 0.2179806, 0.2410215, 
    0.2307246, 0.2539383, 0.2600467, 0.2654922, 0.2292336, 0.2749748, 
    0.230773, 0.1661816, 0.1771001, 0.1653432, 0.1666686,
  0.1709399, 0.1193511, 0.1297816, 0.2009958, 0.1425934, 0.1053138, 
    0.1436288, 0.1947466, 0.2160783, 0.218364, 0.172235, 0.1479426, 
    0.1372142, 0.1614355, 0.1589219, 0.1451403, 0.1125053, 0.1065583, 
    0.1152023, 0.1473956, 0.167436, 0.183081, 0.158541, 0.1160052, 0.1261949, 
    0.1614257, 0.1493453, 0.2178345, 0.2009865,
  0.1293537, 0.09288998, 0.06573919, 0.07024918, 0.09473414, 0.1032302, 
    0.1299089, 0.08259715, 0.1075525, 0.03682569, 0.02334698, 0.03585982, 
    0.07825355, 0.07739355, 0.1663369, 0.09782504, 0.1545232, 0.08784062, 
    0.08231315, 0.05639961, 0.0671384, 0.04867293, 0.03968112, 0.03715996, 
    0.07681198, 0.07050233, 0.1230332, 0.1006177, 0.09584004,
  0.0197835, 0.009998908, 0.03889405, 0.1095909, 0.02811675, 0.01471935, 
    0.01579715, 0.0003386175, 0.003219167, 0.01538482, 0.03813553, 
    0.07609285, 0.1111689, 0.06686781, 0.08962809, 0.02115547, 0.02567981, 
    0.01878456, 0.2448215, 0.1706716, 0.04550887, 0.01059975, 0.0005565524, 
    -1.840322e-05, 0.05198238, 0.04835076, 0.1098127, 0.06827503, 0.06261102,
  6.921649e-08, 0.009250964, 0.02136189, 0.002462663, 0.02492437, 
    5.078403e-05, 0.0005702461, -0.0004729579, 0.001076376, 2.443253e-05, 
    0.03514932, 0.002980596, 0.01525554, 0.0800138, 0.06992008, 0.09972672, 
    0.1480884, 0.09852616, 0.01788009, 0.03344019, 4.051202e-06, 0.007292205, 
    -1.86292e-09, 0.0001335562, 0.05060579, 0.1036968, 0.08195655, 
    -3.751669e-05, 1.819372e-06,
  -1.215045e-05, 0.06621324, 0.02593173, 0.007280948, 0.01919693, 0.03469743, 
    0.03602945, 0.06454537, 0.02105682, 0.0005887668, 0.0022504, 0.00752122, 
    0.06123945, 0.006749808, 0.07587051, 0.1346512, 0.02966727, 7.796301e-05, 
    5.74063e-08, 8.762712e-09, 3.47996e-09, 1.265182e-07, 0.0009588395, 
    0.1545977, 0.06205652, 0.01585409, 2.0509e-05, 2.526801e-07, 0.0005352387,
  0.08750218, 0.2674434, 0.09561626, 0.01086465, 0.01340369, 0.07570411, 
    0.05554925, 0.03813661, 0.03832156, 0.03565412, 0.002533856, 0.009392455, 
    0.006658077, 0.03724335, 0.01087771, 0.003643775, 0.005958226, 
    7.700859e-06, 0.001932661, 2.677804e-07, 1.18404e-07, -8.211789e-06, 
    0.04181338, 0.07379616, 0.009378383, 0.001730697, 0.001915419, 
    0.001570511, 0.01817356,
  0.01953345, 0.01168169, 0.009636922, 0.001985506, 0.001943602, 0.001340511, 
    0.04102148, 0.0705779, 0.1591363, 0.04288325, 0.05710444, 0.1064559, 
    0.1486731, 0.286153, 0.08471934, 0.09698901, 0.1977621, 0.09335595, 
    0.05913297, 0.0668753, 0.1070626, 0.04641014, 0.1090159, 0.0270639, 
    0.05116108, 0.1313471, 0.03840115, 0.01331755, 0.01493838,
  0.006818504, 6.999102e-07, 6.165963e-07, 0.00632122, 1.58263e-08, 
    1.692521e-05, 0.05197922, 0.1086988, 0.0378425, 0.03663322, 0.05774225, 
    0.0733039, 0.0693187, 0.05926517, 0.006193236, 0.006039701, 0.006490634, 
    0.01231441, 0.0001954826, 0.02099042, 0.005931239, 0.06824746, 
    0.01055915, 0.02879107, 0.008714698, 0.009278812, 0.001938392, 
    0.04671157, 0.0002122037,
  0.04953093, 0.03517174, 0.00351, 0.0006268838, 0.002425649, 2.575831e-08, 
    0.002126416, 0.1568396, 0.3318247, 0.1362821, 0.04747077, 0.03857278, 
    0.07202177, 0.01182348, 0.0243599, 0.03349433, 0.02020073, 0.02405571, 
    0.02160818, 0.0005542334, 0.0119951, 0.0271935, 0.04898974, 0.01176759, 
    0.04973055, 0.03152367, 0.04758568, 0.02037948, 0.072396,
  0.08544168, 0.0395369, 0.07254703, 0.04114545, 0.03178423, 0.04802246, 
    0.03384889, 0.03428984, 0.05985149, 0.09089872, 0.0705278, 0.1458284, 
    0.2175984, 0.1676975, 0.1320933, 0.149969, 0.1552354, 0.1461526, 
    0.04258991, 0.0109877, 0.08338914, 0.1083598, 0.1089225, 0.07861928, 
    0.08030181, 0.08784067, 0.1050768, 0.09235892, 0.05403665,
  0.1042256, 0.1841035, 0.2193633, 0.2268897, 0.1384161, 0.1241703, 
    0.05050535, 0.1513012, 0.2108471, 0.1378309, 0.1470275, 0.1940825, 
    0.1732244, 0.1231224, 0.1828085, 0.1974702, 0.1558404, 0.2886724, 
    0.2650308, 0.1290677, 0.1452366, 0.1717279, 0.2195321, 0.2225393, 
    0.1764497, 0.1551033, 0.1816199, 0.1056391, 0.1049865,
  0.247493, 0.2558887, 0.2188956, 0.4069083, 0.3111044, 0.2274601, 0.1818153, 
    0.175049, 0.2630154, 0.259074, 0.1655419, 0.1166222, 0.2550634, 
    0.1707719, 0.228888, 0.2353762, 0.1723561, 0.3159859, 0.2691384, 
    0.1294651, 0.1874162, 0.1816391, 0.2289076, 0.2617349, 0.2517026, 
    0.2548332, 0.1912732, 0.1451434, 0.2300017,
  0.2729241, 0.2934507, 0.248649, 0.3487813, 0.3689471, 0.2641831, 0.3486388, 
    0.3924275, 0.2832626, 0.3299187, 0.2650629, 0.3991298, 0.1882977, 
    0.2349963, 0.2331705, 0.1831569, 0.2380423, 0.2884487, 0.3530079, 
    0.3371953, 0.258731, 0.1756151, 0.1766546, 0.2587689, 0.1615872, 
    0.2248743, 0.1767701, 0.3234055, 0.3341733,
  0.1312369, 0.1194815, 0.1811714, 0.2841806, 0.3187928, 0.2345596, 
    0.2413047, 0.235488, 0.1875663, 0.1392543, 0.1016998, 0.1386637, 
    0.1772238, 0.227898, 0.2742428, 0.2723651, 0.1776599, 0.118406, 
    0.1080948, 0.1386198, 0.1764485, 0.2094298, 0.1689308, 0.2292703, 
    0.1897781, 0.1070362, 0.1199169, 0.1400227, 0.1873434,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001579054, 0.1603593, 0.07443764, 
    0.1129198, 0.162479, 0.1736176, 0.1007719, 0.02997612, 0.01055894, 
    0.008029808, 0.1470956, 0.3678686, 0.3511655, 0.2763898, 0.2167218, 
    0.1695677, 0.005663943,
  0.1754038, 0.1454644, 0.07045449, 0.1239421, 0.009351905, 0.01806614, 
    0.1610946, 0.005917348, -0.001201919, -0.004232503, 0.002912571, 
    0.009261867, 0.1650772, 0.2947083, 0.273362, 0.2214441, 0.297596, 
    0.2629302, 0.2872769, 0.3217592, 0.3406035, 0.3201837, 0.4411099, 
    0.4716852, 0.304056, 0.2197847, 0.2191613, 0.2707835, 0.3286605,
  0.242628, 0.2387335, 0.3026511, 0.3092777, 0.2477473, 0.2119861, 0.1809463, 
    0.1645816, 0.257787, 0.2728463, 0.2357857, 0.2758204, 0.2846265, 
    0.2957913, 0.2804591, 0.2434708, 0.2302169, 0.2641222, 0.2382278, 
    0.2817744, 0.2552153, 0.2698483, 0.2156629, 0.2654373, 0.2234062, 
    0.1625962, 0.1593767, 0.1563998, 0.1594245,
  0.1859264, 0.1495076, 0.1238386, 0.198794, 0.1708663, 0.1059859, 0.167434, 
    0.1984585, 0.2133554, 0.2133409, 0.1712856, 0.1668701, 0.1260198, 
    0.1577918, 0.1656653, 0.1418517, 0.117623, 0.1112529, 0.1156677, 
    0.1449963, 0.1778081, 0.1884641, 0.1610068, 0.1043164, 0.1157329, 
    0.1836788, 0.1519899, 0.1962011, 0.1924131,
  0.1361537, 0.09967059, 0.05719016, 0.07766917, 0.1018668, 0.1126909, 
    0.1287078, 0.09397903, 0.107019, 0.02657063, 0.02257424, 0.02765834, 
    0.07803123, 0.09489442, 0.1705584, 0.08591482, 0.1360105, 0.09165448, 
    0.08408321, 0.05933096, 0.05983785, 0.0547761, 0.05217266, 0.04297611, 
    0.06797472, 0.07674392, 0.1181743, 0.1031165, 0.1052433,
  0.00441794, 0.008623905, 0.03729486, 0.1118223, 0.03763533, 0.01221779, 
    0.01997686, -0.0001723862, 0.004386491, 0.01505807, 0.03046827, 
    0.09358575, 0.1099738, 0.06441651, 0.07783478, 0.0167771, 0.01693773, 
    0.01505954, 0.2337225, 0.1661752, 0.04266373, 0.011211, 0.0001323294, 
    -5.903649e-06, 0.05538977, 0.04218617, 0.1141998, 0.06449258, 0.06979078,
  -1.320361e-08, 0.01874987, 0.03121615, 0.004351093, 0.01975933, 
    -2.231997e-05, 0.0005390336, -0.0002423144, 0.002172725, 9.850268e-06, 
    0.1078444, 0.054492, 0.0141132, 0.09115504, 0.07169629, 0.08512525, 
    0.129278, 0.08010602, 0.02178507, 0.03728395, 1.301237e-05, 0.01346268, 
    6.442248e-09, 0.0001223547, 0.06288087, 0.09162512, 0.09537411, 
    -2.998758e-05, 1.223045e-06,
  0.001969914, 0.07248744, 0.03522778, 0.01645478, 0.01296481, 0.04723538, 
    0.05720552, 0.06403586, 0.02483195, 0.0006783559, 0.002855205, 
    0.01709619, 0.07856634, 0.01193169, 0.1061062, 0.1413538, 0.02986305, 
    0.001279362, 5.705631e-07, 3.203934e-08, 8.172933e-08, 2.501931e-06, 
    0.004196574, 0.1714553, 0.07853663, 0.02917214, 3.046933e-05, 
    5.698521e-08, 3.943048e-06,
  0.1322238, 0.3116516, 0.1588861, 0.01111779, 0.01079623, 0.08524907, 
    0.04514408, 0.03862654, 0.04909826, 0.05011324, 0.003947855, 0.01046318, 
    0.009968303, 0.04837334, 0.01424211, 0.00312614, 0.00309191, 
    4.021326e-05, 0.006227714, 1.297079e-07, 3.459463e-07, -0.0001120949, 
    0.06363929, 0.08738565, 0.006835971, 0.001056635, 0.004213961, 
    0.006592514, 0.07119416,
  0.02435192, 0.01360433, 0.01106492, 0.00490399, 0.00178295, 0.001035712, 
    0.05123395, 0.06868675, 0.1974431, 0.0468859, 0.07929514, 0.1293103, 
    0.1702374, 0.3072356, 0.09689146, 0.1154302, 0.2206164, 0.1171824, 
    0.08956054, 0.06904233, 0.1056971, 0.07054723, 0.1249281, 0.04106911, 
    0.06575004, 0.1418242, 0.03195203, 0.02414189, 0.01531933,
  0.02423321, 8.524757e-05, 5.09644e-07, 0.01137376, 3.73074e-08, 
    0.001502502, 0.05030036, 0.1344341, 0.02919568, 0.03540686, 0.0710222, 
    0.09298977, 0.08066346, 0.07047778, 0.01212701, 0.01395077, 0.008369223, 
    0.007104435, 0.0004966282, 0.02416103, 0.02368912, 0.09795637, 
    0.01652084, 0.03862853, 0.01433749, 0.009830577, 0.005277368, 0.02873729, 
    -6.237296e-05,
  0.03872288, 0.02371924, 0.005207126, -0.0001123256, 0.007280327, 
    5.674071e-08, 0.006132799, 0.1631313, 0.3492742, 0.1138573, 0.04351588, 
    0.0369545, 0.07974873, 0.014163, 0.03019687, 0.03649146, 0.02002599, 
    0.02303129, 0.02220767, 0.002464557, 0.01123052, 0.04841467, 0.05215511, 
    0.01854542, 0.05086933, 0.03528421, 0.05388797, 0.02129822, 0.0701607,
  0.06640527, 0.04469006, 0.0847467, 0.05416673, 0.05850961, 0.04216462, 
    0.03404515, 0.02562416, 0.05183828, 0.08109183, 0.07491124, 0.1496674, 
    0.1953371, 0.1631509, 0.1457497, 0.1533858, 0.1472451, 0.140354, 
    0.03970328, 0.01386076, 0.07387505, 0.1159374, 0.09701176, 0.07918444, 
    0.08219172, 0.0871957, 0.09789582, 0.08861732, 0.02113186,
  0.09247178, 0.2242112, 0.2036499, 0.2139893, 0.1244168, 0.118211, 
    0.0505088, 0.151507, 0.1955572, 0.1257783, 0.1269165, 0.1953392, 
    0.1511255, 0.1267618, 0.1736091, 0.2094752, 0.1485357, 0.2655181, 
    0.228154, 0.1259929, 0.1317866, 0.1693044, 0.2288577, 0.2212763, 
    0.1959994, 0.1512562, 0.1626467, 0.09646357, 0.07683145,
  0.2341879, 0.2631995, 0.2455724, 0.4105937, 0.3215928, 0.2043412, 
    0.1639682, 0.1657476, 0.2379504, 0.2435904, 0.1892234, 0.1182547, 
    0.2602037, 0.1650834, 0.2241023, 0.2260991, 0.1769429, 0.3286726, 
    0.2652303, 0.1092106, 0.2017627, 0.1860932, 0.2382458, 0.2462991, 
    0.3059697, 0.2765659, 0.2180775, 0.1250779, 0.220219,
  0.245971, 0.2900164, 0.2600707, 0.3843844, 0.3669197, 0.2556331, 0.3425104, 
    0.3905838, 0.3016418, 0.3088814, 0.2473412, 0.4075328, 0.1997513, 
    0.2325657, 0.2476307, 0.1945468, 0.2466064, 0.2662475, 0.3487596, 
    0.3398302, 0.2306877, 0.1804236, 0.1248413, 0.2814293, 0.1683427, 
    0.2885604, 0.2434095, 0.3144406, 0.289099,
  0.1163854, 0.148565, 0.1788593, 0.2969938, 0.350937, 0.2252181, 0.2271324, 
    0.2301643, 0.194779, 0.1269415, 0.08936308, 0.1239062, 0.1622137, 
    0.2229295, 0.2641168, 0.2237463, 0.1795778, 0.1190773, 0.104347, 
    0.1380836, 0.1765512, 0.2195456, 0.1585626, 0.2187057, 0.1826577, 
    0.1443479, 0.1536056, 0.1407881, 0.1843804,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  -0.005257796, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.009493772, 0.2007388, 
    0.06226846, 0.09296577, 0.143131, 0.1667809, 0.151532, 0.08995047, 
    0.111309, 0.08349633, 0.2705911, 0.3504965, 0.3276866, 0.2584308, 
    0.1854537, 0.1956538, 0.0492519,
  0.1774332, 0.1507495, 0.06595391, 0.1268112, 0.0185909, 0.0602614, 
    0.1662929, 0.01861854, 0.001745855, 0.01604176, 0.005536756, 0.01389639, 
    0.2238381, 0.2979843, 0.2722447, 0.2203173, 0.2922853, 0.2624553, 
    0.2873138, 0.306019, 0.356575, 0.336682, 0.4364461, 0.5036197, 0.2773753, 
    0.190222, 0.2277209, 0.2597496, 0.2994454,
  0.245445, 0.2489613, 0.3260036, 0.3172048, 0.2424253, 0.222924, 0.1726896, 
    0.1695327, 0.2720754, 0.2752142, 0.2411565, 0.2801066, 0.2782854, 
    0.2789376, 0.284753, 0.2466741, 0.2254384, 0.254135, 0.2433832, 
    0.2825908, 0.2502116, 0.2297331, 0.2128024, 0.2593066, 0.2158978, 
    0.1570113, 0.1351058, 0.1532076, 0.1544414,
  0.2030092, 0.1237319, 0.1434829, 0.2266375, 0.1717698, 0.1077069, 
    0.1626934, 0.1906448, 0.1964948, 0.2276312, 0.1856595, 0.1712738, 
    0.1328538, 0.1635909, 0.1511557, 0.1259123, 0.1101639, 0.117341, 
    0.1167375, 0.1263475, 0.1818718, 0.1806304, 0.1630605, 0.1081483, 
    0.1108247, 0.1899411, 0.1537657, 0.1786251, 0.1868981,
  0.1347901, 0.09895302, 0.05979721, 0.08181488, 0.08837236, 0.1240788, 
    0.1268118, 0.09698393, 0.1113779, 0.02910784, 0.01404687, 0.00911923, 
    0.08106983, 0.10811, 0.1715702, 0.07223292, 0.1266573, 0.0951058, 
    0.09257119, 0.06006625, 0.06710324, 0.05268349, 0.04876752, 0.05375537, 
    0.06414184, 0.08063763, 0.1176601, 0.09857824, 0.1157574,
  0.005942449, 0.001836539, 0.04952934, 0.1303903, 0.06083931, 0.01393539, 
    0.0186668, -0.0003423259, 0.006521369, 0.00951122, 0.0237683, 0.0746376, 
    0.1169581, 0.07561602, 0.06087566, 0.01993078, 0.01866413, 0.01049119, 
    0.2243124, 0.1729541, 0.05371932, 0.005110864, -1.333754e-05, 
    -1.253111e-06, 0.05341623, 0.03861074, 0.1270336, 0.06793655, 0.07262352,
  -1.88405e-05, 0.02111572, 0.06619851, 0.001963376, 0.01863831, 
    -7.661427e-08, 0.001297975, 0.001395689, 0.001861951, 2.756465e-06, 
    0.1527629, 0.04806136, 0.01223272, 0.08847578, 0.07343302, 0.08163139, 
    0.1252975, 0.09501408, 0.02658449, 0.03899495, -0.0001293203, 
    0.0004312084, 2.228244e-09, 6.474633e-06, 0.08058493, 0.1120635, 
    0.09761331, -3.954057e-06, 2.939051e-06,
  0.007203216, 0.1062181, 0.1002492, 0.01398004, 0.01732237, 0.07120931, 
    0.06615331, 0.08017685, 0.02665107, 0.0006781967, 0.00310736, 0.0288529, 
    0.07850327, 0.01914023, 0.1447169, 0.1389341, 0.0361045, 0.006706725, 
    2.754498e-06, 3.815194e-08, 4.594713e-07, 0.0002882766, 0.001219303, 
    0.2029961, 0.1191929, 0.1450314, 2.357761e-05, 1.285708e-08, 3.579116e-07,
  0.1425169, 0.3715082, 0.2156296, 0.007620022, 0.001797659, 0.08308702, 
    0.04887509, 0.04444625, 0.08258918, 0.07002462, 0.006851761, 0.01144892, 
    0.01623455, 0.07358656, 0.02007485, 0.005966499, 0.0001000755, 
    0.002405622, 0.002760575, 9.933883e-08, 9.086591e-06, 0.004309153, 
    0.09949472, 0.1087234, 0.007059064, 0.0008207082, 0.005545771, 
    0.01086001, 0.04226305,
  0.02609747, 0.01569116, 0.009788913, 0.02464126, 0.002195106, 0.001389757, 
    0.05745927, 0.06994285, 0.2154591, 0.04514536, 0.09729781, 0.1419941, 
    0.1881007, 0.3210429, 0.09817391, 0.139472, 0.2256351, 0.1374156, 
    0.1126618, 0.0785714, 0.1172395, 0.09161026, 0.143831, 0.04599173, 
    0.08104099, 0.1624096, 0.03776831, 0.03412519, 0.01758294,
  0.01283424, 2.499225e-05, 8.06795e-07, 0.006609664, 9.09257e-08, 
    0.0008529351, 0.05949362, 0.1264123, 0.03606476, 0.04295497, 0.07519248, 
    0.1144328, 0.07686545, 0.08246154, 0.0143171, 0.02699534, 0.01251277, 
    0.006651337, 0.002629363, 0.04204277, 0.03792379, 0.1300635, 0.01938904, 
    0.03959962, 0.01606776, 0.01607993, 0.007803642, 0.03075584, 4.657317e-05,
  0.01131639, 0.01584068, 0.007870878, -0.0001042481, 0.01004351, 
    3.115739e-07, 0.004749826, 0.1593799, 0.3560004, 0.07626151, 0.04740559, 
    0.04004357, 0.08492672, 0.01788846, 0.03974779, 0.03245026, 0.02155374, 
    0.02543767, 0.02146317, 0.004337863, 0.02303225, 0.06050159, 0.06034126, 
    0.02363791, 0.06281363, 0.04300549, 0.06653832, 0.01340554, 0.06690335,
  0.05442927, 0.04581209, 0.09905472, 0.07022604, 0.07925861, 0.03076996, 
    0.03147266, 0.01810344, 0.04625449, 0.07000729, 0.08708216, 0.1427147, 
    0.1716307, 0.1645135, 0.1499041, 0.1605327, 0.154835, 0.1407755, 
    0.04033803, 0.01747169, 0.07193992, 0.144484, 0.09001714, 0.07294855, 
    0.08871447, 0.09296264, 0.1064415, 0.08112947, 0.03014783,
  0.08943113, 0.2137718, 0.2400316, 0.2129313, 0.1293192, 0.1229521, 
    0.06920575, 0.1434388, 0.186413, 0.1143464, 0.1174586, 0.1865312, 
    0.1596714, 0.1303034, 0.2103727, 0.2121407, 0.1674964, 0.2580653, 
    0.195639, 0.1231706, 0.1289135, 0.1691441, 0.2301816, 0.2216808, 
    0.2047087, 0.1439444, 0.1569551, 0.08782357, 0.06434597,
  0.2230064, 0.2595203, 0.2333462, 0.3829753, 0.3172706, 0.1807956, 
    0.1509895, 0.1762995, 0.222421, 0.2441747, 0.22392, 0.1202449, 0.2681418, 
    0.1692441, 0.2453304, 0.1980545, 0.1972844, 0.3589796, 0.2429402, 
    0.1078314, 0.2150286, 0.1634257, 0.2203051, 0.2404778, 0.3225369, 
    0.2887049, 0.1755353, 0.1415509, 0.2427512,
  0.252112, 0.3251451, 0.2350277, 0.4174662, 0.3803712, 0.3061988, 0.3436948, 
    0.3921725, 0.2820653, 0.3206735, 0.2503736, 0.3932255, 0.2097866, 
    0.2299448, 0.2348609, 0.2099327, 0.2427889, 0.2532895, 0.3366118, 
    0.3561207, 0.2557442, 0.1872349, 0.09959611, 0.2597009, 0.2065415, 
    0.3585636, 0.2798064, 0.2841064, 0.2713033,
  0.1134063, 0.1764052, 0.1786898, 0.2550933, 0.3253339, 0.213851, 0.2233144, 
    0.2391429, 0.194114, 0.119235, 0.07469492, 0.1211688, 0.1633931, 
    0.2249051, 0.2337404, 0.1763007, 0.1913059, 0.1305118, 0.1338796, 
    0.16221, 0.1899367, 0.2388884, 0.1800839, 0.2089432, 0.1754507, 
    0.1709962, 0.2004456, 0.1283518, 0.1735075,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0.01892745, -0.0002736447, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0003249375, 
    0.03343324, 0.2022903, 0.06019291, 0.07828751, 0.1267168, 0.1692871, 
    0.1230481, 0.1662823, 0.2948249, 0.3045217, 0.2973505, 0.344681, 
    0.318479, 0.2223142, 0.1751231, 0.1899797, 0.1242249,
  0.1796667, 0.1633549, 0.06701036, 0.1239841, 0.07143877, 0.1003931, 
    0.1852234, 0.04719172, 0.01177065, 0.06871068, 0.0350985, 0.0774217, 
    0.2138365, 0.2934926, 0.2737397, 0.2226857, 0.2752909, 0.2730152, 
    0.2924754, 0.2964639, 0.3702776, 0.3295942, 0.4401622, 0.5203707, 
    0.277199, 0.1829838, 0.2449753, 0.2680762, 0.2721312,
  0.2710001, 0.2745826, 0.3439331, 0.3095883, 0.2686895, 0.2345977, 
    0.1828122, 0.188311, 0.2747664, 0.2815188, 0.2471816, 0.2970274, 
    0.2871408, 0.2648641, 0.3022887, 0.237417, 0.2307162, 0.2497581, 
    0.2406022, 0.2805679, 0.2428584, 0.2481687, 0.2422604, 0.2648238, 
    0.1966979, 0.1661665, 0.1258203, 0.1793573, 0.1713231,
  0.1933365, 0.1674452, 0.1497879, 0.2127074, 0.1743665, 0.1329224, 
    0.1504426, 0.1897891, 0.2089986, 0.2212386, 0.173682, 0.1869967, 
    0.1321308, 0.1527978, 0.1223858, 0.126396, 0.1017173, 0.1085677, 
    0.1178053, 0.1194244, 0.1663197, 0.1853493, 0.1613369, 0.112751, 
    0.09889975, 0.1688186, 0.1502166, 0.1585535, 0.2041189,
  0.1433758, 0.09621223, 0.06120943, 0.07641877, 0.07616311, 0.1127527, 
    0.1108122, 0.1073634, 0.1180721, 0.04241569, 0.005523418, 0.007265112, 
    0.07697529, 0.09142736, 0.1707904, 0.05638304, 0.127585, 0.09370852, 
    0.09430101, 0.06086025, 0.07633007, 0.05672637, 0.07338979, 0.06420417, 
    0.08121189, 0.08343913, 0.1178238, 0.1036929, 0.1295158,
  5.924015e-05, 0.0001686594, 0.07531308, 0.1265935, 0.06718308, 0.0213976, 
    0.02539017, 0.003762453, 0.004706204, 0.002788706, 0.01524539, 
    0.03190148, 0.1183827, 0.06978273, 0.0464005, 0.02047052, 0.02163645, 
    0.009528951, 0.2214525, 0.2004043, 0.07150242, 0.006475471, 0.0001074298, 
    -1.331027e-06, 0.07052339, 0.03913743, 0.1194207, 0.07227218, 0.07071149,
  7.246041e-09, 0.04000694, 0.1556902, 0.003663647, 0.01721496, 5.790761e-05, 
    0.002962122, 0.001502388, 0.0001989541, 2.256849e-06, 0.1051411, 
    0.0231113, 0.01087379, 0.08059266, 0.04078348, 0.08374627, 0.1198216, 
    0.102149, 0.0349895, 0.03801918, -0.0002480864, 6.636182e-06, 
    3.453817e-08, -1.995959e-05, 0.07572588, 0.1429326, 0.09365249, 
    5.800886e-06, 1.935415e-06,
  0.0102564, 0.07571738, 0.1965511, 0.01940672, 0.03513971, 0.07962763, 
    0.06862851, 0.08003016, 0.0203684, 0.002160404, 0.01162417, 0.02421175, 
    0.07400887, 0.0230698, 0.135158, 0.1285589, 0.03851073, 0.01315583, 
    0.0006201724, 6.056217e-08, 1.161118e-07, 0.0001162621, 0.0001761613, 
    0.1813463, 0.1022631, 0.2650194, 3.329031e-05, 1.003097e-08, 6.635878e-06,
  0.09003644, 0.4408291, 0.2379155, 0.01019603, 0.001684384, 0.08104091, 
    0.05194597, 0.0370896, 0.1189499, 0.09262752, 0.01107434, 0.006295829, 
    0.01578945, 0.0519048, 0.02018092, 0.005232723, 0.0001473406, 
    0.002040741, -8.693893e-05, 4.421239e-05, 0.0005621782, 0.01280048, 
    0.08991863, 0.1031891, 0.02970269, 0.0007088786, 0.01712796, 0.009115919, 
    0.02961518,
  0.01797646, 0.009435204, 0.008279683, 0.0577623, 0.00807537, 0.002434191, 
    0.05766456, 0.05861291, 0.1985953, 0.04265477, 0.08641447, 0.1193519, 
    0.1583085, 0.287244, 0.07683874, 0.1330253, 0.1982456, 0.1368573, 
    0.1259361, 0.08221409, 0.1158992, 0.08430697, 0.1576, 0.05228263, 
    0.07446635, 0.1636497, 0.0425276, 0.02286288, 0.0136948,
  0.001140582, -5.608879e-09, -1.362897e-07, 0.001165222, -1.968875e-06, 
    2.050497e-05, 0.07767601, 0.1233865, 0.04596598, 0.0451297, 0.06111163, 
    0.1300846, 0.06836972, 0.07956077, 0.01989656, 0.03228489, 0.0153412, 
    0.004603917, 0.004472014, 0.06347633, 0.0310689, 0.150355, 0.01843116, 
    0.02836039, 0.01324137, 0.02369912, 0.01702351, 0.0163387, 4.668608e-05,
  0.0003124881, 0.009716035, 0.01922036, -9.090079e-05, 0.005601335, 
    6.243385e-07, 0.005221881, 0.1588384, 0.3611797, 0.03096645, 0.04787442, 
    0.04823487, 0.08361544, 0.01356031, 0.04616437, 0.03332729, 0.02603363, 
    0.02745329, 0.01769165, 0.002314666, 0.02117408, 0.07038838, 0.06281024, 
    0.03547718, 0.07170044, 0.04358758, 0.06661784, 0.007638929, 0.04875318,
  0.0385526, 0.03629297, 0.1263745, 0.09520835, 0.0728454, 0.01750679, 
    0.04012061, 0.01028186, 0.04093955, 0.05719819, 0.09373875, 0.1267005, 
    0.1421868, 0.1647222, 0.1559772, 0.1698888, 0.1648584, 0.1505252, 
    0.04674705, 0.01906551, 0.07762818, 0.1558843, 0.08725081, 0.07213935, 
    0.09559538, 0.1078643, 0.1173337, 0.08128458, 0.0263848,
  0.09484927, 0.2119211, 0.2362732, 0.1946508, 0.1417463, 0.121792, 
    0.07146893, 0.1399444, 0.1778786, 0.1033877, 0.1314164, 0.1819966, 
    0.1737727, 0.1473062, 0.1961199, 0.2380986, 0.1946959, 0.2531552, 
    0.1844516, 0.1296649, 0.1272158, 0.1650108, 0.2598642, 0.2189343, 
    0.2226658, 0.1489045, 0.1718067, 0.07985044, 0.06730319,
  0.1957811, 0.2626581, 0.2399072, 0.3812312, 0.3098792, 0.1803722, 
    0.1555025, 0.1507579, 0.1956748, 0.256723, 0.2279915, 0.1299134, 
    0.2902881, 0.2035062, 0.2796905, 0.2299547, 0.2099197, 0.3879491, 
    0.2445652, 0.09315459, 0.2028577, 0.150335, 0.2327966, 0.2726273, 
    0.2958383, 0.3325565, 0.1794088, 0.1488173, 0.2584856,
  0.2406438, 0.2983623, 0.2469256, 0.4262019, 0.3722429, 0.3263677, 
    0.3085745, 0.3668776, 0.2932993, 0.3160194, 0.2576529, 0.3494469, 
    0.2410283, 0.2285787, 0.2281085, 0.2429574, 0.2234083, 0.2559918, 
    0.3361355, 0.392915, 0.2338992, 0.1914726, 0.1135506, 0.226992, 
    0.2335165, 0.4014393, 0.3068853, 0.2816451, 0.2535129,
  0.1437229, 0.2173993, 0.2284497, 0.2494692, 0.2943382, 0.2429798, 
    0.2568892, 0.2553894, 0.220446, 0.09986687, 0.06066648, 0.09734177, 
    0.1536531, 0.181606, 0.191337, 0.1338971, 0.1317802, 0.09725792, 
    0.1049711, 0.1857442, 0.2032505, 0.256473, 0.1653556, 0.2023356, 
    0.1795681, 0.2138658, 0.1858638, 0.1358202, 0.1835787,
  0.0003883444, 0.0002716848, 0.0001550252, 3.836565e-05, -7.829392e-05, 
    -0.0001949535, -0.0003116131, 1.8472e-05, 3.510201e-05, 5.173203e-05, 
    6.836205e-05, 8.499206e-05, 0.0001016221, 0.0001182521, -0.00172944, 
    -0.001257739, -0.0007860369, -0.0003143351, 0.0001573666, 0.0006290684, 
    0.00110077, 0.001069778, 0.0006981054, 0.0003264332, -4.523903e-05, 
    -0.0004169112, -0.0007885835, -0.001160256, 0.000481672,
  0.1073103, -0.002577145, 0, 0, 0, 0, 0, 0, 0, 0, -0.0004111264, 0.02293323, 
    0.1313919, 0.2047112, 0.06027051, 0.07271164, 0.1162338, 0.1719283, 
    0.1052726, 0.1672231, 0.4194754, 0.5033332, 0.278521, 0.3520322, 
    0.3270951, 0.2185442, 0.1807716, 0.1844323, 0.2010997,
  0.1868028, 0.1562468, 0.0696363, 0.1215226, 0.1283072, 0.1302176, 
    0.2006351, 0.1045716, 0.1055372, 0.1605211, 0.145296, 0.1983785, 
    0.1995226, 0.2996737, 0.2944533, 0.2179013, 0.3053921, 0.2874266, 
    0.2977556, 0.3378297, 0.3878083, 0.3365311, 0.4553547, 0.5752064, 
    0.265335, 0.1981708, 0.2387356, 0.2578351, 0.2608948,
  0.2603263, 0.2573718, 0.3220458, 0.3114115, 0.2685185, 0.2521692, 
    0.1994514, 0.1957828, 0.3051796, 0.3186213, 0.2763502, 0.2873378, 
    0.2990509, 0.2753581, 0.3041978, 0.247015, 0.2262872, 0.2462944, 
    0.2483609, 0.2932527, 0.2854311, 0.2747415, 0.2384966, 0.2561396, 
    0.1967472, 0.141483, 0.1447533, 0.2070658, 0.146315,
  0.2002624, 0.1496743, 0.1531284, 0.222598, 0.1881277, 0.1605801, 0.166585, 
    0.2156802, 0.1899253, 0.2419585, 0.1935907, 0.1998703, 0.1379844, 
    0.1437588, 0.103768, 0.104729, 0.1217479, 0.1143843, 0.1331004, 
    0.1197342, 0.174104, 0.1793253, 0.1547743, 0.1263495, 0.1078291, 
    0.188782, 0.1612509, 0.1359998, 0.2048086,
  0.1425572, 0.1091571, 0.0646213, 0.07766982, 0.09197424, 0.1327694, 
    0.1059111, 0.1089011, 0.1142312, 0.02231871, 0.003983896, 0.01208632, 
    0.09482469, 0.09552986, 0.1803079, 0.049704, 0.1377318, 0.09715402, 
    0.1115246, 0.05825026, 0.07100523, 0.05562799, 0.06922219, 0.07443935, 
    0.07138387, 0.09581713, 0.1187567, 0.1097107, 0.1311785,
  -0.0003518644, 6.189153e-05, 0.09768374, 0.1002459, 0.07752229, 0.06499522, 
    0.03225506, 0.00957196, 0.00601001, 0.0001417868, 0.01026397, 0.01233215, 
    0.1161863, 0.07120714, 0.04012442, 0.02012146, 0.02799816, 0.01133102, 
    0.2300182, 0.2193131, 0.0700332, 0.004373077, 0.001279955, -2.156999e-06, 
    0.07666051, 0.0432927, 0.125423, 0.06752729, 0.06898352,
  1.272206e-07, 0.02626579, 0.1477758, 0.004698731, 0.01229542, 0.001526014, 
    0.00505636, -0.0005730169, -2.647029e-06, 9.27421e-06, 0.03873761, 
    0.006433072, 0.007677861, 0.08297134, 0.01275675, 0.06399089, 0.1096524, 
    0.09175681, 0.03950115, 0.04202814, 0.0001594328, 6.251266e-07, 
    4.054831e-08, -1.04599e-05, 0.08089696, 0.1569652, 0.07408898, 
    1.225547e-05, 9.770235e-07,
  0.00356171, 0.04224688, 0.2003452, 0.03173623, 0.05769379, 0.08251855, 
    0.07052211, 0.07278759, 0.02059879, 0.005247309, 0.01258089, 0.01726901, 
    0.0792407, 0.02582741, 0.1096264, 0.1265131, 0.04413662, 0.02583952, 
    0.002101031, 2.219356e-07, 2.179866e-05, 4.138126e-07, 2.351234e-05, 
    0.1156485, 0.04781817, 0.1832997, 6.62103e-05, 6.219625e-09, 0.0002598268,
  0.04103082, 0.4189194, 0.1383193, 0.01355583, 0.00193231, 0.07773045, 
    0.06611037, 0.02523654, 0.1299376, 0.09649672, 0.01053763, 0.004153282, 
    0.01445193, 0.04127656, 0.02059796, 0.002759601, 0.0001128051, 
    0.003313959, -2.723816e-05, 0.01353514, 0.04063272, 0.02725445, 
    0.06903259, 0.07180508, 0.1276279, 0.0009452623, 0.01163501, 0.004777262, 
    0.01248738,
  0.006993966, 0.002190976, 0.00773509, 0.2107761, 0.01462831, 0.005019031, 
    0.06647488, 0.05204141, 0.196873, 0.04542604, 0.08615987, 0.1101602, 
    0.1212614, 0.2305728, 0.06561368, 0.1300773, 0.1653205, 0.134701, 
    0.1283144, 0.0792296, 0.1109308, 0.08224837, 0.1541153, 0.04890539, 
    0.06998607, 0.1359089, 0.03149972, 0.008624293, 0.006731644,
  5.560528e-05, 1.393398e-06, 4.003012e-07, 0.0002670326, -5.384912e-05, 
    -6.012866e-06, 0.08135927, 0.09793735, 0.06728077, 0.04514771, 
    0.05670377, 0.1376321, 0.06189235, 0.06536725, 0.02502563, 0.03157086, 
    0.01446002, 0.004543138, 0.01400044, 0.05092722, 0.02575688, 0.1632124, 
    0.01699627, 0.024629, 0.01253762, 0.01622252, 0.00104203, 0.02234161, 
    1.841211e-05,
  0.0004191306, 0.009339887, 0.008924491, 0.002562007, 0.002002107, 
    2.225015e-06, 0.006497441, 0.1857759, 0.3539362, 0.009133613, 0.04678997, 
    0.04714448, 0.08908658, 0.01213152, 0.05012625, 0.03884539, 0.02916567, 
    0.02962681, 0.01833063, 0.0004212663, 0.0184228, 0.07006518, 0.04971508, 
    0.04092304, 0.06135252, 0.03046233, 0.05573135, 0.01262391, 0.02374702,
  0.02977329, 0.02462086, 0.1485175, 0.1366739, 0.06614133, 0.008555315, 
    0.04732845, 0.006225374, 0.035457, 0.04096968, 0.1141515, 0.1200236, 
    0.1530743, 0.1620109, 0.1547595, 0.1876232, 0.1733096, 0.1513011, 
    0.04400137, 0.01859339, 0.08622081, 0.1462058, 0.09234904, 0.07374352, 
    0.1126172, 0.1163448, 0.1509692, 0.08194271, 0.02974382,
  0.08624664, 0.212154, 0.260095, 0.1990362, 0.1414803, 0.1202517, 
    0.06396234, 0.1566196, 0.1598366, 0.1065501, 0.1638969, 0.1831918, 
    0.1730775, 0.1431197, 0.1864182, 0.2387281, 0.1818454, 0.2610452, 
    0.1865477, 0.1421485, 0.1425011, 0.1688926, 0.2438415, 0.209788, 
    0.2401806, 0.1552549, 0.1839666, 0.1013333, 0.06362513,
  0.1822578, 0.2599939, 0.2342439, 0.3479295, 0.2834106, 0.1729723, 
    0.1359097, 0.2023061, 0.2054227, 0.2931293, 0.2485423, 0.1629718, 
    0.3629795, 0.2559886, 0.2407323, 0.23293, 0.2667829, 0.4223594, 
    0.2940331, 0.07632264, 0.2129227, 0.1327633, 0.2019784, 0.2379963, 
    0.3056385, 0.3673775, 0.1687883, 0.1486968, 0.2427697,
  0.277393, 0.2948727, 0.2500991, 0.4460714, 0.4180157, 0.3490765, 0.2892903, 
    0.3622597, 0.2894063, 0.3605187, 0.2697627, 0.3397537, 0.2794001, 
    0.268184, 0.2733255, 0.2295657, 0.2157141, 0.258612, 0.3074429, 
    0.3320497, 0.3026544, 0.2741257, 0.1528991, 0.2427662, 0.1833993, 
    0.4446375, 0.318403, 0.2753558, 0.2648224,
  0.2315389, 0.336435, 0.3766279, 0.3490976, 0.3588778, 0.3119942, 0.3041086, 
    0.2836419, 0.2510874, 0.09784202, 0.0781611, 0.1108756, 0.1642131, 
    0.1893649, 0.2081612, 0.1336851, 0.1005723, 0.08731906, 0.08540093, 
    0.1737495, 0.2086109, 0.2757983, 0.2201378, 0.2046907, 0.1773944, 
    0.2177075, 0.1586405, 0.1733675, 0.2338191,
  0.008033142, 0.005041669, 0.002050196, -0.0009412768, -0.00393275, 
    -0.006924223, -0.009915696, 0.0003069507, 0.0005364316, 0.0007659124, 
    0.0009953931, 0.001224874, 0.001454355, 0.001683836, -0.0190103, 
    -0.01320823, -0.007406164, -0.001604097, 0.00419797, 0.01000004, 
    0.0158021, 0.02667755, 0.02363748, 0.02059741, 0.01755733, 0.01451726, 
    0.01147718, 0.008437107, 0.01042632,
  0.2343454, 0.003473091, -2.115594e-05, 0, 0, -1.032009e-05, 0, 0, 0, 0, 
    -0.001800288, 0.08884984, 0.2052138, 0.1960833, 0.07664896, 0.07151219, 
    0.1061553, 0.1603202, 0.1021945, 0.1587681, 0.4371289, 0.59123, 
    0.3227177, 0.3554611, 0.3292209, 0.1855456, 0.1912109, 0.1759536, 
    0.1998805,
  0.2005519, 0.1500974, 0.06986316, 0.1144917, 0.1597798, 0.1517484, 
    0.206652, 0.1818344, 0.2167354, 0.2230927, 0.2321753, 0.2072324, 
    0.1939328, 0.3023799, 0.2814614, 0.2366156, 0.3206004, 0.2749303, 
    0.2968497, 0.3169678, 0.3678926, 0.3261915, 0.4408718, 0.6244727, 
    0.2858095, 0.2038152, 0.2534519, 0.2761756, 0.2504491,
  0.2679082, 0.2985834, 0.3477685, 0.3318263, 0.2966085, 0.2520148, 
    0.2189207, 0.1982782, 0.305998, 0.3438063, 0.2903499, 0.2990516, 
    0.2874248, 0.3010649, 0.3104357, 0.2755579, 0.2781805, 0.2780017, 
    0.2552214, 0.3195238, 0.3098194, 0.2823827, 0.2530354, 0.2830128, 
    0.234542, 0.1864246, 0.1778135, 0.2233303, 0.1974941,
  0.2418248, 0.1694299, 0.1808011, 0.215422, 0.1998984, 0.1799636, 0.1846344, 
    0.2217184, 0.1885029, 0.2326481, 0.2282552, 0.2407065, 0.1735563, 
    0.1449585, 0.1017557, 0.105888, 0.1317079, 0.1484831, 0.1351779, 
    0.1509453, 0.1899598, 0.1792217, 0.1635834, 0.1463127, 0.1300122, 
    0.2159887, 0.18712, 0.1488976, 0.1957954,
  0.1570709, 0.1186437, 0.08040967, 0.08881778, 0.109104, 0.1440766, 
    0.1104358, 0.1245695, 0.1315452, 0.01475805, 0.02020206, 0.01716836, 
    0.1085186, 0.09651349, 0.1850343, 0.07458363, 0.1522967, 0.11309, 
    0.1304617, 0.07768025, 0.07423954, 0.0690162, 0.09691754, 0.09912129, 
    0.07980058, 0.1130473, 0.1146576, 0.1155592, 0.1298543,
  -0.0001132944, 9.887155e-05, 0.07489277, 0.07282854, 0.07890385, 
    0.08173861, 0.04305836, 0.007800989, 0.01015225, 3.482676e-05, 
    0.004549134, 0.009495773, 0.08592727, 0.0670796, 0.04573632, 0.01992586, 
    0.03856444, 0.01526997, 0.2502913, 0.2835881, 0.07626246, 0.00789571, 
    0.008218976, -8.727467e-07, 0.065404, 0.05042996, 0.1354245, 0.07181908, 
    0.1084808,
  2.058725e-07, 0.01216117, 0.04201499, 0.00489695, 0.01588993, 0.004577499, 
    0.007925802, -0.0004985817, -1.061326e-06, 7.86146e-07, 0.007356261, 
    0.001309585, 0.002848145, 0.08006343, 0.0085583, 0.05222948, 0.09002198, 
    0.07574757, 0.05579259, 0.05496596, 0.003484281, 9.74096e-08, 
    1.264688e-08, 1.904586e-06, 0.09027097, 0.1105329, 0.06266113, 
    -1.809608e-05, 2.959115e-07,
  0.0005536901, 0.02204257, 0.1388184, 0.06483806, 0.07327611, 0.09195661, 
    0.0594206, 0.07303014, 0.01689046, 0.005352691, 0.005532497, 0.01528974, 
    0.08593901, 0.02617964, 0.09988994, 0.1228579, 0.0542114, 0.03667168, 
    0.005769643, 0.0004639788, 8.784399e-08, 1.969502e-07, 4.972105e-06, 
    0.1034214, 0.03504092, 0.07215254, 0.0001864126, 1.318528e-09, 2.74476e-07,
  0.01937406, 0.3691401, 0.09305808, 0.03066709, 0.002244304, 0.0703377, 
    0.0671143, 0.02001666, 0.1253241, 0.1086928, 0.009034046, 0.004422589, 
    0.01357984, 0.03692234, 0.02290668, 0.003017498, 0.0005276892, 
    0.0003836901, 8.797834e-05, 0.006468577, 0.01245569, 0.01135645, 
    0.06322657, 0.06908228, 0.1810912, 0.0002100369, 0.008248184, 
    0.007554666, 0.006939507,
  0.001544013, 0.001200797, 0.005090313, 0.233589, 0.008720871, 0.01445775, 
    0.06812436, 0.04926871, 0.2028896, 0.05148333, 0.08106109, 0.1074914, 
    0.09985943, 0.1950261, 0.06712919, 0.1320718, 0.1382019, 0.1439552, 
    0.1431158, 0.08564961, 0.1110915, 0.0844819, 0.1573065, 0.0451143, 
    0.05905871, 0.1012738, 0.03465386, 0.007663111, 0.002634335,
  1.438988e-05, 3.50647e-07, -1.145359e-07, 0.0001771822, -1.620661e-06, 
    -1.142657e-06, 0.08911795, 0.08624613, 0.08475072, 0.05047572, 
    0.05777554, 0.1318946, 0.06190353, 0.05313739, 0.03215395, 0.03294145, 
    0.01394917, 0.01092171, 0.01267673, 0.03875089, 0.01965036, 0.1469902, 
    0.02040013, 0.0284904, 0.01502034, 0.01202075, 0.003570949, 0.004681654, 
    8.784634e-06,
  2.972122e-05, 0.01084907, 0.009898539, 0.007237297, 0.0003560929, 
    1.335143e-06, 0.005523299, 0.1962109, 0.3525368, 0.003574577, 0.04780462, 
    0.05697707, 0.08880098, 0.02060024, 0.06286029, 0.04390885, 0.03168934, 
    0.03158258, 0.01127676, 0.001138677, 0.01829039, 0.05813193, 0.04175191, 
    0.04463397, 0.05503255, 0.02769987, 0.05172575, 0.02395225, 0.00516626,
  0.02546594, 0.02770508, 0.1542556, 0.1383204, 0.05984717, 0.006198009, 
    0.06441692, 0.003644753, 0.0276155, 0.03922572, 0.1379128, 0.1227349, 
    0.1666491, 0.157123, 0.1526577, 0.1930477, 0.1800678, 0.1598303, 
    0.04255616, 0.02003168, 0.07051042, 0.1090924, 0.1006451, 0.08615595, 
    0.1142959, 0.09940173, 0.1706926, 0.08040617, 0.02963913,
  0.08896239, 0.2282852, 0.2505827, 0.1684628, 0.1525834, 0.1222643, 
    0.1081682, 0.1854267, 0.1479422, 0.1211546, 0.1637669, 0.203321, 
    0.1896652, 0.1633206, 0.1855704, 0.2502081, 0.1673848, 0.2700476, 
    0.1933731, 0.1665023, 0.148079, 0.1803363, 0.2845966, 0.2102067, 
    0.2442229, 0.1543238, 0.1898488, 0.1216136, 0.08876225,
  0.1861339, 0.2385842, 0.2577378, 0.380503, 0.3443672, 0.1867824, 0.18679, 
    0.1651028, 0.1959834, 0.2864085, 0.2836829, 0.162395, 0.3750811, 
    0.2585007, 0.2453413, 0.239239, 0.3399148, 0.466657, 0.3171687, 
    0.07411985, 0.1982546, 0.1239779, 0.2114089, 0.2510198, 0.317403, 
    0.3876628, 0.1729602, 0.168335, 0.2578957,
  0.3072746, 0.2902501, 0.2583767, 0.4626774, 0.3955397, 0.3712451, 
    0.3686036, 0.3728362, 0.3373352, 0.3959931, 0.2925304, 0.3726697, 
    0.2215332, 0.2622185, 0.2817943, 0.291171, 0.2461956, 0.2599517, 
    0.340997, 0.4002041, 0.3249669, 0.2645948, 0.1534409, 0.2453616, 
    0.2584301, 0.4750654, 0.3144051, 0.2965719, 0.2515425,
  0.1818312, 0.3135743, 0.3594033, 0.3452849, 0.395813, 0.3910703, 0.2716423, 
    0.388331, 0.221505, 0.2282968, 0.113408, 0.1607529, 0.1885801, 0.1664435, 
    0.1998668, 0.1797337, 0.1430792, 0.1766327, 0.2004664, 0.2154762, 
    0.2211827, 0.3401246, 0.1868007, 0.1970772, 0.1773635, 0.2015585, 
    0.1520052, 0.2109422, 0.2854687,
  0.07106643, 0.06676165, 0.06245687, 0.05815209, 0.05384731, 0.04954252, 
    0.04523774, 0.05715017, 0.06308861, 0.06902706, 0.0749655, 0.08090395, 
    0.08684239, 0.09278084, 0.08916681, 0.09805462, 0.1069424, 0.1158302, 
    0.124718, 0.1336059, 0.1424937, 0.105708, 0.09518655, 0.08466507, 
    0.0741436, 0.06362213, 0.05310066, 0.04257919, 0.07451025,
  0.2541608, 0.07001664, -9.697156e-05, 0, 0, -0.001131532, 0, 0, 0, 
    0.0001033403, 0.02391107, 0.1658704, 0.2840673, 0.1763867, 0.08598953, 
    0.06677085, 0.1072176, 0.1528744, 0.07957271, 0.1638199, 0.4658982, 
    0.6195655, 0.3675808, 0.3557436, 0.3240542, 0.2006285, 0.2167679, 
    0.179245, 0.1935792,
  0.2055891, 0.1294182, 0.05801182, 0.1021111, 0.1883152, 0.1634939, 
    0.2248554, 0.2611062, 0.2910879, 0.2566015, 0.2452841, 0.1940629, 
    0.1883986, 0.2990503, 0.2941987, 0.2116529, 0.3125109, 0.2617776, 
    0.3112907, 0.3061147, 0.346791, 0.3214716, 0.4352809, 0.5940281, 
    0.2929506, 0.1927835, 0.2290509, 0.2866909, 0.2718427,
  0.2589221, 0.2401396, 0.3263748, 0.357423, 0.3123949, 0.2607441, 0.2261719, 
    0.2059668, 0.3168064, 0.3531154, 0.2816631, 0.2899085, 0.2637693, 
    0.3023598, 0.3007577, 0.2826117, 0.2836781, 0.2823934, 0.2693931, 
    0.327641, 0.3164911, 0.2936004, 0.2686411, 0.2744521, 0.2366188, 
    0.1866349, 0.161176, 0.21401, 0.1903295,
  0.24452, 0.2103855, 0.1937125, 0.2243014, 0.2144119, 0.1909474, 0.1768927, 
    0.2205751, 0.2043301, 0.232786, 0.2317401, 0.2756421, 0.2138113, 
    0.1667424, 0.1002742, 0.120587, 0.1540066, 0.1611401, 0.1460441, 
    0.1645383, 0.2116078, 0.2029736, 0.1945806, 0.175411, 0.1350612, 
    0.2351532, 0.1963166, 0.1250746, 0.2138886,
  0.1848593, 0.1333682, 0.1169834, 0.1209925, 0.1375196, 0.1462306, 
    0.1241237, 0.1598496, 0.1529163, 0.01730622, 0.03458012, 0.04453555, 
    0.1171245, 0.1132143, 0.1951652, 0.08341663, 0.1666571, 0.1190588, 
    0.1277718, 0.07971714, 0.09258733, 0.08958088, 0.1207688, 0.1118262, 
    0.06286515, 0.1387242, 0.1217587, 0.1538804, 0.1701729,
  0.005054499, 0.001817932, 0.05105902, 0.06725267, 0.1001969, 0.1013289, 
    0.04816251, 0.01589733, 0.01875306, 8.426361e-05, 0.0005553348, 
    0.002465317, 0.07682408, 0.05560851, 0.06892084, 0.02088552, 0.04952773, 
    0.02916634, 0.239041, 0.2753054, 0.06888396, 0.04023788, 0.0128654, 
    6.106725e-07, 0.04910726, 0.05819241, 0.1324469, 0.06103367, 0.1256396,
  7.807804e-08, 0.005352132, 0.02111153, 0.004292796, 0.02977678, 0.01577222, 
    0.009283586, 0.0001101494, 0.0002021011, 3.779059e-07, 0.0005438274, 
    0.0004585782, 0.001796454, 0.0723963, 0.01086138, 0.04646385, 0.07816024, 
    0.06561106, 0.06704618, 0.06653477, 0.03438516, 0.001673154, 
    1.793912e-06, 8.872514e-06, 0.09059717, 0.06173659, 0.09870293, 
    -4.400191e-06, 3.654621e-07,
  0.0003773532, 0.01622433, 0.04677331, 0.08957081, 0.07479735, 0.09592284, 
    0.06190153, 0.07381374, 0.01689371, 0.00552683, 0.005518771, 0.01025083, 
    0.09196211, 0.02970098, 0.08644199, 0.1158308, 0.06162788, 0.04536073, 
    0.01675028, 0.004533887, 5.111734e-08, 1.231972e-07, 2.959922e-06, 
    0.0943305, 0.0278756, 0.0308014, 0.005022867, 1.257421e-08, 4.316222e-07,
  0.009890425, 0.3387438, 0.07202584, 0.06815542, 0.0024645, 0.06896357, 
    0.06673521, 0.02037962, 0.116896, 0.1332209, 0.009004313, 0.004703392, 
    0.013403, 0.03502483, 0.02370125, 0.008548904, 0.003373635, 0.0006059225, 
    0.0002644147, 0.001956562, 0.001075593, 0.008204469, 0.03820105, 
    0.06992349, 0.1070325, 0.0001714834, 0.007284329, 0.006024322, 0.001424851,
  0.0007863124, 0.0008817278, 0.00221841, 0.1363392, 0.005214427, 0.02872215, 
    0.07125538, 0.04494126, 0.1811737, 0.05450587, 0.08715615, 0.1081738, 
    0.08850871, 0.1746906, 0.06434695, 0.1270352, 0.1260001, 0.1510124, 
    0.1539173, 0.0937375, 0.1080423, 0.08935193, 0.1559444, 0.04397792, 
    0.05028566, 0.07512409, 0.03586638, 0.006534504, 0.001732116,
  5.305789e-06, 1.071643e-07, -0.0002063977, -1.659077e-05, -1.823802e-07, 
    -4.488887e-06, 0.09615165, 0.07962047, 0.09737469, 0.06183188, 
    0.06129815, 0.1327503, 0.06061634, 0.05924046, 0.03778636, 0.04406284, 
    0.02544328, 0.01889493, 0.01602876, 0.02074736, 0.01049501, 0.1554324, 
    0.02243439, 0.03046998, 0.0196893, 0.02577613, 0.01582349, 0.0004417491, 
    4.447415e-06,
  1.405261e-05, 0.0187938, 0.03199903, 0.01524212, 0.0004314788, 
    6.193587e-07, 0.003399797, 0.1438728, 0.3489392, 0.0009774866, 0.0520138, 
    0.08347935, 0.09819327, 0.03038331, 0.06498263, 0.05699398, 0.04685029, 
    0.04130243, 0.01313106, 0.002882301, 0.0153107, 0.05056316, 0.04151388, 
    0.05523672, 0.05807928, 0.02968695, 0.0571272, 0.01736706, 0.001381563,
  0.0157567, 0.03274505, 0.1620407, 0.157345, 0.05627827, 0.007139037, 
    0.06748279, 0.002338683, 0.01888096, 0.04088141, 0.1425917, 0.1281697, 
    0.1801343, 0.1587429, 0.1527165, 0.2049632, 0.1915525, 0.165473, 
    0.05451334, 0.01809519, 0.05691446, 0.08185855, 0.1088353, 0.09375466, 
    0.1120667, 0.1077187, 0.1841891, 0.08044244, 0.02806687,
  0.09239522, 0.2492977, 0.2561109, 0.1888631, 0.1649169, 0.1116002, 
    0.1007158, 0.2144497, 0.1481327, 0.1296438, 0.1495848, 0.2153443, 
    0.2328323, 0.186374, 0.2012088, 0.2717625, 0.1825411, 0.2838328, 
    0.2034231, 0.1815642, 0.1332363, 0.1676347, 0.3012352, 0.2468738, 
    0.2453266, 0.1544817, 0.1992943, 0.1468677, 0.1115122,
  0.2032995, 0.2377533, 0.2650135, 0.4237175, 0.3673889, 0.1869509, 
    0.1777079, 0.1706109, 0.1678744, 0.2741997, 0.2811125, 0.1465315, 
    0.3285248, 0.2509313, 0.2258973, 0.2429779, 0.3354311, 0.4974097, 
    0.3293504, 0.08794358, 0.2021676, 0.09438427, 0.2443401, 0.22699, 
    0.3189608, 0.3970134, 0.2018804, 0.1727444, 0.2773151,
  0.3331628, 0.3003361, 0.2873784, 0.4799301, 0.408717, 0.4080271, 0.3541346, 
    0.4024659, 0.3029446, 0.4002395, 0.2657869, 0.3936965, 0.2116307, 
    0.2809782, 0.2483266, 0.2883806, 0.2445219, 0.2554487, 0.3185082, 
    0.3871258, 0.2602478, 0.2119286, 0.1348483, 0.2567184, 0.3399212, 
    0.5074435, 0.3155248, 0.2917562, 0.245395,
  0.1836194, 0.2755211, 0.2890294, 0.3079635, 0.2964748, 0.3575291, 
    0.2823578, 0.3471926, 0.1461241, 0.1627865, 0.1337095, 0.1353605, 
    0.2404972, 0.2463203, 0.2446946, 0.2233582, 0.2121654, 0.1680239, 
    0.2293104, 0.2238169, 0.2651208, 0.346819, 0.1598502, 0.1836368, 
    0.1956918, 0.1982117, 0.1671943, 0.2316298, 0.2698003,
  0.09580622, 0.08998394, 0.08416166, 0.07833938, 0.0725171, 0.06669482, 
    0.06087254, 0.08773565, 0.1002438, 0.1127519, 0.12526, 0.1377681, 
    0.1502762, 0.1627843, 0.170484, 0.1815898, 0.1926955, 0.2038013, 
    0.2149071, 0.2260128, 0.2371186, 0.2258136, 0.208022, 0.1902304, 
    0.1724388, 0.1546472, 0.1368556, 0.119064, 0.100464,
  0.2487421, 0.1963657, -0.008412168, 0, -4.179243e-06, -0.002561631, 
    0.0004239451, 0, 0, 0.0006716727, 0.1103494, 0.2322884, 0.2968888, 
    0.1390616, 0.05313907, 0.1118373, 0.09008942, 0.1353903, 0.05860334, 
    0.1224708, 0.4948474, 0.6480134, 0.4269962, 0.3570498, 0.335813, 
    0.2129031, 0.2140544, 0.2001493, 0.1860136,
  0.2041278, 0.1127361, 0.05652396, 0.09880789, 0.2324906, 0.1718716, 
    0.2346215, 0.3144179, 0.3347572, 0.2745968, 0.2624646, 0.1761828, 
    0.1703453, 0.2790102, 0.2859225, 0.2118815, 0.2761486, 0.2587255, 
    0.2819094, 0.2912778, 0.3566248, 0.3472162, 0.3996562, 0.5365778, 
    0.2833109, 0.2192414, 0.2683852, 0.3019594, 0.2783074,
  0.1893695, 0.2300858, 0.3303252, 0.3497578, 0.3055487, 0.2959232, 
    0.2033745, 0.1993604, 0.3266849, 0.3719619, 0.3009973, 0.2839912, 
    0.260914, 0.2926251, 0.3144951, 0.303531, 0.2888981, 0.2809399, 
    0.2656566, 0.329887, 0.3198077, 0.3240311, 0.2871313, 0.2600944, 
    0.2026792, 0.128943, 0.1315002, 0.1969239, 0.135484,
  0.2114433, 0.1900954, 0.1963366, 0.2303365, 0.2341359, 0.1669654, 
    0.1737342, 0.2300147, 0.2230244, 0.2664841, 0.2505988, 0.2736523, 
    0.22118, 0.1703672, 0.09874431, 0.1446429, 0.1473266, 0.1749679, 
    0.1773434, 0.187046, 0.2434047, 0.2581695, 0.255515, 0.1732967, 
    0.08535764, 0.1729109, 0.2045921, 0.1176312, 0.2152946,
  0.2078141, 0.1555287, 0.1298381, 0.1424679, 0.153884, 0.1510192, 0.1442524, 
    0.1730148, 0.1832116, 0.04568832, 0.04075694, 0.06653824, 0.144794, 
    0.151232, 0.2446437, 0.1084094, 0.1648849, 0.1573769, 0.1370771, 
    0.09189665, 0.130208, 0.1423209, 0.1346918, 0.127221, 0.05142647, 
    0.1800762, 0.1510376, 0.1721897, 0.19915,
  0.01380572, 0.01170033, 0.02808945, 0.0635007, 0.10979, 0.107783, 
    0.06234799, 0.02721815, 0.03350951, 0.0007550159, -4.607443e-05, 
    0.0004220512, 0.06625049, 0.04888593, 0.07484695, 0.03116279, 0.05922028, 
    0.03495527, 0.2233495, 0.2456985, 0.08733264, 0.06018507, 0.02574211, 
    2.111984e-05, 0.04121467, 0.06871267, 0.1565224, 0.06957103, 0.1588156,
  1.635185e-07, 0.002297332, 0.01148137, 0.008683378, 0.03734996, 0.03992014, 
    0.009306052, 0.008169702, 0.005277565, 2.55789e-07, 0.0001190494, 
    7.72367e-05, 0.00589599, 0.08530698, 0.007231931, 0.03743891, 0.07420263, 
    0.05660175, 0.06553818, 0.07438239, 0.07050252, 0.02094198, 0.00089789, 
    8.953786e-06, 0.06896412, 0.05666633, 0.1216059, 0.006778099, 2.89937e-06,
  9.137902e-06, 0.01350609, 0.02189091, 0.07787573, 0.09694593, 0.1101919, 
    0.06531745, 0.07715002, 0.02594459, 0.00836252, 0.008184987, 0.008519408, 
    0.1002609, 0.03190433, 0.07040257, 0.09215105, 0.05382017, 0.04555744, 
    0.01519038, 0.006757007, -5.081477e-06, 1.298503e-07, 1.848847e-06, 
    0.08767835, 0.02442537, 0.01845752, 0.01752385, -8.577386e-09, 
    7.045095e-07,
  0.005613152, 0.297824, 0.05818786, 0.05986387, 0.004371492, 0.07073246, 
    0.06572086, 0.02034962, 0.09797145, 0.1489242, 0.0103375, 0.005756993, 
    0.01398392, 0.03082095, 0.02380002, 0.01180592, 0.008937881, 0.0016199, 
    0.002664759, 0.001185815, 0.001964853, 0.007963834, 0.02241516, 
    0.07081625, 0.05216735, 0.0003028585, 0.01278531, 0.005383075, 
    0.0004072107,
  0.0008372826, 0.0006872668, 0.001653802, 0.0631585, 0.009092538, 
    0.03114419, 0.07217859, 0.0407735, 0.1566622, 0.05729503, 0.09088805, 
    0.09381761, 0.06895793, 0.1445449, 0.0571142, 0.1129031, 0.1142209, 
    0.1507894, 0.1493753, 0.09020292, 0.114764, 0.0994701, 0.1583415, 
    0.04796001, 0.03923409, 0.05645459, 0.03641086, 0.00494647, 0.001579297,
  2.08018e-06, 3.11631e-08, 9.700258e-05, -2.291852e-05, -6.428411e-09, 
    -2.475334e-06, 0.09529813, 0.06859179, 0.08198921, 0.06802359, 
    0.07355462, 0.1298787, 0.06198639, 0.05839872, 0.03837324, 0.04513846, 
    0.04077901, 0.03959307, 0.01801159, 0.004303051, 0.006343659, 0.1746497, 
    0.02254712, 0.02897654, 0.01999124, 0.02475155, 0.01223978, 2.075573e-05, 
    1.347535e-06,
  6.666804e-06, 0.02746896, 0.05839728, 0.01185604, 0.0003105184, 
    2.478912e-07, 0.0009276383, 0.1120491, 0.3158238, 0.001336007, 
    0.07440363, 0.1011027, 0.1081697, 0.0456279, 0.06630176, 0.06780592, 
    0.05511101, 0.05939258, 0.009988296, 0.004262498, 0.01363001, 0.04742064, 
    0.03503038, 0.06473432, 0.05823054, 0.03691864, 0.08473072, 0.01908143, 
    0.0001262172,
  0.007835721, 0.0515408, 0.151945, 0.1714606, 0.04822763, 0.002374221, 
    0.05571909, 0.001625865, 0.01299175, 0.03679333, 0.1135151, 0.1464562, 
    0.1969759, 0.1948263, 0.1813961, 0.2307287, 0.223645, 0.1516034, 
    0.07876062, 0.02094716, 0.05320114, 0.07938882, 0.1122699, 0.1073692, 
    0.1363994, 0.1212296, 0.1908487, 0.08171289, 0.02630785,
  0.09498367, 0.3135594, 0.2715868, 0.2082236, 0.1628708, 0.1098012, 
    0.07222991, 0.2199797, 0.1542563, 0.1312958, 0.1517736, 0.2474231, 
    0.2515225, 0.2092167, 0.2439563, 0.2890649, 0.2170746, 0.2992751, 
    0.2020126, 0.2018769, 0.1403171, 0.1913712, 0.302246, 0.2798009, 0.23571, 
    0.1792423, 0.2186182, 0.1724626, 0.0903853,
  0.240771, 0.2250443, 0.2738588, 0.4260481, 0.3374254, 0.1968314, 0.1712453, 
    0.1461176, 0.1965129, 0.309833, 0.2956384, 0.1428794, 0.3455245, 
    0.2575265, 0.2025438, 0.2565015, 0.3843594, 0.4868943, 0.3382455, 
    0.101169, 0.1807581, 0.1032839, 0.2453898, 0.2170429, 0.3149461, 
    0.4229931, 0.2240638, 0.1940593, 0.2748457,
  0.3364154, 0.2953475, 0.2631681, 0.4547658, 0.400195, 0.4214958, 0.322791, 
    0.3655385, 0.2950226, 0.5040116, 0.302278, 0.3454234, 0.193199, 
    0.2368555, 0.2871168, 0.2964845, 0.2159103, 0.2095909, 0.2681319, 
    0.3791048, 0.2466516, 0.210462, 0.104662, 0.270191, 0.3359367, 0.5273154, 
    0.3386624, 0.292217, 0.2553897,
  0.1521691, 0.2449556, 0.2348691, 0.2594182, 0.2481385, 0.3055923, 
    0.2511705, 0.2856393, 0.1900342, 0.08934067, 0.2041398, 0.1365438, 
    0.1770231, 0.2262411, 0.2152329, 0.2013723, 0.208978, 0.1309649, 
    0.1406161, 0.2106219, 0.232131, 0.2934405, 0.1914981, 0.1552524, 
    0.2079078, 0.1959892, 0.1736387, 0.2401588, 0.2331402,
  0.1480571, 0.1438056, 0.1395542, 0.1353027, 0.1310512, 0.1267998, 
    0.1225483, 0.1466119, 0.1667297, 0.1868475, 0.2069653, 0.2270831, 
    0.2472009, 0.2673187, 0.3151876, 0.3210359, 0.3268841, 0.3327324, 
    0.3385807, 0.344429, 0.3502772, 0.27527, 0.2535554, 0.2318408, 0.2101261, 
    0.1884115, 0.1666969, 0.1449823, 0.1514582,
  0.2455886, 0.2686774, -0.001209284, -2.381544e-05, -0.0006754231, 
    0.007238225, -0.00120764, -0.0001902238, 0.0003241875, 0.05385225, 
    0.2284512, 0.2094644, 0.3006964, 0.09198166, 0.06841705, 0.1034365, 
    0.1018324, 0.1331667, 0.05940226, 0.1036837, 0.5056963, 0.6473947, 
    0.4926108, 0.3756419, 0.3321243, 0.1790822, 0.2098628, 0.2133397, 
    0.2019621,
  0.225356, 0.09755526, 0.04545339, 0.08785637, 0.2628232, 0.1896385, 
    0.2127615, 0.3435181, 0.3376505, 0.3063892, 0.2541762, 0.1640961, 
    0.1798879, 0.25179, 0.2745329, 0.2324908, 0.3206481, 0.2730847, 
    0.3227125, 0.3209195, 0.374798, 0.3030185, 0.4349777, 0.5460516, 
    0.2971504, 0.1922217, 0.2537155, 0.3173831, 0.2808924,
  0.2197812, 0.2803228, 0.335835, 0.3507554, 0.3448958, 0.3344653, 0.2657977, 
    0.2218472, 0.3355324, 0.3811195, 0.3260809, 0.3128378, 0.304519, 
    0.3119263, 0.3208589, 0.2842917, 0.3265246, 0.3499918, 0.3306192, 
    0.3438582, 0.3464465, 0.3457686, 0.3050504, 0.2558049, 0.1978104, 
    0.1485892, 0.1337868, 0.1848678, 0.1492963,
  0.2541446, 0.2358448, 0.2559304, 0.3192699, 0.2734903, 0.1816473, 
    0.1771857, 0.2529051, 0.2620488, 0.2888695, 0.2797763, 0.320599, 
    0.210958, 0.1719831, 0.1283053, 0.1814081, 0.1614728, 0.2125116, 
    0.2278643, 0.2621643, 0.3003148, 0.2910147, 0.2584193, 0.1584377, 
    0.06778434, 0.1626837, 0.2251464, 0.1372012, 0.2255978,
  0.2086832, 0.2052678, 0.1424596, 0.1886174, 0.1810599, 0.1974933, 
    0.1536823, 0.1862192, 0.2023796, 0.105644, 0.1029848, 0.0827988, 
    0.1610452, 0.1433441, 0.2489442, 0.116052, 0.1710813, 0.2100222, 
    0.2492134, 0.1628852, 0.193838, 0.1891803, 0.154323, 0.1240545, 
    0.07113571, 0.1993716, 0.2125851, 0.1954014, 0.2226698,
  0.03211809, 0.06557658, 0.01976925, 0.08557776, 0.1164704, 0.1220351, 
    0.08009044, 0.05239766, 0.03418478, 0.00448866, -0.000187071, 
    4.12101e-05, 0.05627082, 0.05943408, 0.08757143, 0.0520804, 0.07247013, 
    0.04325107, 0.2645957, 0.2398528, 0.08996056, 0.09825224, 0.06059324, 
    0.0001448789, 0.03971777, 0.09915222, 0.1902219, 0.0875522, 0.1889789,
  2.586257e-06, 0.0005723254, 0.005990225, 0.01321446, 0.03886469, 
    0.05603421, 0.03262964, 0.04331884, 0.01700041, -6.601759e-06, 
    5.386364e-05, 1.297432e-05, 0.006559279, 0.07717127, 0.01186909, 
    0.0318779, 0.06999902, 0.048864, 0.05839339, 0.05759675, 0.04834698, 
    0.1089883, 0.008033372, 5.121819e-06, 0.05671721, 0.04791007, 0.1332597, 
    0.04745274, 0.0005421222,
  1.067722e-06, 0.01411503, 0.0153618, 0.05626747, 0.09463296, 0.1017652, 
    0.05833018, 0.0830754, 0.02898126, 0.01162801, 0.01017327, 0.009172357, 
    0.1060247, 0.03238688, 0.05116395, 0.07334535, 0.04731724, 0.04314113, 
    0.01473836, 0.008169377, 0.001098689, 1.887263e-06, 7.260034e-07, 
    0.07948282, 0.02211832, 0.01221885, 0.03160514, 4.394691e-06, 2.435673e-06,
  0.004430531, 0.2573964, 0.05010802, 0.05115192, 0.005579442, 0.0675801, 
    0.05644453, 0.02043323, 0.08106481, 0.1700251, 0.01681487, 0.008119877, 
    0.0161176, 0.02556433, 0.02388954, 0.01404758, 0.009459315, 0.005371007, 
    0.008077037, 0.0005047191, 0.002792582, 0.01851568, 0.01890555, 
    0.0639703, 0.02401897, 0.0009639767, 0.01737457, 0.005976437, 0.0006688745,
  0.0008762667, 0.0004979398, 0.0006322856, 0.02031095, 0.01654766, 
    0.02476246, 0.07826465, 0.03490519, 0.1422601, 0.04949103, 0.08496824, 
    0.06544076, 0.05318562, 0.1184541, 0.04780244, 0.09268969, 0.09669397, 
    0.1324032, 0.1359539, 0.08115245, 0.1034654, 0.08843727, 0.1639869, 
    0.05896661, 0.03019405, 0.04173043, 0.03338838, 0.004243609, 0.001627362,
  1.062838e-06, 2.27033e-08, 0.0001097296, -6.103183e-05, -1.474481e-11, 
    0.01719347, 0.08590213, 0.06164267, 0.0934889, 0.09706622, 0.1060899, 
    0.1177292, 0.05830039, 0.04880382, 0.04981589, 0.04858991, 0.04888338, 
    0.09160237, 0.02260393, 0.004344882, 0.004709947, 0.2103955, 0.02528867, 
    0.02515724, 0.02359228, 0.02255582, 0.0115255, 1.162071e-05, 3.458274e-07,
  2.998837e-06, 0.02151969, 0.03977293, 0.004139778, 0.0001478291, 
    9.364999e-08, -0.0004001808, 0.08356215, 0.3012932, 0.003685394, 
    0.1569313, 0.100838, 0.119659, 0.07130183, 0.07494602, 0.07255433, 
    0.08821081, 0.08953815, 0.02506028, 0.01052801, 0.01529238, 0.04868307, 
    0.03334937, 0.07264623, 0.04927936, 0.04305646, 0.09164635, 0.02914972, 
    4.103745e-05,
  0.00556923, 0.07512647, 0.1397701, 0.1644741, 0.03913831, 0.0002583481, 
    0.05795145, 0.0002723957, 0.01118995, 0.02994418, 0.1240876, 0.145787, 
    0.2307548, 0.2275373, 0.2234844, 0.2888385, 0.2669479, 0.2074955, 
    0.106658, 0.02463841, 0.04351544, 0.08874562, 0.1398326, 0.1179341, 
    0.162746, 0.1249033, 0.1904027, 0.08916428, 0.02286002,
  0.1294901, 0.3661709, 0.2990049, 0.239486, 0.176785, 0.127792, 0.07503634, 
    0.234503, 0.1365946, 0.1134844, 0.1587483, 0.3057669, 0.3002127, 
    0.2569948, 0.3306819, 0.3614636, 0.2502941, 0.3028655, 0.2268714, 
    0.1998607, 0.1759178, 0.2313885, 0.349962, 0.3129401, 0.2480465, 
    0.237776, 0.2287283, 0.193257, 0.07805278,
  0.2761893, 0.214706, 0.2616217, 0.3879803, 0.3579459, 0.1749728, 0.1847698, 
    0.1617299, 0.197335, 0.3591489, 0.3723739, 0.1664713, 0.3661194, 
    0.2771439, 0.2788431, 0.3775952, 0.3756804, 0.4711447, 0.3123421, 
    0.07479021, 0.2272132, 0.1244257, 0.2479281, 0.2151153, 0.3490008, 
    0.4304968, 0.2636486, 0.215518, 0.3072036,
  0.3617587, 0.2956292, 0.267722, 0.4636491, 0.4069914, 0.3926715, 0.2934565, 
    0.427523, 0.31529, 0.4737158, 0.3369733, 0.3327093, 0.2104413, 0.2191294, 
    0.3155639, 0.2785622, 0.2336647, 0.1920145, 0.2467327, 0.4239451, 
    0.2836448, 0.2619842, 0.1986596, 0.2905144, 0.3952447, 0.5250599, 
    0.3257815, 0.302374, 0.3312753,
  0.1503021, 0.2382241, 0.2761872, 0.2129894, 0.2121737, 0.3021942, 
    0.3168629, 0.305247, 0.1833626, 0.1292973, 0.1731043, 0.1127865, 
    0.1610195, 0.2089942, 0.181309, 0.1562705, 0.1362883, 0.136401, 
    0.09982453, 0.1838441, 0.2270123, 0.2263454, 0.2026963, 0.1552875, 
    0.2048544, 0.2120544, 0.1947674, 0.2316216, 0.245227,
  0.1537506, 0.1504861, 0.1472215, 0.143957, 0.1406924, 0.1374279, 0.1341633, 
    0.1520905, 0.1772152, 0.2023398, 0.2274644, 0.252589, 0.2777137, 
    0.3028383, 0.3683217, 0.3682153, 0.368109, 0.3680026, 0.3678962, 
    0.3677899, 0.3676835, 0.2580721, 0.2363184, 0.2145647, 0.192811, 
    0.1710573, 0.1493035, 0.1275498, 0.1563622,
  0.2547307, 0.2704693, 0.09977525, -0.0001673625, 0.004401582, 0.03563887, 
    0.007072197, -0.0007674049, 0.001305092, 0.08558834, 0.279682, 0.2220322, 
    0.2925076, 0.0564118, 0.04452482, 0.06145627, 0.09590095, 0.1231163, 
    0.04992534, 0.1060204, 0.5441527, 0.7045745, 0.554491, 0.4051265, 0.3455, 
    0.2006269, 0.2296203, 0.2384897, 0.2242391,
  0.2215812, 0.09434689, 0.0480173, 0.05631582, 0.255478, 0.2211616, 
    0.1682837, 0.3507829, 0.3545669, 0.3141842, 0.2523654, 0.1642033, 
    0.1792939, 0.2221991, 0.2604554, 0.2138639, 0.3113552, 0.2884819, 
    0.3507099, 0.4457265, 0.3969286, 0.3321742, 0.4090879, 0.5635759, 
    0.3065377, 0.1751134, 0.2594665, 0.3391972, 0.3170777,
  0.3083803, 0.330451, 0.3949697, 0.4128684, 0.4455537, 0.3923557, 0.3135572, 
    0.2512802, 0.3482366, 0.3843624, 0.3043904, 0.3006073, 0.3291392, 
    0.3282691, 0.3161051, 0.2825436, 0.3607861, 0.3780724, 0.3315502, 
    0.3200433, 0.3329231, 0.2989328, 0.2845481, 0.2715591, 0.2163742, 
    0.224018, 0.1540688, 0.2171545, 0.1943376,
  0.322814, 0.4070578, 0.3309231, 0.3105649, 0.2648969, 0.2060845, 0.1868203, 
    0.255193, 0.2586256, 0.3118964, 0.298679, 0.3582887, 0.2610576, 
    0.1879244, 0.1836409, 0.2023363, 0.2143787, 0.2395059, 0.2622933, 
    0.2715395, 0.3277507, 0.2999583, 0.2497519, 0.1574018, 0.06060521, 
    0.2007318, 0.2450386, 0.1708559, 0.2679725,
  0.2597545, 0.2834422, 0.1836058, 0.2688752, 0.2376799, 0.2393677, 0.181002, 
    0.2183942, 0.2518676, 0.166388, 0.1602987, 0.1618174, 0.168286, 
    0.1399149, 0.2403953, 0.1940342, 0.3056286, 0.2898593, 0.298667, 
    0.1970768, 0.2663515, 0.1997973, 0.1861387, 0.1306597, 0.07527306, 
    0.2331334, 0.2491316, 0.2056545, 0.2755362,
  0.1638581, 0.1061212, 0.01677841, 0.1117889, 0.170293, 0.1791026, 
    0.0793215, 0.08764122, 0.06902143, 0.01239793, -0.0003491418, 
    3.741195e-05, 0.0332999, 0.0883968, 0.07994301, 0.06053337, 0.1134178, 
    0.07708112, 0.2848331, 0.2498787, 0.1781405, 0.1445642, 0.1670903, 
    0.0001685337, 0.04774565, 0.1345337, 0.2795795, 0.1384711, 0.2393661,
  0.001673824, 0.0002997452, 0.003682522, 0.02086116, 0.04677087, 0.0595947, 
    0.1454091, 0.1302172, 0.134386, -1.679623e-05, 2.138565e-05, 
    2.073474e-06, 0.03258996, 0.06807825, 0.02638044, 0.03337976, 0.0759767, 
    0.04127894, 0.05873956, 0.04924905, 0.0757833, 0.2674701, 0.1103771, 
    7.50567e-06, 0.06732117, 0.05599197, 0.1321002, 0.1283615, 0.04515053,
  5.602201e-06, 0.0142318, 0.01189986, 0.03493234, 0.08530115, 0.07966656, 
    0.05483658, 0.07850568, 0.04331464, 0.01559156, 0.01102062, 0.01692491, 
    0.108386, 0.03571742, 0.03659864, 0.06463598, 0.04383127, 0.0375786, 
    0.0183279, 0.01875309, 0.02485171, 0.003271382, 3.206005e-06, 0.07178318, 
    0.0188667, 0.005796834, 0.06711692, 0.007256943, 0.000107044,
  0.02012306, 0.2433217, 0.04489433, 0.047065, 0.009775924, 0.0633862, 
    0.05256741, 0.02081715, 0.07450057, 0.1927894, 0.02239442, 0.01057724, 
    0.02072421, 0.02273771, 0.02835488, 0.02232664, 0.01240731, 0.01116572, 
    0.01840965, 0.01090432, 0.002329576, 0.009714991, 0.02454595, 0.05585836, 
    0.01143325, 0.006428488, 0.02620151, 0.01094759, 0.004945635,
  0.0005391045, 0.0002958229, 0.0002239314, 0.004847963, 0.02242259, 
    0.03100831, 0.08255092, 0.03467937, 0.1276591, 0.0481706, 0.07618643, 
    0.06666944, 0.04305079, 0.1070023, 0.04069878, 0.07788481, 0.07959152, 
    0.107347, 0.1189057, 0.07624203, 0.08967756, 0.07467096, 0.1706716, 
    0.05511884, 0.028525, 0.03870676, 0.03463763, 0.004841855, 0.0008703788,
  6.728139e-07, 1.874682e-08, 4.694075e-06, -2.808801e-05, 1.158848e-10, 
    0.004268451, 0.06905279, 0.05895206, 0.1015832, 0.1622117, 0.09114455, 
    0.1059504, 0.05347556, 0.04909515, 0.04733913, 0.05627249, 0.05747157, 
    0.09349817, 0.08181904, 0.01713841, 0.004460006, 0.2236969, 0.03646773, 
    0.02381131, 0.03037924, 0.0320869, 0.02218266, -1.161144e-05, 1.715843e-07,
  1.469676e-06, 0.007698518, 0.0404891, 0.0003138013, 4.577018e-05, 
    4.116137e-08, -0.0006948098, 0.06702614, 0.3269471, 0.008350707, 
    0.2525879, 0.1620338, 0.1828169, 0.09803097, 0.1350869, 0.08966509, 
    0.0962721, 0.09997012, 0.08512726, 0.008326967, 0.01161178, 0.04837586, 
    0.04710461, 0.1055628, 0.06106708, 0.05377984, 0.104396, 0.03042696, 
    1.744267e-05,
  0.01261257, 0.06790657, 0.1231457, 0.1819968, 0.05962466, -0.0001107551, 
    0.05771774, 2.322984e-05, 0.01753673, 0.02410809, 0.1252885, 0.1444833, 
    0.2620185, 0.280986, 0.3299882, 0.3213436, 0.2992682, 0.2582639, 
    0.1711176, 0.02677135, 0.03045243, 0.1122401, 0.126672, 0.1471372, 
    0.2166196, 0.1455236, 0.1942392, 0.09036396, 0.01730935,
  0.170137, 0.3728346, 0.3156927, 0.2768051, 0.1744633, 0.1092495, 
    0.09726442, 0.278349, 0.1576932, 0.1085302, 0.1166878, 0.307015, 
    0.3729488, 0.378754, 0.3732667, 0.3706107, 0.2818362, 0.3284095, 
    0.264394, 0.1769002, 0.1763464, 0.2345984, 0.3447437, 0.3191666, 
    0.2798522, 0.297261, 0.2645864, 0.2176918, 0.1291599,
  0.3575826, 0.1970774, 0.2853845, 0.4154471, 0.4008621, 0.1692117, 0.195179, 
    0.2379525, 0.271718, 0.4268676, 0.3850029, 0.2237663, 0.3306712, 
    0.3544169, 0.4560688, 0.4972229, 0.4006811, 0.4657325, 0.329521, 
    0.09199747, 0.308307, 0.2037031, 0.2856406, 0.2781504, 0.3893506, 
    0.4096875, 0.2958859, 0.2991681, 0.3565691,
  0.3394549, 0.2545694, 0.34938, 0.4213496, 0.4127973, 0.4138266, 0.3246461, 
    0.4575399, 0.3294088, 0.5039181, 0.3974345, 0.3479205, 0.2093898, 
    0.2782907, 0.3109113, 0.257823, 0.231915, 0.2280668, 0.3092688, 
    0.4523254, 0.3282985, 0.3374484, 0.3591423, 0.2929674, 0.3728029, 
    0.5256091, 0.3245422, 0.2650708, 0.479742,
  0.1582853, 0.2407654, 0.2923999, 0.2097169, 0.3465958, 0.4168252, 
    0.4899644, 0.3726155, 0.2634816, 0.1299478, 0.1479324, 0.1391359, 
    0.1689944, 0.2114095, 0.2012508, 0.1441842, 0.1289223, 0.1995848, 
    0.1720588, 0.2393058, 0.2405953, 0.2708275, 0.1868805, 0.178893, 
    0.2208684, 0.2190777, 0.2199566, 0.2581587, 0.2930642,
  0.1418939, 0.1407577, 0.1396215, 0.1384853, 0.1373491, 0.1362129, 
    0.1350767, 0.1518921, 0.1761358, 0.2003795, 0.2246232, 0.2488669, 
    0.2731106, 0.2973543, 0.3475796, 0.3437681, 0.3399567, 0.3361453, 
    0.3323338, 0.3285224, 0.3247109, 0.2391396, 0.2198436, 0.2005475, 
    0.1812515, 0.1619555, 0.1426594, 0.1233634, 0.1428028,
  0.2596151, 0.275584, 0.1314534, -0.0006528808, 0.0207417, 0.06824689, 
    0.02734991, -0.001642398, 0.01794983, 0.1234756, 0.2894039, 0.2474974, 
    0.2803645, 0.02710425, 0.03998328, 0.0563242, 0.09523909, 0.09749609, 
    0.04028799, 0.08980345, 0.5917917, 0.713694, 0.6050204, 0.3638094, 
    0.3346069, 0.1966214, 0.2422668, 0.2833096, 0.2481836,
  0.2340681, 0.09155261, 0.05116142, 0.0279093, 0.2314721, 0.2510308, 
    0.1082578, 0.3629832, 0.3488615, 0.3210222, 0.2659618, 0.1653399, 
    0.158933, 0.1926399, 0.2583608, 0.2096892, 0.2930034, 0.3344571, 
    0.3570498, 0.439543, 0.4413343, 0.3876741, 0.4187269, 0.5830541, 
    0.3009137, 0.2024303, 0.3031322, 0.3943957, 0.3838835,
  0.3740248, 0.3737338, 0.4522081, 0.5020847, 0.5121489, 0.465649, 0.3073156, 
    0.3322541, 0.3602986, 0.3558046, 0.3073237, 0.2577825, 0.3572135, 
    0.3522843, 0.3237309, 0.29445, 0.3640338, 0.3699994, 0.314391, 0.3132963, 
    0.307138, 0.2554072, 0.2568034, 0.2763437, 0.2735195, 0.2875384, 
    0.256851, 0.2910435, 0.2883987,
  0.4498899, 0.4700688, 0.4169709, 0.3470459, 0.2959675, 0.2143303, 
    0.2460617, 0.3047595, 0.3330748, 0.3682738, 0.3024723, 0.3016291, 
    0.2699603, 0.2509082, 0.222659, 0.275258, 0.2770306, 0.3148953, 
    0.3548051, 0.3270107, 0.3087847, 0.3338576, 0.2808139, 0.1781565, 
    0.07506416, 0.296161, 0.3509966, 0.2054689, 0.372396,
  0.2959245, 0.2728106, 0.154966, 0.2652552, 0.2577944, 0.2423199, 0.2524694, 
    0.3337273, 0.3719311, 0.2230715, 0.1907607, 0.1406807, 0.1338962, 
    0.1608482, 0.2189865, 0.2467427, 0.3509808, 0.276697, 0.301722, 
    0.2853466, 0.3222744, 0.212973, 0.221541, 0.1339318, 0.04208482, 
    0.2029852, 0.2433838, 0.2264803, 0.3099445,
  0.3021685, 0.07688748, 0.01478514, 0.1465643, 0.173738, 0.1652129, 
    0.1790631, 0.1463005, 0.1631085, 0.05420151, 0.002787594, 5.037091e-05, 
    0.02586789, 0.112822, 0.1382269, 0.1275392, 0.2266825, 0.1385753, 
    0.3135432, 0.2455682, 0.170877, 0.1526952, 0.2003866, 0.001560152, 
    0.05325586, 0.1620917, 0.2459951, 0.1654647, 0.2980592,
  0.2427641, 0.0002028766, 0.001129695, 0.02567628, 0.05379147, 0.06462133, 
    0.1675171, 0.2251486, 0.3053853, 0.01348699, 8.687418e-06, 2.854601e-09, 
    0.1039564, 0.130947, 0.06072894, 0.07785788, 0.07555719, 0.0681157, 
    0.06771154, 0.06671124, 0.0986217, 0.4055285, 0.2487151, -3.900853e-06, 
    0.1151351, 0.07565895, 0.1329306, 0.1825563, 0.3451368,
  0.003056635, 0.007397712, 0.009025648, 0.02721991, 0.06679688, 0.0696459, 
    0.06332523, 0.1434275, 0.07281189, 0.02258343, 0.01479063, 0.02130788, 
    0.1369002, 0.05221328, 0.03501399, 0.06124838, 0.06696684, 0.06772482, 
    0.0505482, 0.04644259, 0.1285145, 0.07302666, -1.359757e-05, 0.06042551, 
    0.01444706, 0.001465315, 0.09454051, 0.06180989, 0.01069834,
  0.05142736, 0.2268483, 0.03337752, 0.03369226, 0.02377971, 0.06872961, 
    0.05553976, 0.02568373, 0.07130808, 0.2000558, 0.0791443, 0.01715233, 
    0.03540426, 0.02530047, 0.04264219, 0.06271017, 0.02570295, 0.008167899, 
    0.02168893, 0.0531848, 0.006694889, 0.004764626, 0.01061083, 0.04339459, 
    0.005660663, 0.01858042, 0.04476568, 0.02772191, 0.01151993,
  0.0001980483, 0.0001393668, 9.688153e-05, 0.0008069513, 0.02059192, 
    0.0806332, 0.09106222, 0.04306375, 0.1338571, 0.0551817, 0.06308374, 
    0.08795387, 0.04755138, 0.1032819, 0.04319899, 0.06822116, 0.0698295, 
    0.09416474, 0.1108218, 0.07319684, 0.08374824, 0.06841768, 0.1667652, 
    0.06249807, 0.03551384, 0.04224608, 0.03975311, 0.01000549, 0.0002465569,
  4.781259e-07, 1.848101e-08, 9.927337e-09, 0.001129253, 1.401743e-10, 
    -8.594683e-05, 0.04909371, 0.05911097, 0.1133291, 0.208743, 0.08028416, 
    0.1008784, 0.05415105, 0.06029647, 0.07128463, 0.07056586, 0.07989995, 
    0.09774842, 0.146265, 0.05681346, 0.02408752, 0.2230722, 0.06577431, 
    0.02937005, 0.04864212, 0.05484726, 0.05890442, 0.006263537, 1.309499e-07,
  7.445348e-07, 0.006406981, 0.03368009, -2.560847e-07, -4.045046e-05, 
    2.286245e-08, -0.0006448093, 0.05670619, 0.3312184, 0.008113743, 
    0.1540964, 0.1119659, 0.2181274, 0.1548362, 0.2107939, 0.1635297, 
    0.1176375, 0.1232172, 0.2175541, 0.01856126, 0.006014052, 0.04781221, 
    0.06301682, 0.0866388, 0.08320548, 0.09474657, 0.1127695, 0.04246156, 
    2.014545e-05,
  0.02263366, 0.02175288, 0.09981329, 0.2046735, 0.04624782, 0.0004839229, 
    0.04920697, -3.945802e-05, 0.02151292, 0.01645771, 0.1220433, 0.1525029, 
    0.2985244, 0.3792609, 0.3645859, 0.3136494, 0.2881918, 0.2319368, 
    0.2252095, 0.02103882, 0.02392183, 0.08665071, 0.1659999, 0.1157363, 
    0.1821742, 0.208099, 0.2042443, 0.1245921, 0.01792265,
  0.2540301, 0.3743815, 0.3005454, 0.2588294, 0.1411503, 0.09615201, 
    0.1126764, 0.2836967, 0.1414255, 0.09275264, 0.1035118, 0.3166149, 
    0.4017346, 0.3913144, 0.3496617, 0.3741243, 0.2812862, 0.3163815, 
    0.2811972, 0.1852825, 0.1688707, 0.214234, 0.3479461, 0.3214722, 
    0.2993822, 0.3969805, 0.3424951, 0.3662232, 0.245162,
  0.3273711, 0.185457, 0.3010062, 0.4264089, 0.381663, 0.2016509, 0.2355416, 
    0.3050215, 0.3306461, 0.4210538, 0.4366648, 0.2816746, 0.2974367, 
    0.3514513, 0.6202184, 0.4209546, 0.4479917, 0.4683407, 0.3991514, 
    0.1205799, 0.2872577, 0.261765, 0.2388644, 0.3335678, 0.4228613, 
    0.3787251, 0.3420627, 0.3192032, 0.3445896,
  0.2992081, 0.1828321, 0.3557302, 0.3702007, 0.4119249, 0.4428854, 
    0.4626154, 0.4875593, 0.3837807, 0.4223191, 0.4401932, 0.4164867, 
    0.2116679, 0.2993145, 0.311881, 0.290703, 0.3110913, 0.3298518, 
    0.3424547, 0.474332, 0.4642889, 0.3349722, 0.3064412, 0.2982697, 
    0.3015398, 0.5450065, 0.3069139, 0.262108, 0.3765111,
  0.2888272, 0.2892714, 0.3228789, 0.2615552, 0.4435863, 0.4884493, 0.511293, 
    0.4648416, 0.4130595, 0.3243386, 0.2102235, 0.1997993, 0.1811985, 
    0.1956259, 0.2178066, 0.1796246, 0.1676306, 0.2164719, 0.2249618, 
    0.2850598, 0.320517, 0.3108763, 0.1919831, 0.2252164, 0.2176072, 
    0.2212821, 0.2255686, 0.277814, 0.3628593,
  0.1262513, 0.1254863, 0.1247213, 0.1239564, 0.1231914, 0.1224264, 
    0.1216614, 0.142972, 0.1670952, 0.1912185, 0.2153418, 0.239465, 
    0.2635883, 0.2877116, 0.3260635, 0.3188774, 0.3116913, 0.3045053, 
    0.2973192, 0.2901332, 0.2829471, 0.2090539, 0.1928817, 0.1767095, 
    0.1605373, 0.1443651, 0.1281929, 0.1120206, 0.1268633,
  0.281264, 0.2809329, 0.1686208, -0.0008395698, 0.03305781, 0.0864804, 
    0.04930173, -0.00275325, 0.03150155, 0.1598093, 0.282005, 0.2817313, 
    0.2679362, 0.01240965, 0.03087528, 0.04426314, 0.08566971, 0.07945448, 
    0.03669596, 0.06887218, 0.6283323, 0.7383608, 0.5972399, 0.3072329, 
    0.3292884, 0.1996309, 0.2361692, 0.2856682, 0.2929522,
  0.2321722, 0.0754426, 0.0509559, 0.01321925, 0.1866232, 0.2444951, 
    0.05434056, 0.3539909, 0.3315383, 0.3123146, 0.2634378, 0.1694382, 
    0.1149643, 0.1646831, 0.2654914, 0.2584646, 0.3222389, 0.3754754, 
    0.4057647, 0.3845602, 0.4561057, 0.3528927, 0.4058206, 0.5883167, 
    0.2994032, 0.2508065, 0.4036206, 0.4500234, 0.4074036,
  0.416218, 0.4149694, 0.5253346, 0.5457556, 0.4688865, 0.4797953, 0.3396311, 
    0.3764026, 0.390067, 0.3221506, 0.2466793, 0.2454094, 0.357686, 
    0.3424044, 0.3209235, 0.3074346, 0.3564457, 0.373152, 0.377735, 
    0.2961664, 0.2589032, 0.2316533, 0.2392532, 0.2970669, 0.3067977, 
    0.3038625, 0.3386987, 0.375685, 0.4459119,
  0.4954306, 0.4831595, 0.4459847, 0.4009444, 0.3856152, 0.348577, 0.3296631, 
    0.3106308, 0.3398455, 0.3809679, 0.2858422, 0.2620604, 0.2451129, 
    0.2362633, 0.196426, 0.3188309, 0.307114, 0.4214389, 0.4392955, 
    0.3979094, 0.3245402, 0.2886484, 0.286883, 0.1888606, 0.08030386, 
    0.3359765, 0.4709816, 0.2970147, 0.4785114,
  0.2633393, 0.1875447, 0.1193609, 0.2329767, 0.201577, 0.1896466, 0.2658475, 
    0.376058, 0.3497838, 0.2380908, 0.1565684, 0.1368926, 0.1028687, 
    0.2119189, 0.2238617, 0.3451373, 0.3522053, 0.3525381, 0.3236624, 
    0.2295677, 0.2041612, 0.173442, 0.2382738, 0.1617, 0.02394326, 0.1731095, 
    0.2251894, 0.2411539, 0.2310638,
  0.2878446, 0.06656194, 0.01454919, 0.1327518, 0.1535307, 0.1434748, 
    0.281556, 0.3894759, 0.235637, 0.0383796, 0.01041963, 4.954677e-05, 
    0.01680834, 0.1406655, 0.1890579, 0.2259957, 0.1971609, 0.2006374, 
    0.3214973, 0.2178577, 0.1137645, 0.1204127, 0.1630546, 0.0003897764, 
    0.04084611, 0.2051637, 0.1834644, 0.1072348, 0.2447727,
  0.3867689, -0.0003264207, 0.0002224116, 0.06096238, 0.1011498, 0.03938981, 
    0.08288991, 0.1372005, 0.2033479, 0.03922818, 4.701734e-06, -1.04425e-07, 
    0.09659999, 0.1524021, 0.05666856, 0.1010718, 0.09173286, 0.07214441, 
    0.1022242, 0.045625, 0.06813633, 0.251471, 0.4181249, -0.0001205565, 
    0.1111366, 0.07046348, 0.1672899, 0.1452938, 0.4247722,
  0.05675582, 0.01493659, 0.004624462, 0.02268454, 0.07503732, 0.08721844, 
    0.08142453, 0.1123796, 0.1083147, 0.07911913, 0.01820607, 0.05934196, 
    0.1443287, 0.05840975, 0.04280965, 0.06958094, 0.0791737, 0.06772472, 
    0.1024472, 0.06956788, 0.1460125, 0.5041195, 0.04600662, 0.0401178, 
    0.008604634, 0.0004568554, 0.1390088, 0.3267561, 0.244331,
  0.08640535, 0.1929008, 0.02005846, 0.02910979, 0.09151052, 0.2319116, 
    0.05829677, 0.04072286, 0.05589421, 0.1433832, 0.1047365, 0.1377853, 
    0.1270628, 0.03741123, 0.05957368, 0.09725229, 0.03543748, 0.01580557, 
    0.03182489, 0.05150675, 0.07382289, 0.02651784, 0.04704492, 0.02792775, 
    0.002102026, 0.09584372, 0.06202701, 0.107003, 0.02811984,
  8.64212e-05, 5.947427e-05, 3.937808e-05, 7.7864e-05, 0.01876373, 0.1449383, 
    0.1033482, 0.07184133, 0.134269, 0.06470714, 0.04830348, 0.07408269, 
    0.06457011, 0.0936124, 0.05812404, 0.06763227, 0.07338677, 0.1138688, 
    0.1310726, 0.09682398, 0.1350843, 0.07020564, 0.2395576, 0.07745191, 
    0.1100651, 0.05001027, 0.07746711, 0.0722974, 0.0001695923,
  3.685437e-07, 1.803403e-08, -3.01815e-08, 0.003251413, 1.383667e-10, 
    -0.0002093453, 0.03663626, 0.1444052, 0.06787053, 0.1274273, 0.04660275, 
    0.08471205, 0.08452109, 0.05252502, 0.04927764, 0.05309227, 0.08950641, 
    0.08577768, 0.1528452, 0.2082084, 0.07320476, 0.2134815, 0.1037001, 
    0.05704906, 0.06052764, 0.09772208, 0.1322634, 0.05177004, 1.175448e-07,
  3.794488e-07, 0.01241479, 0.006813716, -5.734691e-05, -0.0001398057, 
    1.320588e-08, -0.0004639978, 0.05308489, 0.3133571, 0.0007779046, 
    0.1534772, 0.1008812, 0.1941554, 0.130529, 0.1393659, 0.1523598, 
    0.08983366, 0.1388254, 0.237137, 0.01011193, 0.004591044, 0.03990781, 
    0.05027071, 0.05514806, 0.04816038, 0.06148099, 0.112217, 0.1039296, 
    0.0002250578,
  0.04651498, 0.0192902, 0.09613105, 0.2175601, 0.03158937, 0.004308937, 
    0.04976097, 0.0001568326, 0.0172155, 0.01542048, 0.1204363, 0.1238699, 
    0.2505784, 0.3640004, 0.2851741, 0.300687, 0.2945513, 0.3040726, 
    0.3005274, 0.01533422, 0.01771191, 0.06727226, 0.1858481, 0.09327057, 
    0.1390856, 0.1778669, 0.2049513, 0.1300807, 0.01976193,
  0.3112333, 0.3693408, 0.3317212, 0.2753825, 0.1415528, 0.1202425, 
    0.1146822, 0.2535687, 0.1290274, 0.09088664, 0.09000178, 0.3851289, 
    0.3975229, 0.3173583, 0.322888, 0.3607259, 0.2651635, 0.3173814, 
    0.2893191, 0.2051966, 0.1665631, 0.1765473, 0.3335151, 0.3297684, 
    0.2747853, 0.3809072, 0.4317119, 0.4056252, 0.3494697,
  0.2537734, 0.1943596, 0.31829, 0.5081378, 0.4132102, 0.1746762, 0.2833133, 
    0.3057583, 0.4104477, 0.4294289, 0.4224874, 0.3913308, 0.3242134, 
    0.4174907, 0.4770484, 0.2910586, 0.472712, 0.4765807, 0.3919495, 
    0.08661609, 0.3061453, 0.3313624, 0.2544137, 0.4608922, 0.4856071, 
    0.3663719, 0.335646, 0.3437485, 0.374557,
  0.2232039, 0.1252001, 0.2760906, 0.3201144, 0.417403, 0.4391684, 0.5452539, 
    0.5421788, 0.39589, 0.4309288, 0.4787112, 0.4452136, 0.3076344, 
    0.3085313, 0.2771995, 0.4085956, 0.3846878, 0.3961644, 0.4363469, 
    0.4850636, 0.4503395, 0.3570392, 0.2811875, 0.366447, 0.274532, 
    0.6167458, 0.3055777, 0.246185, 0.3155611,
  0.3482069, 0.3423001, 0.3298505, 0.2994476, 0.4325116, 0.4608034, 
    0.4801421, 0.508233, 0.3178972, 0.5094576, 0.3153457, 0.2829163, 
    0.2404139, 0.2245121, 0.2557255, 0.2301444, 0.2513123, 0.2658876, 
    0.2883847, 0.3353803, 0.3872375, 0.3078391, 0.252879, 0.2628258, 
    0.2261921, 0.2257782, 0.262455, 0.3146373, 0.3375142,
  0.1132192, 0.1117519, 0.1102847, 0.1088174, 0.1073502, 0.1058829, 
    0.1044157, 0.1140643, 0.136595, 0.1591256, 0.1816562, 0.2041869, 
    0.2267175, 0.2492481, 0.2843918, 0.2747316, 0.2650714, 0.2554112, 
    0.245751, 0.2360907, 0.2264305, 0.1777242, 0.1663211, 0.1549179, 
    0.1435147, 0.1321116, 0.1207084, 0.1093052, 0.114393,
  0.3080943, 0.2932978, 0.1543645, 0.001124181, 0.04341831, 0.1019519, 
    0.07164619, 0.002705211, 0.03243441, 0.1350578, 0.2695448, 0.337139, 
    0.3188917, -0.00712925, 0.03568517, 0.04203487, 0.07082275, 0.07049537, 
    0.03582789, 0.09003742, 0.6219528, 0.7216404, 0.5773456, 0.2656536, 
    0.3061293, 0.2293136, 0.2262159, 0.2716772, 0.3287408,
  0.2326753, 0.06125122, 0.04385129, 0.004138701, 0.1389631, 0.2107148, 
    0.02810327, 0.3143154, 0.3080222, 0.277417, 0.2305294, 0.1778313, 
    0.05998614, 0.137907, 0.2623836, 0.2970552, 0.3631673, 0.3940248, 
    0.4269267, 0.3810286, 0.4343266, 0.3658237, 0.4169137, 0.5922614, 
    0.2965612, 0.3033271, 0.4510951, 0.538571, 0.4448643,
  0.562488, 0.5195694, 0.5709913, 0.4762004, 0.4102906, 0.4547261, 0.3335533, 
    0.3696454, 0.3815234, 0.2923739, 0.1918074, 0.2230927, 0.3220595, 
    0.3279318, 0.2933405, 0.342169, 0.4081841, 0.4406582, 0.3989094, 
    0.2740872, 0.2206354, 0.2126671, 0.2284484, 0.2784724, 0.3258277, 
    0.3640658, 0.4012429, 0.4202048, 0.5621699,
  0.4377044, 0.4234122, 0.4273262, 0.399064, 0.4077209, 0.3805239, 0.3371517, 
    0.2778595, 0.2985123, 0.3476612, 0.2637172, 0.2636266, 0.2348404, 
    0.2108476, 0.2040302, 0.3239743, 0.3639798, 0.4329394, 0.4274229, 
    0.3761131, 0.3013668, 0.2633023, 0.2375038, 0.1704258, 0.05065888, 
    0.292152, 0.5582676, 0.3776114, 0.4946643,
  0.2165756, 0.1738354, 0.1116802, 0.194142, 0.1805999, 0.1808068, 0.2501986, 
    0.3220208, 0.3092129, 0.1688524, 0.07548571, 0.05136415, 0.08564716, 
    0.1885184, 0.2400392, 0.3035634, 0.3590554, 0.3276343, 0.2349963, 
    0.1501407, 0.1347428, 0.1413356, 0.1831287, 0.155864, 0.01908629, 
    0.1354625, 0.1663901, 0.1672841, 0.1966804,
  0.1508268, 0.05061591, 0.01482225, 0.1023963, 0.1591447, 0.1508449, 
    0.1736183, 0.2552794, 0.1910956, 0.01669024, 0.01153699, -9.594645e-06, 
    0.01057638, 0.06042734, 0.1879618, 0.1211428, 0.1441608, 0.09946191, 
    0.3136958, 0.2007879, 0.1046235, 0.04327082, 0.06346829, 0.007919575, 
    0.04826582, 0.1416074, 0.1407345, 0.05957411, 0.162642,
  0.3508915, -0.0004651336, 1.143535e-05, 0.06560939, 0.07198826, 
    0.006707974, 0.02200981, 0.04764527, 0.07388934, 0.03043717, 
    1.302828e-06, -1.709537e-08, 0.08367443, 0.09720309, 0.05336328, 
    0.05081734, 0.07288998, 0.1145726, 0.05545889, 0.01825004, 0.01893792, 
    0.07526831, 0.3575978, 0.02986567, 0.09119501, 0.07353482, 0.1071057, 
    0.07502714, 0.2067783,
  0.5104324, 0.09145913, 0.001688363, 0.03265525, 0.03129009, 0.04126491, 
    0.0359746, 0.05945909, 0.04618587, 0.1661259, 0.02338858, 0.02875016, 
    0.1156441, 0.1003649, 0.04940008, 0.04754257, 0.027622, 0.04058792, 
    0.01896136, 0.01559583, 0.0437578, 0.2530604, 0.4776749, 0.02714035, 
    0.002384231, 0.0002787818, 0.03756977, 0.1479873, 0.447992,
  0.2754237, 0.1700495, 0.0173908, 0.0294875, 0.2044861, 0.07493553, 
    0.02904681, 0.05080556, 0.05570236, 0.08192036, 0.02876948, 0.1387058, 
    0.02463091, 0.02075882, 0.01131583, 0.01491223, 0.01966952, 0.01706339, 
    0.02237652, 0.04833464, 0.2274957, 0.4130366, 0.1440198, 0.01216703, 
    0.0006744454, 0.03768278, 0.0319711, 0.08262932, 0.4159417,
  5.146061e-05, 2.251525e-05, 3.507303e-05, -0.0002718845, 0.01586651, 
    0.03794713, 0.07135821, 0.040068, 0.06702517, 0.03478816, 0.02403431, 
    0.03130399, 0.04393631, 0.0605075, 0.03569893, 0.06024791, 0.05786611, 
    0.07210957, 0.1109873, 0.1425941, 0.112763, 0.05648404, 0.284957, 
    0.07177772, 0.03569153, 0.02638261, 0.0524161, 0.1296363, 9.477245e-05,
  3.025027e-07, 1.608428e-08, -1.874997e-08, 0.0002571176, 1.324126e-10, 
    0.006080223, 0.02755882, 0.0549468, 0.03092119, 0.0427893, 0.02183269, 
    0.04301835, 0.03875435, 0.03461984, 0.01547295, 0.0171256, 0.01907717, 
    0.0418616, 0.1133364, 0.1775754, 0.05066359, 0.2097735, 0.02154426, 
    0.019944, 0.02407905, 0.05923593, 0.0798972, 0.08438166, 1.088809e-07,
  2.091103e-07, 0.01198344, 0.0006632438, 0.0001166942, -0.0002102805, 
    8.795662e-09, -0.0003616473, 0.05340595, 0.2872573, -0.000104943, 
    0.1018437, 0.07091138, 0.1726698, 0.09283223, 0.06367151, 0.1054746, 
    0.04878986, 0.09489347, 0.1841046, 0.02165946, 0.002949686, 0.03631696, 
    0.03896243, 0.03955747, 0.02408101, 0.0334012, 0.05607449, 0.07340587, 
    -0.0003671054,
  0.02847517, 0.008896211, 0.08591042, 0.2483511, 0.025284, 0.00443521, 
    0.0489182, 0.0006008961, 0.01763293, 0.01443029, 0.1472373, 0.09923008, 
    0.1928208, 0.2985914, 0.2343871, 0.2684851, 0.2794683, 0.4108498, 
    0.2715751, 0.01586529, 0.01499823, 0.06840079, 0.1899363, 0.0800502, 
    0.09410021, 0.1056065, 0.1638266, 0.1262344, 0.01808324,
  0.2644203, 0.3933437, 0.3399713, 0.2752475, 0.1624442, 0.09675723, 
    0.1102806, 0.2544411, 0.1262736, 0.09349356, 0.08360583, 0.4170176, 
    0.306437, 0.2555893, 0.2766187, 0.3227917, 0.2220099, 0.3052178, 
    0.2781976, 0.2151409, 0.147016, 0.1577274, 0.3028021, 0.3428384, 
    0.2365331, 0.3287204, 0.374111, 0.39821, 0.3853235,
  0.1912457, 0.2174434, 0.3281024, 0.5423563, 0.4410825, 0.2070205, 
    0.3245212, 0.2626897, 0.4049918, 0.3830505, 0.3692445, 0.4863337, 
    0.3566101, 0.3773412, 0.3238228, 0.2111769, 0.5241752, 0.4722181, 
    0.3654781, 0.09072305, 0.3025478, 0.3614537, 0.2126094, 0.4720972, 
    0.4390458, 0.3234089, 0.2864933, 0.3167028, 0.2993149,
  0.1738475, 0.09119841, 0.237972, 0.2510548, 0.37077, 0.4178941, 0.5732868, 
    0.496813, 0.3062126, 0.3858268, 0.4675612, 0.4479536, 0.3963783, 
    0.3458986, 0.2568605, 0.5163381, 0.3836488, 0.3659983, 0.5248946, 
    0.4443497, 0.4130184, 0.5065883, 0.2655039, 0.4759215, 0.2329128, 
    0.643796, 0.3055898, 0.2134266, 0.2397902,
  0.3750318, 0.377361, 0.3854253, 0.3310969, 0.4249927, 0.464702, 0.4362527, 
    0.4548194, 0.2644966, 0.5675048, 0.5217511, 0.4383935, 0.4009377, 
    0.3366205, 0.3790792, 0.3465992, 0.3468017, 0.3691313, 0.358487, 
    0.418691, 0.4179776, 0.3205805, 0.2680426, 0.2872647, 0.2228859, 
    0.199835, 0.2688222, 0.3243402, 0.354651,
  0.09338196, 0.09071989, 0.08805783, 0.08539577, 0.08273371, 0.08007164, 
    0.07740957, 0.06431968, 0.08602139, 0.1077231, 0.1294248, 0.1511265, 
    0.1728282, 0.1945299, 0.2383488, 0.2274456, 0.2165424, 0.2056392, 
    0.1947359, 0.1838327, 0.1729295, 0.146331, 0.1381945, 0.1300581, 
    0.1219217, 0.1137853, 0.1056489, 0.0975125, 0.09551162,
  0.3187168, 0.2886704, 0.1422607, -0.0007444991, 0.04289641, 0.107171, 
    0.07639468, 0.01642817, 0.03561177, 0.059902, 0.2358191, 0.3806417, 
    0.3750287, -0.01507832, 0.06471682, 0.07433524, 0.135124, 0.06717192, 
    0.03235918, 0.1208467, 0.5802772, 0.7089478, 0.5706217, 0.2689874, 
    0.2593323, 0.2533021, 0.2343808, 0.2568457, 0.349263,
  0.2289545, 0.04816006, 0.03125549, -0.0005300305, 0.08910819, 0.1817485, 
    0.009474302, 0.2496246, 0.2756616, 0.2255481, 0.1907623, 0.1804764, 
    0.02321101, 0.1114417, 0.2802739, 0.3199671, 0.4053659, 0.4195276, 
    0.4426819, 0.45582, 0.4416326, 0.3760503, 0.4227954, 0.5727921, 
    0.3075578, 0.3859167, 0.5337607, 0.5498825, 0.4439977,
  0.6008882, 0.5799072, 0.5572793, 0.4198255, 0.3476262, 0.3829026, 
    0.2833858, 0.3003508, 0.3381702, 0.2472121, 0.1516523, 0.2027014, 
    0.2949636, 0.3060602, 0.2672136, 0.312335, 0.3916021, 0.4399329, 
    0.352999, 0.2424459, 0.1948121, 0.178941, 0.1988179, 0.2489724, 
    0.2666168, 0.4137357, 0.4066851, 0.4521811, 0.5453027,
  0.3904518, 0.3777761, 0.342927, 0.3715993, 0.3583489, 0.3244181, 0.2864883, 
    0.2397541, 0.2784344, 0.3126077, 0.2378168, 0.2664065, 0.2006067, 
    0.1726432, 0.166691, 0.3228601, 0.4064053, 0.3575228, 0.3885749, 
    0.3563365, 0.2623613, 0.22906, 0.2033318, 0.1460753, 0.04574489, 
    0.2521782, 0.5663174, 0.3341842, 0.3990743,
  0.187045, 0.1570517, 0.1146229, 0.1678167, 0.165585, 0.2074136, 0.272108, 
    0.3150556, 0.2762958, 0.1581879, 0.03513802, 0.02877506, 0.06479447, 
    0.2662342, 0.2380465, 0.2874594, 0.2868263, 0.2873578, 0.1812544, 
    0.1165639, 0.110893, 0.08614025, 0.1333714, 0.1369566, 0.01291229, 
    0.1272372, 0.1069576, 0.1207158, 0.1650647,
  0.06473687, 0.1096151, 0.01493166, 0.08147658, 0.1325879, 0.09020781, 
    0.09045848, 0.08220568, 0.08520163, 0.006484775, 0.006541765, 
    -8.20663e-05, 0.007694693, 0.02775344, 0.1419688, 0.07613602, 0.1014588, 
    0.04487628, 0.2571939, 0.1773661, 0.03991036, 0.01459702, 0.02288219, 
    0.01759847, 0.04432035, 0.1262978, 0.1412369, 0.04180983, 0.106796,
  0.1933278, 0.003813213, -7.445261e-05, 0.0307394, 0.008356315, 
    0.0002426372, 0.00481006, 0.01676779, 0.02689083, 0.01008619, 
    4.942139e-08, 4.872126e-08, 0.03375852, 0.06725425, 0.02605024, 
    0.04415549, 0.04319053, 0.04920764, 0.02339738, 0.006490031, 0.002705575, 
    0.02271754, 0.1357621, 0.01945425, 0.06973492, 0.07424962, 0.05077317, 
    0.01239192, 0.05867194,
  0.4654574, 0.1763665, 0.0005775173, 0.08310664, 0.01472287, 0.01576508, 
    0.01280249, 0.03983717, 0.01293193, 0.03344967, 0.008791142, 0.01682936, 
    0.09588124, 0.02107911, 0.01446742, 0.02682789, 0.005862036, 0.005761788, 
    0.003815882, 0.002268493, 0.009045929, 0.07881732, 0.458903, 0.03162068, 
    0.0009140254, 8.919622e-05, 0.004715709, 0.04661418, 0.1764362,
  0.1955163, 0.1412056, 0.01725105, 0.03045273, 0.05540633, 0.03810174, 
    0.01538439, 0.01724749, 0.05776571, 0.04309305, 0.004738788, 0.0187143, 
    0.003960575, 0.002635589, 0.001363995, 0.002604979, 0.004112761, 
    0.01076491, 0.01028075, 0.02708603, 0.1181332, 0.4240336, 0.4889812, 
    0.007725241, 0.0003091958, 0.007736998, 0.005545493, 0.03930445, 0.223545,
  2.977776e-05, 2.599016e-05, 2.102162e-05, 1.891844e-05, 0.02325954, 
    0.006536827, 0.0389169, 0.01471708, 0.03369722, 0.007592909, 0.0122733, 
    0.01175329, 0.02517554, 0.0330844, 0.01764421, 0.03542096, 0.04463066, 
    0.05313521, 0.07802369, 0.05378233, 0.04694263, 0.02265487, 0.310264, 
    0.05932463, 0.007572867, 0.01144933, 0.01020248, 0.05747202, 3.519976e-05,
  2.580744e-07, 1.262193e-08, -1.611279e-08, 7.695372e-06, 1.318837e-10, 
    0.05438704, 0.0224314, 0.01876443, 0.02623457, 0.01540595, 0.01160257, 
    0.01989007, 0.01531569, 0.01760653, 0.003854286, 0.00329355, 0.004094169, 
    0.01887569, 0.03576246, 0.07202426, 0.02003777, 0.1658607, 0.003889855, 
    0.0009800576, 0.004454559, 0.01357068, 0.01947709, 0.07939699, 
    1.053592e-07,
  1.545262e-07, 0.008855902, 0.0001887223, 0.0007034257, 0.0001928867, 
    6.842531e-09, -0.0002819454, 0.04676973, 0.2610387, -0.0001071588, 
    0.08006518, 0.04391747, 0.1143173, 0.05339406, 0.03696565, 0.05389685, 
    0.01156929, 0.03677031, 0.08239038, 0.01820946, 0.002456632, 0.03523995, 
    0.03041003, 0.01204259, 0.008476366, 0.01125244, 0.02763085, 0.02762375, 
    -0.0007499395,
  0.02589393, 0.006104154, 0.05729711, 0.2519625, 0.007628831, 0.002813052, 
    0.0445268, 0.0008337297, 0.01437973, 0.0137626, 0.1508203, 0.08241996, 
    0.1707659, 0.248386, 0.1953778, 0.2417576, 0.33072, 0.3807185, 0.2290142, 
    0.01616418, 0.01273407, 0.07075936, 0.1658877, 0.07193274, 0.0693645, 
    0.08539192, 0.1754479, 0.1588585, 0.01261705,
  0.1635164, 0.3986903, 0.3226238, 0.2529191, 0.1398797, 0.08937816, 
    0.08561602, 0.2595424, 0.121588, 0.1026153, 0.07203066, 0.3862493, 
    0.2217729, 0.2116506, 0.2160283, 0.2524668, 0.1810748, 0.3057584, 
    0.2755144, 0.2377184, 0.1338468, 0.1275358, 0.2646111, 0.3386283, 
    0.2046463, 0.2948721, 0.3013169, 0.3832863, 0.2970476,
  0.1476493, 0.2456495, 0.3094761, 0.5506433, 0.4570368, 0.2157482, 
    0.3326217, 0.247548, 0.3798018, 0.3328359, 0.3930694, 0.4784118, 
    0.3402825, 0.3054261, 0.2319341, 0.1570433, 0.5970244, 0.4409909, 
    0.4328733, 0.123106, 0.3001256, 0.3465571, 0.1820219, 0.37496, 0.3588887, 
    0.2822083, 0.2460714, 0.2512324, 0.2192848,
  0.1367829, 0.0690162, 0.2181653, 0.1832513, 0.3156935, 0.3731948, 
    0.6667923, 0.5094729, 0.2639143, 0.259585, 0.4762491, 0.4563533, 
    0.4265186, 0.4180823, 0.2855038, 0.4524801, 0.4164205, 0.3826949, 
    0.5340681, 0.3481306, 0.4270333, 0.6126787, 0.439627, 0.5297961, 
    0.1794107, 0.628203, 0.3037798, 0.1726273, 0.1782372,
  0.3251563, 0.4396713, 0.4496278, 0.3407545, 0.4245855, 0.4853863, 0.417852, 
    0.4498578, 0.3414164, 0.5652834, 0.5461918, 0.5046849, 0.4972459, 
    0.4210435, 0.4772235, 0.4327649, 0.3771068, 0.4190868, 0.4641101, 
    0.5201852, 0.4912809, 0.2935736, 0.2839576, 0.3505313, 0.199268, 
    0.1975775, 0.2923255, 0.3388992, 0.3981402,
  0.05107618, 0.04976555, 0.04845492, 0.04714429, 0.04583367, 0.04452304, 
    0.04321241, 0.03557192, 0.05345465, 0.07133737, 0.0892201, 0.1071028, 
    0.1249856, 0.1428683, 0.1710559, 0.1631553, 0.1552548, 0.1473543, 
    0.1394538, 0.1315533, 0.1236528, 0.1187856, 0.110114, 0.1014424, 
    0.09277084, 0.08409926, 0.07542767, 0.06675608, 0.05212468,
  0.3126582, 0.2743697, 0.09098388, 0.0002195216, 0.0270917, 0.08218889, 
    0.03692235, 0.02025953, 0.02625014, 0.01903494, 0.1317505, 0.3219119, 
    0.420167, -0.0141301, 0.08152571, 0.1437405, 0.2591218, 0.1131801, 
    0.03733232, 0.1179553, 0.5361602, 0.7094759, 0.4911294, 0.2605903, 
    0.2387604, 0.2914798, 0.2207943, 0.2387469, 0.3508524,
  0.2276814, 0.03937365, 0.02724021, 0.0001678167, 0.04595086, 0.1455964, 
    0.00150257, 0.1763527, 0.2399702, 0.1699218, 0.1428766, 0.1964539, 
    0.01269431, 0.09826992, 0.3052064, 0.3732514, 0.4868752, 0.4356474, 
    0.4255233, 0.4977305, 0.4132169, 0.3435282, 0.3432639, 0.5108615, 
    0.2971654, 0.4421369, 0.5677218, 0.5189943, 0.4416913,
  0.5494302, 0.5185256, 0.5294983, 0.3534955, 0.2798797, 0.3005768, 
    0.2515011, 0.2351353, 0.2550364, 0.1931163, 0.118267, 0.1728315, 
    0.2559151, 0.2751672, 0.2270508, 0.275212, 0.3359371, 0.3641642, 
    0.292476, 0.2026449, 0.1637415, 0.1475372, 0.1689072, 0.2195512, 
    0.2152219, 0.4451921, 0.413521, 0.4720172, 0.4651639,
  0.3510231, 0.3328008, 0.2737598, 0.3448471, 0.3237376, 0.2646513, 
    0.2360987, 0.1925989, 0.2517995, 0.2670433, 0.1974687, 0.2424217, 
    0.1498246, 0.1294023, 0.1351191, 0.3042761, 0.3552279, 0.2921321, 
    0.3218794, 0.3101577, 0.2181256, 0.1798919, 0.1717138, 0.1155088, 
    0.04621084, 0.2481316, 0.5272442, 0.275173, 0.3494864,
  0.1646304, 0.1200984, 0.09690008, 0.1577641, 0.1261557, 0.1742193, 
    0.2125266, 0.2717275, 0.2276368, 0.1130931, 0.01902508, 0.01617908, 
    0.04896145, 0.1803396, 0.2014048, 0.2682931, 0.2199073, 0.2161648, 
    0.1697788, 0.08883867, 0.07977268, 0.04900995, 0.08939146, 0.1180877, 
    0.02026544, 0.110039, 0.06777162, 0.08866722, 0.1383196,
  0.02929517, 0.0428727, 0.00985116, 0.05992025, 0.1050195, 0.0411994, 
    0.04297413, 0.03351851, 0.03887758, 0.003190285, 0.004336068, 
    -0.0002601331, 0.007850519, 0.01746863, 0.09266253, 0.03710995, 
    0.08411013, 0.02850229, 0.1932604, 0.1487848, 0.02100556, 0.005019303, 
    0.009265821, 0.01314381, 0.03379664, 0.086147, 0.1300355, 0.02930374, 
    0.07210726,
  0.08137705, 0.008471222, -5.824822e-05, 0.006412382, 0.0005852965, 
    4.522125e-05, 0.001193555, 0.006918148, 0.01218906, 0.005099745, 
    6.376075e-08, 2.861219e-08, 0.01040467, 0.03179952, 0.01011006, 
    0.03208094, 0.02346305, 0.01692146, 0.01280478, 0.00227509, 0.0006524332, 
    0.009136897, 0.05727942, 0.03104622, 0.04332363, 0.06284536, 0.02517306, 
    0.004661942, 0.02035721,
  0.1849156, 0.05616174, 0.0003213401, 0.1336862, 0.004284808, 0.004941241, 
    0.0026033, 0.02096082, 0.002691861, 0.009474825, 0.004221548, 
    0.002104368, 0.05443752, 0.003767892, 0.00166214, 0.010012, 0.001589168, 
    0.001013891, 0.00176685, 0.0008879109, 0.002715275, 0.02610886, 
    0.2060518, 0.03280807, 0.0005016181, 5.692275e-05, 0.00141139, 
    0.01707196, 0.06849131,
  0.05624056, 0.1401252, 0.01386306, 0.02456129, 0.01244304, 0.02100507, 
    0.009010407, 0.002515166, 0.06098307, 0.02907979, 0.001748463, 
    0.00543705, 0.000921764, 0.0003284464, 0.0004342965, 0.0009856328, 
    0.0005186269, 0.001490033, 0.0008587856, 0.003997395, 0.04307477, 
    0.1937283, 0.3172081, 0.006542974, 0.0002170017, 0.001790483, 
    0.000790661, 0.005848489, 0.06950407,
  2.497832e-05, 1.892038e-05, 9.715644e-06, 0.0003677577, 0.04341925, 
    0.001993122, 0.01943827, 0.007652137, 0.01905789, 0.0008267552, 
    0.008017171, 0.005323386, 0.01260351, 0.02105791, 0.006119431, 
    0.009135919, 0.02549444, 0.0281009, 0.02916588, 0.01392969, 0.02714639, 
    0.005219004, 0.2858795, 0.04478578, 0.002598544, 0.005445975, 
    0.002749486, 0.008691497, 1.476227e-05,
  2.294226e-07, 8.926808e-09, -1.194046e-08, 1.992186e-05, 1.002179e-10, 
    0.0235181, 0.02225204, 0.005081235, 0.01821796, 0.006326815, 0.005651071, 
    0.007313051, 0.005596214, 0.007428156, 0.0005199102, 0.0006398743, 
    0.001198216, 0.009512754, 0.01212962, 0.0321587, 0.01006121, 0.1245919, 
    0.001436022, -0.0003752375, 0.0009104564, 0.004525501, 0.007335198, 
    0.02736836, 1.025463e-07,
  1.370611e-07, 0.004604532, 6.035516e-05, 0.0004838335, 5.563406e-05, 
    6.14442e-09, -0.0002462735, 0.04514221, 0.2355035, -0.0001112188, 
    0.06644409, 0.01901558, 0.06380063, 0.02391233, 0.03008315, 0.01835919, 
    0.004232899, 0.01604041, 0.05032815, 0.005323722, 0.001603863, 0.0287724, 
    0.02944567, 0.003284015, 0.003474033, 0.003963079, 0.01201814, 0.0109426, 
    1.962958e-05,
  0.02297556, 0.001496147, 0.03302442, 0.2496865, 0.001873466, 0.001180826, 
    0.03625954, 0.0009691452, 0.01588189, 0.01266274, 0.134907, 0.05813835, 
    0.1323335, 0.2030383, 0.1578424, 0.2161743, 0.3344817, 0.2971972, 
    0.174085, 0.0117126, 0.01085231, 0.06275013, 0.1414874, 0.06433203, 
    0.04188043, 0.06734265, 0.141686, 0.1313109, 0.005396893,
  0.09209804, 0.3576047, 0.2725696, 0.2368331, 0.1032821, 0.1004717, 
    0.05583493, 0.235759, 0.09989942, 0.08776574, 0.0606938, 0.3447672, 
    0.1767984, 0.1660845, 0.1713359, 0.1879762, 0.1704059, 0.2935583, 
    0.2454762, 0.2530396, 0.1259754, 0.1013109, 0.2291349, 0.3289305, 
    0.1766273, 0.2739939, 0.2739344, 0.3223006, 0.2141518,
  0.1297237, 0.2451113, 0.2872978, 0.5226452, 0.4651877, 0.2354192, 
    0.3010395, 0.2158591, 0.346946, 0.3184075, 0.3378397, 0.4584658, 
    0.3036179, 0.2601881, 0.1729933, 0.1245739, 0.6008868, 0.3886682, 
    0.4872186, 0.1324167, 0.3015349, 0.3415263, 0.1563319, 0.3138888, 
    0.3004892, 0.2362187, 0.2286083, 0.2162738, 0.1776423,
  0.1047357, 0.04889, 0.2071916, 0.1289489, 0.2615004, 0.3142368, 0.6861098, 
    0.5040672, 0.2117413, 0.1980916, 0.4311889, 0.4232351, 0.4212993, 
    0.3762996, 0.3841012, 0.3835938, 0.4368877, 0.4172218, 0.5103418, 
    0.2640722, 0.4315473, 0.6258748, 0.509249, 0.5711117, 0.1256494, 
    0.6149898, 0.3130469, 0.1297102, 0.1403857,
  0.399143, 0.3972571, 0.5399946, 0.3684922, 0.4663485, 0.4877909, 0.4906499, 
    0.4857101, 0.4127479, 0.5635521, 0.5182444, 0.5542998, 0.5428053, 
    0.4420243, 0.5275494, 0.5068488, 0.4481654, 0.4942122, 0.5216148, 
    0.5926877, 0.5504225, 0.2517241, 0.3067074, 0.4441093, 0.2051913, 
    0.2068348, 0.2982432, 0.3837582, 0.4299474,
  0.02197386, 0.01974013, 0.01750641, 0.01527268, 0.01303895, 0.01080522, 
    0.008571495, 0.0065023, 0.01411693, 0.02173157, 0.0293462, 0.03696083, 
    0.04457546, 0.0521901, 0.0476786, 0.04893797, 0.05019734, 0.05145671, 
    0.05271608, 0.05397544, 0.05523481, 0.07519098, 0.0685507, 0.06191042, 
    0.05527015, 0.04862988, 0.04198961, 0.03534933, 0.02376084,
  0.2898149, 0.2412924, 0.04960679, 0.001169458, 0.004012011, 0.05783533, 
    0.02330606, 0.01200943, 0.00780157, 0.003758901, 0.0504301, 0.232202, 
    0.3929246, -0.008112356, 0.1325637, 0.2859482, 0.3592539, 0.2149498, 
    0.04563717, 0.1062891, 0.4608218, 0.6681904, 0.3898919, 0.2264913, 
    0.2086017, 0.2872649, 0.1878048, 0.2210472, 0.3330356,
  0.2203482, 0.03436279, 0.02806342, 0.000367783, 0.02307894, 0.1159288, 
    0.0002507779, 0.1259925, 0.1610393, 0.1207891, 0.09409433, 0.1813223, 
    0.006165835, 0.07248565, 0.3063363, 0.3610024, 0.4767734, 0.4291933, 
    0.38135, 0.4748833, 0.3274012, 0.2857797, 0.2694346, 0.4386896, 
    0.2447921, 0.4540371, 0.5151215, 0.4558858, 0.4233141,
  0.4538279, 0.413502, 0.4484487, 0.2751611, 0.2058182, 0.2315796, 0.2326705, 
    0.1796432, 0.1821301, 0.1448504, 0.08651732, 0.1309609, 0.2096965, 
    0.2223075, 0.1719939, 0.2161835, 0.2751851, 0.2796843, 0.228396, 
    0.1637141, 0.1292633, 0.1272817, 0.1381342, 0.1702177, 0.2038425, 
    0.4378106, 0.3925372, 0.4224738, 0.3833113,
  0.3121633, 0.2847663, 0.2230201, 0.298547, 0.2813671, 0.2097052, 0.1730378, 
    0.1542825, 0.1996668, 0.2107798, 0.1403997, 0.1762419, 0.08808973, 
    0.0873559, 0.1052259, 0.2353147, 0.2642153, 0.2229392, 0.2363225, 
    0.2165892, 0.1680489, 0.1259208, 0.120493, 0.08816708, 0.04471034, 
    0.2243162, 0.4474338, 0.24878, 0.3215577,
  0.1402926, 0.07214128, 0.0784818, 0.1384953, 0.09374958, 0.1223093, 
    0.1341973, 0.2079715, 0.1627983, 0.0691907, 0.01476915, 0.009658935, 
    0.03548082, 0.1221988, 0.1649162, 0.2095622, 0.1674756, 0.1838861, 
    0.1522705, 0.06773799, 0.051043, 0.02989168, 0.05532263, 0.09865563, 
    0.02102304, 0.08823677, 0.04630266, 0.06669137, 0.1009655,
  0.01494419, 0.02323397, 0.007014661, 0.03710739, 0.06038875, 0.02249134, 
    0.01899014, 0.01904835, 0.02285115, 0.001977207, 0.00238094, 
    -0.0003415685, 0.003368202, 0.01020046, 0.06222466, 0.02210086, 
    0.05804193, 0.02137631, 0.1375023, 0.1052841, 0.00929956, 0.00299015, 
    0.005235252, 0.008713537, 0.02361527, 0.0557121, 0.09404641, 0.01857517, 
    0.04051207,
  0.04332291, 0.008976307, -2.959494e-05, 0.002666739, -0.0002874301, 
    1.901305e-05, 0.0005670834, 0.003634912, 0.007132197, 0.003179133, 
    5.998194e-08, 3.154382e-08, 0.005050154, 0.0113104, 0.002071332, 
    0.01055956, 0.01095026, 0.006643797, 0.01041629, 0.0003311978, 
    0.0002974599, 0.004856558, 0.02977316, 0.01252015, 0.02499333, 
    0.05262433, 0.01188057, 0.002536672, 0.01008912,
  0.09415611, 0.02450617, 0.0001537166, 0.12815, 0.000670352, 0.001229309, 
    0.0004461579, 0.0074617, 0.0009836684, 0.004465987, 0.001751332, 
    0.0006008952, 0.02908538, 0.001436055, 0.000620914, 0.005060578, 
    0.0005537001, 0.0004748873, 0.001068279, 0.0004928519, 0.001315765, 
    0.01251398, 0.1131193, 0.03349112, 0.0002902596, 2.847587e-05, 
    0.001002784, 0.008836855, 0.03379646,
  0.02476824, 0.1377153, 0.01306472, 0.01647749, 0.005636636, 0.009211536, 
    0.003318459, 0.0008375984, 0.04665506, 0.02432353, 0.0009719259, 
    0.002739759, 0.0004580754, 0.0001960164, 0.0001755353, 0.0005252769, 
    0.0002647103, 0.0002623018, 0.0002407775, 0.001021944, 0.0132513, 
    0.09022606, 0.1841759, 0.01007462, 0.0001169113, 0.0009060453, 
    7.247164e-05, 0.001958882, 0.03070939,
  8.455555e-07, 3.485985e-06, 6.540235e-06, 0.000162515, 0.03320139, 
    0.001118384, 0.006834997, 0.004567454, 0.008484219, 6.032827e-05, 
    0.004172034, 0.002569458, 0.004600095, 0.01170481, 0.001983169, 
    0.002367517, 0.01128417, 0.01466496, 0.01282181, 0.004940951, 0.02208832, 
    0.0006796038, 0.2235718, 0.03229412, 0.001231289, 0.001800131, 
    0.001118432, 0.003144643, 1.515494e-07,
  2.094179e-07, 7.519972e-09, -8.527661e-09, 1.661567e-05, 1.259818e-10, 
    0.01028092, 0.01473649, 0.002243495, 0.01329932, 0.002589371, 
    0.002887932, 0.002853237, 0.002377627, 0.003073994, 0.0002131836, 
    0.0002589902, 0.0005342014, 0.003177256, 0.004617203, 0.01829273, 
    0.005367524, 0.09850822, 0.0008107444, -0.0006366564, 0.0004235635, 
    0.002381491, 0.003965775, 0.01537841, 1.012974e-07,
  1.256592e-07, 0.004135725, 3.82392e-05, 0.0001034898, -9.924062e-05, 
    5.809786e-09, -0.0001772109, 0.0423155, 0.2091953, 0.0001923218, 
    0.04381328, 0.01039544, 0.035364, 0.009237499, 0.01260088, 0.00766211, 
    0.002073637, 0.007244422, 0.03580025, 0.002392577, 0.00172789, 
    0.02230157, 0.0219028, 0.001257788, 0.000703926, 0.001621891, 
    0.004966451, 0.005494207, 0.005302788,
  0.01723113, 0.000654558, 0.01799443, 0.2346818, 3.699669e-05, 0.0005971771, 
    0.02643494, 0.0008553958, 0.01134716, 0.01038003, 0.1236963, 0.04161717, 
    0.09273977, 0.1656441, 0.1237803, 0.1820034, 0.2620977, 0.2069169, 
    0.1160329, 0.008846731, 0.007684239, 0.04685116, 0.1189203, 0.05227152, 
    0.02013109, 0.03809821, 0.0949344, 0.09061421, 0.001073898,
  0.05499074, 0.2977253, 0.2114938, 0.1960036, 0.07974576, 0.08431202, 
    0.04203675, 0.1957634, 0.0792447, 0.0662695, 0.05306293, 0.2996973, 
    0.1404118, 0.1262463, 0.1278851, 0.1353411, 0.1641684, 0.2685516, 
    0.1958098, 0.2634217, 0.117632, 0.06773166, 0.1832468, 0.302528, 
    0.1376558, 0.2620424, 0.2596454, 0.2761424, 0.1605396,
  0.1124102, 0.2346231, 0.2521551, 0.4633204, 0.423338, 0.2220566, 0.2485581, 
    0.1642916, 0.2886676, 0.2795499, 0.2698607, 0.4277098, 0.2701201, 
    0.2451767, 0.1298981, 0.08492988, 0.5965456, 0.3337236, 0.4448359, 
    0.1077629, 0.2916428, 0.3231384, 0.122107, 0.2610847, 0.2569644, 
    0.1884362, 0.2164522, 0.1817996, 0.1460034,
  0.07912725, 0.03111082, 0.2131064, 0.08927791, 0.197931, 0.2403458, 
    0.6701924, 0.4464636, 0.1716306, 0.1603599, 0.3618818, 0.422925, 
    0.4342511, 0.3477258, 0.4030575, 0.3224589, 0.4234141, 0.4305197, 
    0.4101842, 0.2011808, 0.3891153, 0.5853611, 0.5219827, 0.5620282, 
    0.105089, 0.5362214, 0.365921, 0.1006148, 0.1096661,
  0.3967714, 0.3261477, 0.6111372, 0.4589721, 0.4435437, 0.4843043, 
    0.5621275, 0.5381909, 0.4976722, 0.6148762, 0.5719906, 0.6382038, 
    0.5911634, 0.4616576, 0.57522, 0.6012988, 0.5183623, 0.4962991, 
    0.5436729, 0.5353705, 0.5542439, 0.2563363, 0.3429752, 0.4907917, 
    0.1992763, 0.2238827, 0.273483, 0.3867991, 0.4301828,
  0.004051184, 0.003536265, 0.003021346, 0.002506427, 0.001991509, 
    0.00147659, 0.0009616712, 0.001004457, 0.003810836, 0.006617216, 
    0.009423596, 0.01222998, 0.01503635, 0.01784273, 0.0202607, 0.02199587, 
    0.02373103, 0.0254662, 0.02720136, 0.02893652, 0.03067169, 0.03722743, 
    0.03320081, 0.02917418, 0.02514756, 0.02112093, 0.01709431, 0.01306768, 
    0.004463119,
  0.2746014, 0.2083342, 0.01659939, 0.0005202598, 0.004654234, 0.0359421, 
    0.004763685, -9.145874e-05, 0.001463019, 0.003135997, 0.02228054, 
    0.111597, 0.288616, -0.005821587, 0.1771394, 0.4121339, 0.4044406, 
    0.2338977, 0.04260492, 0.1268824, 0.3748804, 0.6476714, 0.3080634, 
    0.1802965, 0.1801014, 0.3006893, 0.1673064, 0.1952564, 0.3093567,
  0.2182901, 0.03538722, 0.0288497, 0.0002420038, 0.01031203, 0.09140437, 
    -0.0001033551, 0.09768487, 0.09101739, 0.08598219, 0.08138752, 0.1451119, 
    0.00291166, 0.04689323, 0.2912062, 0.3499449, 0.4303305, 0.3767285, 
    0.329987, 0.4015269, 0.2485667, 0.2166982, 0.1914721, 0.3660864, 
    0.2159523, 0.4259869, 0.4327028, 0.3728714, 0.393819,
  0.3528851, 0.3279329, 0.3597886, 0.2083166, 0.1557321, 0.1750011, 0.188944, 
    0.1355894, 0.1322447, 0.1079607, 0.05990876, 0.09812852, 0.15723, 
    0.1751076, 0.1249874, 0.1637095, 0.2196755, 0.216506, 0.1785348, 
    0.1260114, 0.1002001, 0.09856432, 0.1002052, 0.1234211, 0.1727314, 
    0.3630088, 0.3188925, 0.3389618, 0.3023246,
  0.2641741, 0.2239043, 0.1868794, 0.2473934, 0.234934, 0.1604288, 0.1277584, 
    0.1220683, 0.1540539, 0.1547148, 0.0917377, 0.1162018, 0.04871492, 
    0.05389314, 0.07469238, 0.1529377, 0.1847716, 0.1436956, 0.1510586, 
    0.1463152, 0.1121157, 0.08241334, 0.07901341, 0.07053553, 0.03675564, 
    0.1657855, 0.3632273, 0.2071868, 0.2830581,
  0.1007592, 0.0446112, 0.05976751, 0.0947189, 0.05911468, 0.07850073, 
    0.08027612, 0.138572, 0.1012735, 0.04091842, 0.01508855, 0.006431868, 
    0.0243442, 0.08403629, 0.1336206, 0.1432486, 0.116168, 0.1393023, 
    0.1220554, 0.04632399, 0.03211493, 0.01924992, 0.03323748, 0.08530235, 
    0.01960175, 0.06376684, 0.0276919, 0.04611696, 0.06703176,
  0.00885377, 0.01522285, 0.004914716, 0.0167371, 0.02541487, 0.0106808, 
    0.01073255, 0.01299104, 0.01597102, 0.001397958, 0.001428247, 
    -0.0003635403, 0.003214649, 0.004866006, 0.04875319, 0.01338445, 
    0.03378265, 0.0111311, 0.08504914, 0.06939688, 0.00400943, 0.002236241, 
    0.00371393, 0.005700117, 0.01560988, 0.0360713, 0.06217203, 0.01026368, 
    0.0191617,
  0.02811444, 0.007491164, -1.735393e-05, 0.001587088, -0.0001687164, 
    1.124344e-05, 0.0003445609, 0.002290602, 0.004889461, 0.002289828, 
    5.635532e-08, 2.985498e-08, 0.003203794, 0.003673165, 0.0008524319, 
    0.004538835, 0.00421074, 0.003485427, 0.007192813, 6.429372e-05, 
    0.0001736908, 0.003086986, 0.01898157, 0.007596021, 0.01390505, 
    0.04102646, 0.005545296, 0.001517647, 0.006199533,
  0.05850318, 0.01235712, 8.711997e-05, 0.08974199, 0.0001461343, 
    0.0004573253, 0.000135656, 0.00298859, 0.0005862855, 0.003302344, 
    0.0004898124, 0.0003215442, 0.01495305, 0.0008843569, 0.0003211705, 
    0.001887653, 0.0002736806, 0.0003030402, 0.0007401428, 0.000322781, 
    0.0008174255, 0.007553784, 0.07321284, 0.02480455, 0.0001901259, 
    1.695568e-05, 0.0008083959, 0.005614739, 0.02074154,
  0.01498542, 0.116629, 0.01340517, 0.01168955, 0.003444876, 0.004258249, 
    0.001461759, 0.0005482964, 0.02960812, 0.0312413, 0.0006428258, 
    0.001685996, 0.000272062, 0.0001022825, 8.004467e-05, 0.0003357826, 
    0.0001676764, 0.0001525619, 0.0001238709, 0.0005544567, 0.006429911, 
    0.05236836, 0.1199207, 0.01454324, 6.08409e-05, 0.0005798468, 
    -5.242676e-06, 0.001059434, 0.01817061,
  -4.015819e-05, 3.250747e-07, 8.031137e-06, 0.0002215704, 0.01535752, 
    0.0007540442, 0.002849761, 0.002480272, 0.003901004, -1.874713e-05, 
    0.001617583, 0.0007806736, 0.001762528, 0.005720187, 0.0005664432, 
    0.0006493292, 0.004403429, 0.006744216, 0.006308225, 0.002358909, 
    0.01245477, 0.0001253849, 0.184149, 0.02851574, 0.0007339169, 
    0.0006982719, 0.0005612727, 0.001730437, -1.558615e-05,
  1.952072e-07, 6.965228e-09, -6.496343e-09, 1.493524e-05, 1.228767e-10, 
    0.006024655, 0.004844611, 0.001156805, 0.006522731, 0.001300065, 
    0.0008291684, 0.001308214, 0.001055589, 0.001072278, 0.0001405978, 
    0.000163693, 0.0003500141, 0.0006770623, 0.002218567, 0.01236635, 
    0.003622888, 0.07793231, 0.0005382208, -0.0005902609, 0.0002621554, 
    0.001515456, 0.002571396, 0.009737695, 1.010708e-07,
  1.203686e-07, 0.001862863, 3.301519e-05, -1.192303e-05, -7.695851e-05, 
    5.604243e-09, -0.0001340983, 0.04076668, 0.1837565, 0.0004911852, 
    0.01954561, 0.004634304, 0.01736376, 0.00366931, 0.004834957, 
    0.004446815, 0.001254716, 0.003681801, 0.02491967, 0.001445604, 
    0.0009804287, 0.02051863, 0.01557179, 0.0008282718, 0.0003347137, 
    0.0008914263, 0.002073402, 0.00348711, 0.004913833,
  0.0133385, 0.0002329344, 0.01085968, 0.2187708, -0.0003772852, 
    0.0003659248, 0.01807612, 0.0006889628, 0.006077408, 0.009053282, 
    0.1081164, 0.0281996, 0.06084298, 0.1294091, 0.08645909, 0.1330367, 
    0.185845, 0.1219174, 0.07021588, 0.007895244, 0.004847502, 0.03178023, 
    0.09180955, 0.03986857, 0.008151415, 0.01905006, 0.05620913, 0.05701607, 
    -0.0002802074,
  0.03765092, 0.2381033, 0.1567066, 0.141589, 0.05548451, 0.0666076, 
    0.03402579, 0.158932, 0.0622717, 0.05156614, 0.04536574, 0.2558407, 
    0.1075047, 0.08662685, 0.0907936, 0.08735808, 0.1269128, 0.206545, 
    0.1363225, 0.2572879, 0.09738117, 0.04551232, 0.1412514, 0.2695554, 
    0.1036041, 0.2497484, 0.2233381, 0.2234582, 0.1187768,
  0.07690454, 0.2241222, 0.2193717, 0.3980115, 0.3589264, 0.1927658, 
    0.2057346, 0.1317917, 0.2209403, 0.2144556, 0.2205527, 0.3711909, 
    0.2418774, 0.2073509, 0.09753326, 0.05236212, 0.5640966, 0.2841321, 
    0.3906871, 0.09123193, 0.260035, 0.2972786, 0.08922292, 0.2056445, 
    0.2132533, 0.1456795, 0.1712929, 0.1309025, 0.1013516,
  0.05820784, 0.01728012, 0.209457, 0.06484276, 0.1487983, 0.1841514, 
    0.5836433, 0.3871743, 0.154686, 0.1264475, 0.2873806, 0.3248049, 
    0.4279981, 0.2905897, 0.3545077, 0.2782855, 0.3558241, 0.3750288, 
    0.3288107, 0.1591569, 0.3326611, 0.5445181, 0.4939124, 0.5134207, 
    0.07839978, 0.4471641, 0.4518313, 0.07794034, 0.08408431,
  0.3733396, 0.2690133, 0.6237263, 0.4777766, 0.3955718, 0.4629947, 
    0.5213113, 0.4807036, 0.4772777, 0.5725589, 0.5486633, 0.5794213, 
    0.5690317, 0.4196434, 0.4690842, 0.571634, 0.4739441, 0.4697957, 
    0.4934394, 0.5215512, 0.508163, 0.2400512, 0.3822973, 0.5316184, 
    0.1895218, 0.2659409, 0.2607937, 0.3677644, 0.4370263,
  0.001986551, 0.001687597, 0.001388643, 0.001089688, 0.000790734, 
    0.0004917796, 0.0001928253, 0.001431668, 0.002866327, 0.004300985, 
    0.005735643, 0.007170301, 0.00860496, 0.01003962, 0.01342644, 0.01419735, 
    0.01496826, 0.01573917, 0.01651007, 0.01728098, 0.01805189, 0.01791029, 
    0.01600368, 0.01409707, 0.01219045, 0.01028384, 0.008377228, 0.006470616, 
    0.002225715,
  0.2511431, 0.09400836, 0.01772259, 0.0004134012, 0.002435744, 0.02235826, 
    0.002720215, -3.537614e-05, 6.594363e-05, 0.002974506, 0.01419324, 
    0.06084324, 0.159081, -0.004394894, 0.2354107, 0.412125, 0.4069834, 
    0.2279518, 0.04350082, 0.1670123, 0.3034405, 0.6224028, 0.2590379, 
    0.1481027, 0.1763749, 0.3133805, 0.1852323, 0.1703988, 0.2684582,
  0.2007191, 0.03620718, 0.03140713, 0.0005056514, 0.01153691, 0.07806088, 
    -0.0002460864, 0.07740083, 0.06134168, 0.06814684, 0.07269952, 0.1273589, 
    0.001854039, 0.02807408, 0.2710553, 0.3116941, 0.3655946, 0.3318883, 
    0.2884319, 0.3403027, 0.1848344, 0.1735192, 0.1543569, 0.3101572, 
    0.1980013, 0.3719288, 0.3595671, 0.3075468, 0.3635884,
  0.287265, 0.2632316, 0.2960149, 0.1660214, 0.121138, 0.1372369, 0.1595172, 
    0.1110418, 0.1058226, 0.0854671, 0.04722565, 0.07798388, 0.1243009, 
    0.1468747, 0.09944734, 0.1321769, 0.1865297, 0.182208, 0.1498033, 
    0.10225, 0.08359914, 0.0790459, 0.07649688, 0.09659027, 0.1464052, 
    0.2943633, 0.2685319, 0.2712066, 0.2517588,
  0.2246554, 0.1801761, 0.1632718, 0.2137807, 0.1995225, 0.1345575, 
    0.1041594, 0.09722611, 0.1210099, 0.1225217, 0.0667216, 0.0819506, 
    0.03100411, 0.03716474, 0.0497082, 0.1051255, 0.1381896, 0.09768578, 
    0.1069449, 0.1033002, 0.07599912, 0.05815022, 0.05682532, 0.05956644, 
    0.02596977, 0.1308024, 0.289939, 0.1747894, 0.2372869,
  0.06295331, 0.02714267, 0.04041355, 0.06492106, 0.03642493, 0.04752627, 
    0.05230568, 0.09605046, 0.06433841, 0.02876243, 0.013229, 0.005059999, 
    0.0156411, 0.05862467, 0.1091672, 0.1001287, 0.08001559, 0.1052801, 
    0.08573736, 0.03063004, 0.02143033, 0.01212615, 0.02351682, 0.07583682, 
    0.01944874, 0.04416775, 0.01716909, 0.03011889, 0.04418657,
  0.006446914, 0.01169515, 0.003367034, 0.009516364, 0.01320534, 0.005312135, 
    0.006529339, 0.009812449, 0.01240703, 0.001087866, 0.001032992, 
    -0.0003226972, 0.002867508, 0.003057973, 0.03126133, 0.007213458, 
    0.01789425, 0.007002707, 0.04611033, 0.04392217, 0.002477422, 
    0.001807442, 0.00288795, 0.004483549, 0.01101735, 0.02029845, 0.0367513, 
    0.005888321, 0.01055174,
  0.02086974, 0.004900001, -1.196058e-05, 0.001131081, 8.005465e-05, 
    7.979937e-06, 0.0002448542, 0.001659595, 0.003740596, 0.001808743, 
    5.428628e-08, 2.866383e-08, 0.002373867, 0.001826856, 0.0005609184, 
    0.002409878, 0.002053465, 0.002327114, 0.003919949, 3.787988e-05, 
    0.0001197132, 0.002247959, 0.01386427, 0.005474587, 0.008528162, 
    0.03382672, 0.002782248, 0.001041567, 0.004414305,
  0.04208074, 0.007560634, 0.0001159747, 0.06352809, 8.730721e-05, 
    0.0002804974, 7.90813e-05, 0.001347697, 0.0004115179, 0.002731656, 
    0.0002756811, 0.0002110148, 0.00720698, 0.0006314642, 0.0001736183, 
    0.0009465636, 0.0001735721, 0.0002261728, 0.0005679526, 0.0002394667, 
    0.0005910171, 0.005344988, 0.05431035, 0.01830897, 0.0005919687, 
    5.196608e-06, 0.0006419006, 0.004092687, 0.014798,
  0.01064268, 0.09430165, 0.01003262, 0.009127833, 0.002462521, 0.002226703, 
    0.0007962834, 0.0004154595, 0.02041783, 0.03831182, 0.0004792424, 
    0.001201145, 0.000183644, 5.990769e-05, 3.717097e-05, 0.0002438421, 
    0.0001241601, 0.0001081971, 8.188304e-05, 0.0003802168, 0.004171033, 
    0.03638181, 0.08867437, 0.006916325, 7.736935e-05, 0.0004220644, 
    3.102558e-05, 0.0007107883, 0.01267987,
  -0.0001671998, 2.52972e-08, 5.548631e-05, 0.0002737199, 0.007981341, 
    0.0005672906, 0.0006906739, 0.00116161, 0.001983166, -6.2975e-06, 
    0.0007914505, 0.0003603209, 0.0008272087, 0.002931248, 0.0002362339, 
    0.0003501564, 0.001927988, 0.002960705, 0.003172987, 0.001418224, 
    0.00649241, 0.0001117861, 0.1545455, 0.02923636, 0.0005158688, 
    0.0003871456, 0.0003598211, 0.00117128, -8.193353e-05,
  1.849536e-07, 6.64836e-09, -5.009605e-09, 1.412737e-05, -1.420787e-11, 
    0.004277098, 0.001694696, 0.0006407744, 0.003385172, 0.0007770566, 
    0.0003666706, 0.0006944404, 0.0006507122, 0.0004270944, 0.0001061603, 
    0.0001247888, 0.0002661383, 0.0003130167, 0.001551373, 0.00938751, 
    0.002770599, 0.06471919, 0.0004025726, -0.0007747322, 0.0001890751, 
    0.001101704, 0.001895286, 0.00707062, 1.015537e-07,
  1.178298e-07, 0.0007953221, 2.612565e-05, -2.154043e-05, -4.525657e-05, 
    5.45054e-09, -0.0001298093, 0.0501813, 0.1717471, 0.0007779077, 
    0.01171415, 0.002303159, 0.009624516, 0.00191457, 0.002715987, 
    0.003083517, 0.0009208276, 0.002211899, 0.01647853, 0.001025158, 
    0.0003924903, 0.02996599, 0.01543744, 0.0006267239, 0.0002525221, 
    0.000655162, 0.001194799, 0.00258604, 0.004399797,
  0.01204935, 2.353963e-06, 0.008300253, 0.2078764, -0.000422653, 
    0.0002665664, 0.01254276, 0.0005325651, 0.003889305, 0.007610807, 
    0.09844704, 0.01755418, 0.03938136, 0.1012938, 0.06223645, 0.09946585, 
    0.1259034, 0.07330538, 0.04198439, 0.007819123, 0.003840692, 0.02294026, 
    0.07041624, 0.02915474, 0.004820287, 0.01216691, 0.02938405, 0.03981493, 
    -0.0006781849,
  0.02758862, 0.1961196, 0.1215536, 0.1091078, 0.0429562, 0.05489954, 
    0.02809926, 0.1352363, 0.05211976, 0.04347987, 0.04258831, 0.2266413, 
    0.08493946, 0.05755867, 0.06919631, 0.05811378, 0.09169975, 0.1528063, 
    0.09305441, 0.2463257, 0.08087742, 0.03617507, 0.1125266, 0.2449844, 
    0.08002568, 0.2124151, 0.1798567, 0.1711208, 0.0893679,
  0.05037691, 0.2234854, 0.194254, 0.3434602, 0.3216031, 0.1736983, 
    0.1946714, 0.115936, 0.1911775, 0.179887, 0.1925182, 0.341758, 0.2234502, 
    0.1776085, 0.07685532, 0.03629753, 0.5338018, 0.2540345, 0.3645282, 
    0.08327582, 0.2395931, 0.2746532, 0.06715821, 0.1721996, 0.1755958, 
    0.1151516, 0.1244939, 0.09395616, 0.07205432,
  0.04250782, 0.01202203, 0.2220942, 0.05010959, 0.1198898, 0.1476021, 
    0.5254229, 0.3386096, 0.1551545, 0.1198005, 0.2405416, 0.2690791, 
    0.3643055, 0.2448954, 0.3044906, 0.2482502, 0.3140647, 0.3286498, 
    0.2696543, 0.1267918, 0.2846113, 0.4985094, 0.4354715, 0.4755161, 
    0.0615198, 0.3789133, 0.5562015, 0.06907083, 0.06638519,
  0.3639317, 0.2309282, 0.5100788, 0.4415416, 0.3432788, 0.3915924, 
    0.4136986, 0.3821922, 0.3897402, 0.4519497, 0.424199, 0.4346191, 
    0.4523625, 0.2957345, 0.3462496, 0.4343148, 0.365711, 0.3529118, 
    0.3661428, 0.3846584, 0.4173948, 0.2126903, 0.4076576, 0.5446542, 
    0.1977219, 0.2400873, 0.2714649, 0.3696538, 0.337609,
  0.001809807, 0.001398553, 0.0009873, 0.0005760467, 0.0001647934, 
    -0.0002464599, -0.0006577132, -0.003228507, -0.002229742, -0.001230976, 
    -0.0002322108, 0.0007665546, 0.00176532, 0.002764085, 0.00648501, 
    0.007537538, 0.008590065, 0.009642593, 0.01069512, 0.01174765, 
    0.01280017, 0.01356096, 0.01192092, 0.01028088, 0.008640844, 0.007000805, 
    0.005360765, 0.003720726, 0.002138809,
  0.2245727, 0.04111981, 0.01359705, 2.639707e-05, 0.001744294, 0.02036073, 
    0.002333286, -9.129529e-05, 6.75598e-05, 0.002257227, 0.01114273, 
    0.0588641, 0.1359673, -0.003294671, 0.3068175, 0.413423, 0.3996394, 
    0.2448706, 0.04540059, 0.192064, 0.2581198, 0.5879805, 0.2391487, 
    0.1355568, 0.1990618, 0.313818, 0.2166135, 0.1580038, 0.2355806,
  0.1996502, 0.05143648, 0.06061349, 0.001217458, 0.009398077, 0.07230517, 
    -0.0008073981, 0.07496605, 0.06414659, 0.06465667, 0.07273329, 0.126339, 
    0.007943328, 0.02971567, 0.2467388, 0.2832707, 0.3371407, 0.3070149, 
    0.2565765, 0.2980251, 0.1547693, 0.1555344, 0.1433297, 0.2834093, 
    0.1861398, 0.3442679, 0.3156087, 0.2717525, 0.3389685,
  0.2534989, 0.2284428, 0.2634032, 0.1461934, 0.1068956, 0.1210746, 
    0.1505774, 0.100616, 0.09284397, 0.07328101, 0.04167466, 0.06842716, 
    0.1108122, 0.1325067, 0.0880295, 0.1187978, 0.1615818, 0.1637637, 
    0.1325641, 0.08838108, 0.07508072, 0.06921399, 0.06295663, 0.08208016, 
    0.123952, 0.262274, 0.2568457, 0.2346795, 0.2241792,
  0.1915065, 0.1521854, 0.1388548, 0.17953, 0.1704445, 0.116935, 0.08915861, 
    0.08316385, 0.1041913, 0.1068977, 0.05476002, 0.06601381, 0.02367183, 
    0.0277522, 0.03799487, 0.0815255, 0.1073492, 0.07496083, 0.08558547, 
    0.08060417, 0.05695729, 0.04549132, 0.04487347, 0.06600796, 0.02156044, 
    0.1002482, 0.2337497, 0.1500943, 0.1951096,
  0.04587001, 0.01952202, 0.03078254, 0.04820818, 0.02467057, 0.03460986, 
    0.03850699, 0.06734471, 0.04465878, 0.02336489, 0.01078497, 0.004365752, 
    0.01151121, 0.04444433, 0.100697, 0.07638799, 0.05754476, 0.07524211, 
    0.05969044, 0.02406556, 0.01575314, 0.008198001, 0.01729931, 0.0740523, 
    0.01826601, 0.0289414, 0.0127319, 0.02228347, 0.03291292,
  0.005372829, 0.009588053, 0.004989857, 0.005990198, 0.008473559, 
    0.00368048, 0.004843725, 0.00819705, 0.01055586, 0.0009174935, 
    0.0007849363, -0.0002654175, 0.005010284, 0.001421306, 0.01709164, 
    0.004891997, 0.01063538, 0.005227059, 0.02831886, 0.02663267, 
    0.001809613, 0.001566542, 0.002474998, 0.003844163, 0.01291066, 
    0.01214131, 0.02128348, 0.003897781, 0.006885265,
  0.01734377, 0.003935551, -4.017749e-05, 0.0009195699, -7.678216e-05, 
    6.614683e-06, 0.0002049094, 0.001376879, 0.003173127, 0.001548139, 
    5.425043e-08, 2.763687e-08, 0.001976701, 0.001278541, 0.000448425, 
    0.001647128, 0.001391728, 0.00183893, 0.002159342, 2.859306e-05, 
    9.681422e-05, 0.001869632, 0.01147904, 0.004456861, 0.007668104, 
    0.05394028, 0.001843595, 0.0008400786, 0.003589579,
  0.03408339, 0.005309715, 0.00172051, 0.06205847, 6.601613e-05, 
    0.0002207547, 6.350762e-05, 0.0008537501, 0.0003342028, 0.001997035, 
    0.000208762, 0.0001673138, 0.004265271, 0.0005087102, 0.0001263127, 
    0.0006570155, 0.0001354356, 0.0001874677, 0.0004832913, 0.0001986819, 
    0.0004883664, 0.004360649, 0.0448125, 0.08253741, 0.005947402, 
    -1.568354e-05, 0.0005499291, 0.003372271, 0.01200058,
  0.008541656, 0.120227, 0.01033408, 0.008176392, 0.001983634, 0.001591522, 
    0.0005601014, 0.000273162, 0.03637862, 0.06390946, 0.0003983506, 
    0.0009861552, 0.0001454635, 4.519151e-05, 2.682486e-05, 0.0002001738, 
    0.0001036636, 8.890861e-05, 6.49125e-05, 0.0003058357, 0.003175614, 
    0.02842525, 0.07293667, 0.01187314, 0.003206009, 0.0003544537, 
    4.636747e-05, 0.000560333, 0.01009111,
  -0.0003778369, -5.2598e-05, 0.0005019726, 0.0003061602, 0.005494222, 
    0.0004696289, -0.0009110589, 0.0006620451, 0.0005735363, 3.593855e-06, 
    0.0005363188, 0.0002569778, 0.0005559734, 0.002025283, 0.0001533174, 
    0.0002579407, 0.001230216, 0.001734673, 0.001878237, 0.001113186, 
    0.003917199, 0.0001185054, 0.2339206, 0.03495217, 0.0004163036, 
    0.0002801081, 0.0002790047, 0.0008593516, -0.0007177857,
  1.781476e-07, 6.403926e-09, -3.481289e-09, 3.899401e-07, -3.159002e-10, 
    0.003417465, 0.004323268, 0.0004679297, 0.002462542, 0.0002409567, 
    0.0002456658, 0.0004685973, 0.0004944592, 0.0002730367, 9.007443e-05, 
    0.0001065177, 0.0002102685, 0.0002243398, 0.001249648, 0.007848518, 
    0.002325771, 0.05845244, 0.0003351183, -0.001346612, 0.0001543228, 
    0.0009072244, 0.00156192, 0.005762997, 1.042653e-07,
  1.17487e-07, 0.0005325195, 1.321608e-05, -1.06276e-05, -4.566056e-05, 
    5.460283e-09, -0.0002451981, 0.06962897, 0.1755748, 0.001084593, 
    0.008405144, 0.001601707, 0.006157587, 0.001283999, 0.002013447, 
    0.002506348, 0.0007573114, 0.001718091, 0.01191454, 0.000837722, 
    0.0002531651, 0.07191586, 0.02063855, 0.000526212, 0.0002173466, 
    0.0005421441, 0.0009201039, 0.002141563, 0.003464975,
  0.01666955, -0.0002083156, 0.006366328, 0.2045709, -0.0004727931, 
    0.0002205289, 0.009294837, 0.0004745311, 0.004052672, 0.006675228, 
    0.1099871, 0.01263718, 0.02753457, 0.07386822, 0.0461186, 0.06709543, 
    0.09059239, 0.05105107, 0.02782296, 0.007704804, 0.003963395, 0.02637739, 
    0.066342, 0.02159949, 0.003789225, 0.008885436, 0.01767652, 0.03058535, 
    -0.0009718133,
  0.02180574, 0.2040061, 0.1111903, 0.1070411, 0.0348108, 0.04726307, 
    0.02412112, 0.1307781, 0.0534362, 0.03868469, 0.05273194, 0.2368628, 
    0.06939183, 0.04200814, 0.05332802, 0.04344136, 0.07309872, 0.1154358, 
    0.06892936, 0.2525748, 0.07572529, 0.03177902, 0.1232081, 0.2564778, 
    0.07266602, 0.1739114, 0.1366103, 0.1324027, 0.06886186,
  0.03823762, 0.2507586, 0.2096361, 0.3412149, 0.3432402, 0.1919414, 
    0.2095025, 0.1313683, 0.1963017, 0.1944451, 0.199292, 0.3639503, 
    0.231256, 0.1998124, 0.06709766, 0.02947791, 0.5407681, 0.2462346, 
    0.4092284, 0.08598582, 0.2450422, 0.2724752, 0.05607663, 0.1688427, 
    0.1479174, 0.1010164, 0.09654147, 0.07376521, 0.05528603,
  0.03569981, 0.01001352, 0.2736686, 0.04105508, 0.1026445, 0.12411, 
    0.5087608, 0.3284029, 0.1890019, 0.1336501, 0.2507027, 0.2401779, 
    0.3187093, 0.2129846, 0.2811607, 0.2331166, 0.3000199, 0.3157699, 
    0.2388877, 0.1088392, 0.2587824, 0.4580208, 0.4040383, 0.4562759, 
    0.04629343, 0.3526334, 0.6136554, 0.06504256, 0.0559487,
  0.3497979, 0.2125242, 0.4673252, 0.3805221, 0.3064586, 0.3257843, 
    0.3308556, 0.3030222, 0.3176813, 0.3605712, 0.3267037, 0.3428708, 
    0.3633319, 0.2231982, 0.2702672, 0.3465581, 0.2863278, 0.2764228, 
    0.3240412, 0.3235088, 0.3536806, 0.2003309, 0.4159078, 0.5322804, 
    0.2200127, 0.2223815, 0.2916982, 0.3954227, 0.2738242,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -4.954702e-06, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0008251527, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, -6.271177e-06, 0, 0, 0, 0, 0, 0, 0, -0.0001175386, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.0003204219, 0, 0, 0,
  0, 0, -1.13965e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, -2.090035e-05, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.0007870967, -5.327915e-05, 0.001581971, 0, 
    -6.515444e-07, 0.0008662037, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3.672994e-05, -8.001684e-07, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0.0002111749, -3.77435e-05, 0, 0, 0, 0, 0, 0, 0, -0.0001988136, 
    -2.723663e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, -4.288225e-05, 0.002199712, 0, 
    0, 0,
  0, 0, -2.866954e-05, 0, 0, 0, 0, 0, 7.544798e-06, 0, 0, 0, 0, 
    -3.965341e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.099267e-05, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.00227801, -0.0001622717, 0.004560962, -4.510288e-05, 
    0.0001229582, 0.001591074, 0.0001286336, 0, 0, 0.0004814128, 0, 0, 
    -5.58423e-05, -8.245673e-05, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -5.092964e-05, -1.944676e-06, -2.131265e-05, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0.0006400415, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, -1.883469e-06, 0, 0, 0,
  0, 0, -1.950752e-05, 0, 0.0005310062, 5.442087e-05, 0.002631418, 
    -4.129605e-05, 0, 0, 0, 0, 0, -0.000189297, -7.137992e-05, -5.133168e-05, 
    0, 0, 0, 0, 0, 0, 0, -7.679454e-08, -9.140798e-05, 0.005686537, 0, 0, 0,
  0, 0, -2.855553e-05, 0, 0, 0.001212848, 0, 0, -6.008521e-05, -5.608389e-05, 
    0, 0, 0, 0.0001147859, 0, -1.223459e-06, 0, 0, 0, 0, 0, 0, 0, 
    -2.449136e-05, 0, 0, 6.919583e-05, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.006283578, -0.0003102303, 0.009508011, 0.002325651, 
    0.002024822, 0.003490037, 0.002482031, 0.0005214345, 0, 0.004725255, 
    0.0001885848, -3.821963e-05, -0.0001463529, 0.004895335, 0, 0, 0, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0003517914, -2.155753e-06, -5.904976e-05, 
    0.0009102497, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, -9.747487e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, -2.073661e-05, 0, 0, 0,
  0, 0, 0.003032253, 0, -1.42609e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, -8.351135e-05, 0, 0, 0,
  0, 0, -0.0001084161, 0, 0.002405482, 0.005812394, 0.005211085, 
    0.0002267944, -1.549124e-05, 0, 0, 0, 0, 0.0003030052, -0.0002752577, 
    -9.221906e-05, 0, 0, 0, 0, 0, 0, 0, 4.858511e-06, -0.0002106905, 
    0.008502989, 0, 0, 0,
  0, 0, 0.000384557, 0, 0, 0.001932089, 0, 0, -0.000210781, -0.0001497611, 
    -1.490287e-05, 0, -1.795409e-06, 0.0006798919, 0, 2.667694e-05, 
    -2.147711e-05, 0, 0, 0, 0, 0, 0, -5.065805e-05, 0, 0, 0.0004531548, 0, 0,
  0, 0, 0, 0, 0, -6.37561e-06, 0, 0.01362446, -5.154502e-05, 0.02035251, 
    0.004382352, 0.003448504, 0.008379173, 0.004328317, 0.001341067, 
    -7.452878e-06, 0.005897429, 0.0009891094, 0.0003304804, -0.000230651, 
    0.0207812, -1.077627e-05, -7.481362e-05, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0.000218756, 0, 0.003908889, -1.126152e-05, 
    -6.477616e-05, 0.002263756, 0, 0, 0, 0, 0, 0, 0, 0, 0.0009892328, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -3.01728e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -4.109701e-08, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -7.616509e-07, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, -1.482184e-06, 0, 0, 0,
  0, 0, 0, 0.0001037176, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.373621e-05, 0, 0, 0, 
    0, 0, -9.61254e-06, 0, 0, 0, 0, -6.150461e-05, 0.000901162, 0, 0, 0,
  0, 0, 0.004791455, 0.0005951847, -3.11393e-05, 0.001478019, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.001310419, 0, 0, -3.500959e-05, 0, 0, 0, 0, 0, 
    -2.189271e-05, -2.156946e-05, 0.0001951633, 0, 0,
  0, 0, -0.0001895246, -6.166042e-10, 0.003988993, 0.01014091, 0.01015225, 
    0.001127079, -3.098247e-05, 0, 0, 0, 0, 0.001059706, -0.0005020144, 
    -0.0002866606, -4.88868e-06, 0, 0, 0, 0, 0, 0, -2.196624e-05, 
    0.0007831771, 0.01029822, 0, 0, 0,
  0, 0, 0.001677622, 0, 0, 0.002018571, 0, 0, 0.004129824, -0.0002229474, 
    -4.47086e-05, 2.73046e-05, -1.694239e-05, 0.001346935, -4.902336e-06, 
    7.817036e-05, -9.534807e-05, 0, 0, 0, 0, 0, 0, -6.736117e-05, 
    6.336463e-05, 0.0005346485, 0.0005871645, 0, 0,
  0, 0, 0, 0, 0, -2.607558e-05, -6.243836e-05, 0.02233179, 0.005813565, 
    0.04122732, 0.00826993, 0.00371751, 0.01308238, 0.009495128, 0.004039722, 
    -0.0001001864, 0.007416434, 0.003538817, 0.001286132, -0.0006912503, 
    0.04022647, -3.002134e-05, -0.0001163767, 0, 0, -1.437039e-07, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0.0002522088, 0, 0.005802486, 4.988989e-05, 
    -7.557671e-05, 0.0031672, 0, 0, 0, 0, 0, 0, 0, 0.0002177431, 0.005034491, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -5.352573e-05, -1.551295e-05, 
    0.000581191, 0, 0, 0, 0, 0, 0, 0, 0.001139306, -2.743613e-06, 0, 
    0.0005304645, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0004801341, 0, -1.048891e-05, 
    0.000891608, 0, 0, 0, 0, 0, 0, 0, -8.087161e-06, -7.341774e-06, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, -6.236651e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, -5.367149e-05, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.0003580676, 0.001701285, -8.115748e-05, 0, 0,
  0, 0, -4.059235e-06, 0.0003102635, 3.753717e-05, 0, 0, 0, 0, 0, 0, 
    0.0006163734, 0, -0.0001134817, 0, 0, 0, 0.001360136, -9.484559e-05, 
    -0.0001055298, 0, 0, 0, 0, 0.0004612012, 0.004715836, 0, 0, 0,
  0, 0, 0.006740841, 0.001488461, -0.0001078343, 0.005535892, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.002410151, 0, -3.611661e-05, 0.0002670607, 0, 0, 0, 0, 0, 
    -7.091038e-05, 0.003341901, 0.001237264, 0, 0,
  0, 0, -0.0002562176, -1.890969e-08, 0.007444295, 0.01261289, 0.0172008, 
    0.004184233, 0.0002810458, 0, 0, 0, 0, 0.003500489, 0.000815735, 
    -0.0001766145, -5.944022e-05, 0, 0, 0, 0, 0, 0, 0.0002110816, 
    0.002213451, 0.01219379, 0, 0, 0,
  -3.076231e-05, 0, 0.003270106, 0, -9.744193e-06, 0.004578185, 0, 0, 
    0.007344851, 0.001795108, -6.448235e-05, 4.367763e-05, -7.145924e-05, 
    0.01024296, -2.454032e-05, 1.979995e-05, -0.0002837705, 0, -2.151585e-05, 
    0, 0, 0, 0, -8.075035e-05, 4.529551e-05, 0.002475319, 0.0005830638, 0, 0,
  0, 0, 0, 0, 0, 3.94258e-05, -0.0001200449, 0.03430549, 0.01662183, 
    0.06447767, 0.01600943, 0.007984004, 0.02110842, 0.02258063, 0.00872754, 
    -0.0002853379, 0.01186697, 0.006962501, 0.001505953, -0.001374763, 
    0.06440446, -2.172277e-05, -0.0003073101, 0, -5.023628e-06, 6.87611e-05, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0.002265744, 0, 0.009485468, 0.0009763713, 
    -0.0001755332, 0.003151362, 0, 0, 0, -3.166548e-06, -6.254662e-06, 0, 
    -2.718042e-06, 0.003525567, 0.007712469, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.004533172, 0.002118865, 0.004586464, 
    0, 0, 0, 0, 0, 0, 1.801163e-05, 0.00420699, -5.746516e-05, 0, 
    0.002393614, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -7.966552e-07, 0.003312907, 
    -3.039489e-05, 0.002124578, 0.002537173, 0, 0, 0, 0, 0, 0, 0, 
    0.001048731, 3.817324e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, -9.734036e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, -2.921837e-05, -1.78339e-05, 0, 0,
  0, 0, 0, 0.001946282, 0.001424572, 0.0003440448, 0, 0, 0, 0, 0, 0, 
    -1.64473e-05, 0.001380696, -3.434021e-06, 0, 0, 0, 0, -0.0001311078, 0, 
    0, 0, 0, 0.003359251, 0.006201142, 0.003456556, 0, 0,
  0, 0, 7.681078e-05, 0.00344835, 0.004157082, -9.26508e-05, 0, 0, 0, 0, 0, 
    0.004524142, -5.693854e-06, 0.002562027, 0, -3.316436e-06, 0, 
    0.009403303, 0.002652497, -0.0001813417, 0, 0, 0, 0, 0.005945095, 
    0.01610433, -9.127109e-08, -3.32253e-05, 0,
  0, 0, 0.01525193, 0.002727836, -0.0001562444, 0.01012014, -4.748216e-05, 0, 
    0, 0, -5.758722e-06, -3.560041e-08, 0, 0, -8.138883e-06, 0.008538725, 
    -7.564252e-06, 0.001986844, 0.003021439, 0, 0, 0, 0, -1.308245e-06, 
    0.001005968, 0.007509634, 0.005509499, 0, 0,
  0, 0, 0.0004449298, -9.887614e-06, 0.01922516, 0.02581805, 0.030532, 
    0.01387162, 0.001195671, 0, 0, 0, 0, 0.006820752, 0.002582189, 
    0.003942403, -0.0002020862, 0, 0, 0, 0, 0, 0, 0.0009064657, 0.008682114, 
    0.01600014, 0.0006327971, 0, 0,
  -4.002035e-05, 0, 0.01897469, -2.432186e-09, -3.753838e-05, 0.009852399, 
    -5.33426e-10, 0, 0.01167463, 0.006240416, 0.0003901376, 3.375742e-05, 
    -0.0001454118, 0.03165442, 0.001343612, 0.004215856, 0.0005087474, 
    3.153029e-06, 2.048682e-05, 0, 0, 0, 0, 0.003841741, 0.002743162, 
    0.004402543, 0.004845854, 0, 0,
  0, 0, 0, 0, -1.550853e-05, 0.0009632391, -0.0003525191, 0.04190522, 
    0.02670988, 0.09615953, 0.02946709, 0.01896486, 0.03776026, 0.03615946, 
    0.01660301, -0.0001198157, 0.02269075, 0.02257217, 0.004932927, 
    0.003069456, 0.1028031, -0.0002317211, -0.00102901, 0, -3.861402e-05, 
    0.0003305415, 0.0005767016, 0, 0,
  0, 0, 0, 0, 0, -2.261684e-06, 0, -7.336653e-06, 0.005174896, 0, 0.01408459, 
    0.006386482, 0.0002005832, 0.003255545, -6.57723e-06, 0, 0, 
    -7.569026e-05, -2.501865e-05, 0, 0.001596645, 0.007235433, 0.01274429, 0, 
    3.019419e-07, -1.290902e-05, 0, 0, 0,
  0, 0, 0, 0.0007540449, 0, 0, 0, 0, 0, 0, 0, -8.750779e-05, 0.005611707, 
    0.005662406, 0.007147373, 0, 0, 0, 0, 0, 0, 0.00424814, 0.007593501, 
    -0.0001504433, -5.53754e-05, 0.006299224, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0001397327, 0.006136945, 
    0.0005130512, 0.01072766, 0.004996285, 0.0009757314, -5.835487e-08, 
    -3.113991e-05, 0, 0, 0, -2.487872e-05, 0.003369251, 0.0009465045, 
    0.0003704653, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3.012009e-05, 
    -6.791722e-05, 0, 0, 0, 0, 0, 0.001582832, -2.997543e-06, 0.00315804, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -4.45469e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -1.34356e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.613128e-06, 
    0, 0, 0, 0, 0, 0, 0, 0,
  -1.875367e-05, -3.038348e-06, 0, 0, -8.686048e-05, 0.0004946779, 0, 0, 0, 
    0, 0, 0, 0, -2.24193e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0003786662, 
    -2.241914e-05, 8.971774e-06, -6.490588e-06,
  0, 0, 0, 0.0102185, 0.00920063, 0.007653547, -4.037576e-05, 0, 0, 0, 0, 
    -6.225898e-07, 0.0009234072, 0.00971758, 4.650073e-05, -9.031179e-06, 0, 
    0, 0, 0.002260146, 4.711381e-05, 0.002568043, 0, 0, 0.008411258, 
    0.01751779, 0.01260646, 0, -6.029258e-05,
  -1.837862e-06, 0, 0.001343931, 0.01191756, 0.01078852, 0.00317789, 
    3.347121e-05, 0, 0.0001290659, 9.191102e-06, 0, 0.007154637, 
    -3.304849e-05, 0.01215028, -3.899305e-05, -5.709876e-05, -0.0001488978, 
    0.0247, 0.02237939, -0.0004119718, -2.106439e-05, 0, 0, 0, 0.02115962, 
    0.02582122, 0.0005737991, -8.36695e-05, 0,
  0, 2.068553e-08, 0.02136192, 0.008362638, -0.0003163449, 0.01813748, 
    0.001775719, -1.008145e-07, 0, 9.874622e-07, -5.441043e-05, -9.39816e-06, 
    -2.823634e-10, -3.427896e-05, -0.0002852529, 0.01669042, 0.001288915, 
    0.0171775, 0.005608549, -4.43103e-06, 0, 0, 0, -6.054821e-05, 
    0.007113873, 0.01630545, 0.01784994, 4.702726e-05, 0,
  0, -2.681765e-05, 0.006010303, 0.0004708311, 0.03683618, 0.05366374, 
    0.0606382, 0.02820481, 0.002875446, -1.984988e-08, 0, -5.207233e-05, 
    -3.427834e-10, 0.04452328, 0.0232126, 0.01270793, 0.0005536469, 
    -2.63366e-10, 0, 0, 0, 0, 0, 0.01174584, 0.04762817, 0.0255664, 
    0.001747805, -2.509091e-09, 0,
  0.001290051, 0.001736126, 0.04404658, 0.000144515, -0.0001423012, 
    0.02677643, 1.656725e-06, -6.674936e-05, 0.03470143, 0.02404879, 
    0.005805368, 0.00168042, 0.0007813341, 0.0914354, 0.003473406, 
    0.008381633, 0.002806995, 4.919847e-06, 0.001417452, 0, 0, 7.509361e-09, 
    7.188237e-09, 0.02511821, 0.02067188, 0.006102168, 0.009323422, 
    -6.036341e-06, 0,
  0, 6.9459e-07, 0, 0, 0.0004541413, 0.001436365, 0.0005265686, 0.05812635, 
    0.03261847, 0.1262477, 0.04593166, 0.0316708, 0.08149969, 0.06539315, 
    0.02380003, 0.0008855704, 0.03789051, 0.04890068, 0.01968888, 0.01585695, 
    0.1431485, 0.001828356, 0.009727544, 0, -4.067549e-05, 0.0008487143, 
    0.0046813, 2.213861e-08, 0,
  0, 0, 0, 0, 0, -6.205794e-05, -4.762774e-06, -8.588837e-06, 0.009521919, 
    -1.940878e-06, 0.02608144, 0.02043301, 0.002830144, 0.004987338, 
    -1.147112e-05, 0, -3.982483e-05, -0.0001817096, -5.473704e-05, 
    -5.314127e-06, 0.00778431, 0.01756292, 0.01643561, 0, 9.83486e-05, 
    -1.008688e-05, 0, 0.0005883676, 0,
  0, 0, 0, 0.005009647, -5.091545e-06, 2.419885e-05, 0, 0, 0, 0, 
    2.848363e-07, -1.606575e-05, 0.006235494, 0.02120867, 0.01269601, 
    -2.320943e-08, 0.001022078, -9.441927e-06, 0, 0, -3.266401e-05, 
    0.01386809, 0.0151395, 0.0008399725, 0.001251051, 0.01656658, 0, 
    -6.23537e-05, 0,
  0, 0, 0, 5.804349e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0.0003306606, 0.01489532, 
    0.006720128, 0.02050925, 0.009134658, 0.006222547, 0.001634093, 
    0.0003294561, 0, 0, 0, -0.0001036687, 0.005726183, 0.002669178, 
    0.004312116, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -4.755406e-08, 0, 3.792136e-05, 0, 
    -7.195945e-05, 0.002963962, -2.123544e-05, -1.548031e-05, 0, 0, 0, 
    0.005704704, 0.0002521814, 0.006564423, -7.666667e-06, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -6.109159e-06, 0, 
    0, 0, 0, 0.001079577, 0.002870276, 0.00243989, 0, 3.173625e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -0.0001150767, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001153166, 0, 
    0, 0, 0, 0, 0, 0.0003567294, -1.247757e-05,
  0.003740207, 0.0001287526, -6.581405e-06, -6.625301e-05, 0.00324212, 
    0.002349998, 0.002106204, 0.004134176, -2.674689e-07, 0, 0, 
    -5.550784e-06, -7.271763e-06, 0.002680046, -7.793007e-06, 0.0005735473, 
    0.000113648, 0, -1.5639e-05, -6.690373e-05, 0, 0, 0, 0, -5.260281e-06, 
    0.004361048, 0.0006371081, 0.002805886, 0.001729278,
  -1.96365e-05, 0, -1.693519e-08, 0.02915853, 0.02114263, 0.02050002, 
    0.003354586, -8.02693e-05, -1.633367e-05, -6.028351e-05, 2.800823e-14, 
    -2.58893e-05, 0.003400127, 0.02132874, 0.004816475, 0.001280687, 0, 
    -1.124558e-05, -4.483698e-05, 0.008909622, 0.005015119, 0.01188201, 
    -7.07275e-05, -5.3976e-05, 0.02049077, 0.03167275, 0.03310662, 
    0.00163589, 0.0052065,
  -2.301635e-05, 0.0004384918, 0.005202848, 0.03611374, 0.02463109, 0.018983, 
    0.0002389573, 0.004765838, 0.002954297, 0.0001032971, -2.860135e-05, 
    0.0118458, -0.0002173897, 0.01725083, 0.002211494, 0.01276239, 
    0.002977935, 0.04255446, 0.05699868, 0.001323863, 0.003275487, 0, 0, 
    1.638007e-07, 0.031276, 0.03980508, 0.01412307, -0.000167778, 
    -9.433282e-06,
  2.562365e-08, 0.000181107, 0.06791972, 0.02270394, 0.002750908, 0.02508378, 
    0.01099851, 0.0005498833, 1.977729e-06, 0.0001596251, 0.001753583, 
    -4.009543e-05, -3.313664e-07, -4.68732e-05, 0.01163133, 0.03010506, 
    0.007494808, 0.04162095, 0.01485895, 0.0004060875, -4.476211e-10, 0, 0, 
    0.02246878, 0.0707856, 0.02899591, 0.03393842, 0.0004233837, -1.472263e-06,
  -4.422764e-11, 0.00849955, 0.04742683, 0.007087753, 0.04593288, 0.07048558, 
    0.1113396, 0.06285059, 0.01140515, -9.935185e-06, 1.252289e-06, 
    0.01044883, 0.001313109, 0.1285944, 0.1198332, 0.08420274, 0.002447208, 
    2.785845e-08, -1.664423e-08, -3.565811e-08, -1.172501e-08, 7.975465e-08, 
    -0.000143697, 0.06693155, 0.2044088, 0.07932063, 0.01418243, 
    0.0007834113, 6.448993e-09,
  0.005874776, 0.0125424, 0.1220703, 0.0007099456, -2.525254e-05, 0.03034457, 
    0.001155483, 6.454332e-05, 0.09609824, 0.07975656, 0.08585561, 
    0.03668619, 0.02249506, 0.1347563, 0.03905327, 0.02285357, 0.003975128, 
    -7.182883e-05, 0.00607218, 7.400185e-06, 2.295393e-06, 0.000128985, 
    0.0001501114, 0.1396324, 0.1917696, 0.009166745, 0.01194575, 
    -7.475317e-06, 0,
  -3.57103e-11, -9.209394e-05, -9.36999e-06, 0, 0.001462341, 0.01560365, 
    0.009451972, 0.07822575, 0.04983885, 0.2436959, 0.1558286, 0.1064319, 
    0.1824912, 0.1761735, 0.09416457, 0.02043523, 0.06029745, 0.0894689, 
    0.03518797, 0.04756565, 0.1935929, 0.02729672, 0.02062936, 0.001218973, 
    -6.506895e-05, 0.01187043, 0.007888572, 8.790406e-05, 0.0007722398,
  -1.478675e-06, 0, -3.457047e-09, 6.91207e-06, 0, 0.0006865326, 0.001142504, 
    0.0004747049, 0.01025634, -5.484931e-05, 0.07027469, 0.1240349, 
    0.04995586, 0.0269203, -5.513353e-05, 6.115117e-07, -9.710342e-05, 
    0.0008524745, 0.002824331, 0.005336012, 0.01621037, 0.0486293, 
    0.02358616, -5.640931e-05, 0.000137736, 0.0008544424, 0, 0.01014089, 
    -3.525831e-05,
  0, 0, 0, 0.009214593, 4.22568e-05, 0.005486727, -2.401517e-10, 0, 0, 
    0.0008989141, -1.995861e-06, 0.002402666, 0.03028681, 0.03795185, 
    0.02616699, 0.0009252583, 0.009746672, 0.001187931, 0.0002682132, 0, 
    -0.0001484967, 0.01887412, 0.04524383, 0.009712474, 0.005350229, 
    0.0282297, 0, -0.0001780564, 0,
  9.592339e-06, 0, 0, 0.001146621, -4.795828e-05, 0, 0, 0, 0, 0, 0, 
    -6.865176e-06, 0.008120947, 0.03038424, 0.01297606, 0.04897691, 
    0.02376376, 0.017219, 0.01485884, 0.001275244, 0, 0, 0, 0.007553624, 
    0.02568288, 0.008234063, 0.01106936, 0, 0,
  -1.104527e-05, 0, 0.0005112089, 0.001208398, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -0.0002599991, -1.007334e-07, 0.0008241602, 0, 0.004426427, 0.01112769, 
    -4.55205e-06, 0.00243966, 0, 0, 0.001739736, 0.01195252, 0.00128329, 
    0.0178246, 0.004719393, 0.0006535237,
  0.001072148, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.000270508, 0, 0, 0, 0, 0.006297116, 0.01402717, 0.006467094, 
    0.002528898, 0.00996557,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -3.697651e-05, -0.0001334577, 0, 0, 0, 0,
  0.0001554988, 0, -7.368421e-06, -3.31449e-06, 0, 0, 0, 0, 0, -7.828617e-07, 
    0, 0, 0, 0, 0, 0, 0, -6.252506e-06, 0, 0, 0.003566106, 0, 0, 0, 0, 0, 
    -1.453315e-05, 0.002444477, -8.952375e-05,
  0.01076776, 0.005268042, 0.000366166, 0.0006784419, 0.009709624, 
    0.00749501, 0.004398439, 0.01116947, 5.490446e-05, -8.503394e-08, 0, 
    -7.892521e-05, -3.663357e-05, 0.004226753, -4.165873e-05, 0.007505354, 
    0.0008031221, 0, -2.61266e-05, 0.000218779, 0, 0, 0.0003263787, 
    -2.3617e-06, 0.0003514467, 0.0077357, 0.006174792, 0.007331784, 
    0.007138398,
  0.008025887, -9.212475e-05, 0.000518959, 0.04968889, 0.07845191, 
    0.06216262, 0.0401977, 0.003929075, 0.0002564037, -0.000141265, 
    0.0001829655, -3.559686e-05, 0.009820119, 0.03287198, 0.01123, 
    0.004768496, 0.004642824, 1.164942e-05, 1.670924e-05, 0.03691727, 
    0.02136672, 0.03306147, 0.001898511, -6.310539e-05, 0.03925287, 
    0.0580776, 0.05929982, 0.02680711, 0.01819032,
  0.004816074, 0.004701349, 0.009889981, 0.1135021, 0.0742313, 0.08287819, 
    0.04306573, 0.01132566, 0.04550884, 0.03297481, 0.003253212, 0.02338343, 
    0.002262205, 0.02778368, 0.01037963, 0.02552914, 0.01392061, 0.09884863, 
    0.1215129, 0.04712928, 0.01680518, 0.001031628, 2.347231e-05, 
    2.331933e-05, 0.0667548, 0.121921, 0.05077785, 0.0100047, 0.02870894,
  0.0003966634, 0.004506301, 0.2938239, 0.06752072, 0.04680417, 0.0794851, 
    0.04894108, 0.003732258, 0.003647648, 0.02882892, 0.08675539, 
    -0.0001834297, 0.0006003434, 0.001317173, 0.05444065, 0.1131222, 
    0.1347119, 0.1986714, 0.1658065, 0.06718893, 0.0001273429, 0, 
    1.343094e-06, 0.05985807, 0.08974257, 0.1297449, 0.151964, 0.08458403, 
    0.03642458,
  1.456046e-06, 0.01056814, 0.3281356, 0.08314263, 0.07539208, 0.1096643, 
    0.1751336, 0.09559701, 0.05701135, 0.001981982, 0.0001023167, 0.03085193, 
    0.01928929, 0.1874728, 0.1687824, 0.1228075, 0.04000711, 0.0003901512, 
    9.093382e-08, -1.319538e-05, 4.051033e-07, -3.639161e-09, 1.629152e-05, 
    0.3797666, 0.2873378, 0.3714566, 0.09403146, 0.09058347, 0.0002415185,
  0.01546591, 0.1549133, 0.425423, 0.01827183, 0.01712717, 0.09697255, 
    0.03964818, 0.02359308, 0.2925806, 0.2423889, 0.1638321, 0.08854581, 
    0.06173537, 0.1402722, 0.02778196, 0.01385951, 0.005560545, 0.0001509889, 
    0.007326812, 1.568602e-05, 2.140401e-06, 0.0004480761, 0.01071784, 
    0.4539517, 0.3999971, 0.04396066, 0.01965826, 0.03275187, 5.893405e-07,
  7.872868e-07, 0.0010671, 0.005377447, -7.907386e-07, 0.007497771, 
    0.06654577, 0.06755011, 0.1145539, 0.06186572, 0.2876026, 0.1439973, 
    0.1033324, 0.2203377, 0.1781211, 0.08328594, 0.0537151, 0.1182423, 
    0.1916217, 0.08695163, 0.1277161, 0.2773388, 0.05756617, 0.100541, 
    0.009690759, 0.01004707, 0.08223042, 0.1722928, 0.02791287, 0.001863947,
  0.0007723938, 0.001083315, 0.0001426325, 3.590501e-05, -2.442657e-08, 
    0.01909045, 0.05718249, 0.04385236, 0.03782967, 0.004774961, 0.06754103, 
    0.08852608, 0.04228104, 0.05510524, 0.0003875746, 0.0001338441, 
    0.004184616, 0.01373547, 0.02855915, 0.06245377, 0.09230363, 0.1145101, 
    0.1478017, 0.1072589, 0.07892017, 0.04302141, 0.01232277, 0.1392265, 
    0.01112997,
  4.862785e-07, 0.0004984278, -1.312623e-06, 0.01957522, 0.000138349, 
    0.009741807, 0.0003348404, 0, -8.053058e-06, 0.08060164, 0.006851504, 
    0.01208529, 0.05139978, 0.08587327, 0.1056794, 0.06217799, 0.04684307, 
    0.008117273, 0.002860142, 0.0003338157, -0.0002059043, 0.02946303, 
    0.09726091, 0.06449431, 0.04963077, 0.06000888, 0.0002653739, 
    0.0007471933, -7.696152e-05,
  0.002952884, 0.002959773, 0, 0.002174477, -0.0005190375, -9.175997e-06, 0, 
    0, 0, 0, 0, -0.000159627, 0.02380385, 0.06184671, 0.03975942, 0.09577779, 
    0.04506159, 0.0402504, 0.03175554, 0.004289344, 0, 0, -1.262276e-06, 
    0.02145109, 0.04999487, 0.02007654, 0.02888784, 0.0008630113, 0,
  -1.868866e-05, -1.445897e-05, 0.004181766, 0.002186071, 0, 0, 0, 0, 0, 0, 
    0, 0, -0.0001663668, 0.00226397, 0.003931551, 0.006358494, 0.001405512, 
    0.02020851, 0.0210812, 0.004231137, 0.003375329, -1.295895e-07, 0, 
    0.007560736, 0.02414345, 0.008657781, 0.02651706, 0.0132767, 0.005060207,
  0.004673984, 7.843074e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -2.27239e-05, 0.001239228, 0.0006386964, -1.208111e-05, 0, 0.0004009787, 
    0.01143899, 0.03330597, 0.01564437, 0.01173144, 0.01875792,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2.578581e-06, -0.0001627109, 0.002243165, 0, 0, 0, 0,
  0.008659071, 9.092537e-05, 6.465008e-05, -4.082897e-05, 8.265464e-05, 
    -1.872644e-05, 0.001554154, 3.151779e-05, 4.391294e-05, 0.002231956, 
    -1.395021e-06, -6.833215e-06, 0, 0, -0.0001110072, -3.828433e-05, 
    8.922166e-05, 0.0005880031, 0.002418682, -3.053805e-05, 0.006087746, 
    -4.760985e-05, -5.327143e-06, 0, 0, 0, 0.0001002097, 0.003560809, 
    0.006159277,
  0.03045572, 0.01421994, 0.007513675, 0.002421389, 0.01759134, 0.02094441, 
    0.02660605, 0.02173089, 0.02498958, 0.008583684, 0.001312889, 
    2.654807e-05, 0.001837608, 0.01097006, 0.0007612581, 0.01013352, 
    0.01205081, 0.008353434, -0.0001010471, 0.00531673, 0.005384744, 
    -1.240804e-05, 0.002108499, 1.471309e-05, 0.002322501, 0.02021431, 
    0.0404448, 0.04044396, 0.0356401,
  0.02093539, 0.004523375, 0.02038264, 0.08983311, 0.1305717, 0.1201972, 
    0.08671548, 0.01899313, 0.02664459, 0.01871417, 0.04368904, 0.02404488, 
    0.03606716, 0.04552817, 0.0305546, 0.04271226, 0.01982331, 0.005195023, 
    0.02968983, 0.1186774, 0.09300931, 0.08182205, 0.01561993, 0.000376591, 
    0.06860007, 0.1321121, 0.1189801, 0.07653578, 0.07737871,
  0.01360103, 0.0431223, 0.04717094, 0.09136803, 0.09815906, 0.09506576, 
    0.07566839, 0.08163811, 0.1082288, 0.1058603, 0.08323286, 0.08824385, 
    0.04710558, 0.05347407, 0.04011267, 0.07297069, 0.06878182, 0.1687846, 
    0.3443878, 0.1968797, 0.1129044, 0.08487926, 0.008074822, 0.00567111, 
    0.07784537, 0.1068765, 0.1008221, 0.06952322, 0.06967559,
  -1.219564e-05, 0.0009439497, 0.3064454, 0.05809986, 0.0332898, 0.07264819, 
    0.02442744, 0.009094932, 0.0007120072, 0.04425474, 0.08191695, 
    0.01336826, 0.004068125, 0.00708559, 0.07054061, 0.1275969, 0.1226353, 
    0.2246041, 0.1368353, 0.0575902, 0.002797584, 1.641956e-05, 
    -1.379094e-09, 0.05280044, 0.07897534, 0.1373253, 0.1543925, 0.1142618, 
    0.02980757,
  1.118115e-07, 0.004378519, 0.2925869, 0.06841445, 0.05841985, 0.08590499, 
    0.125441, 0.07579558, 0.0497682, 0.002036888, 6.323379e-05, 0.01050214, 
    0.01101171, 0.1470302, 0.1362743, 0.09326728, 0.02813209, 0.002001502, 
    -8.661013e-07, 3.20127e-07, 5.090902e-08, 1.668911e-09, 5.152373e-06, 
    0.289963, 0.2381396, 0.3328467, 0.08037004, 0.09358747, 3.84076e-05,
  0.01203472, 0.115356, 0.3589218, 0.01194757, 0.007160728, 0.05676498, 
    0.01631056, 0.01172925, 0.2336246, 0.1852177, 0.1047778, 0.05420517, 
    0.02545814, 0.1234351, 0.0249228, 0.01549186, 0.003815608, 7.786136e-05, 
    0.001749879, 6.382476e-06, 2.16758e-07, 1.323718e-06, 0.01434706, 
    0.3655283, 0.2999607, 0.03232428, 0.02195846, 0.01132167, 4.114681e-07,
  6.162768e-07, 0.001044591, 0.0001383623, 1.112549e-06, 0.001454116, 
    0.05111759, 0.04692981, 0.09076073, 0.05755567, 0.2412467, 0.1142232, 
    0.07780132, 0.1928709, 0.1462752, 0.06472564, 0.03240473, 0.09352824, 
    0.1306351, 0.07342921, 0.09517115, 0.2326274, 0.02876434, 0.0737231, 
    0.004204443, 0.005886056, 0.04903048, 0.1259908, 0.02299369, 0.003223338,
  0.07571788, 0.01589895, 7.701507e-06, 6.279794e-06, 1.88595e-08, 
    0.006971437, 0.07209388, 0.03304332, 0.02642912, 0.002912074, 0.06266247, 
    0.06000317, 0.02692653, 0.03797192, 0.002014232, 0.01164439, 0.002801437, 
    0.01422211, 0.01286532, 0.04417153, 0.06412129, 0.1137527, 0.1150132, 
    0.06057466, 0.04181134, 0.06876171, 0.07932207, 0.1512955, 0.07756981,
  0.009303592, 0.005812969, 0.003587182, 0.04107188, 0.0005294054, 
    0.01770786, 0.008678513, 0, 0.0006397555, 0.08685955, 0.01395037, 
    0.03759871, 0.0664504, 0.1145301, 0.1452237, 0.1262353, 0.1663871, 
    0.08975916, 0.08434916, 0.03630435, 0.005641822, 0.06003262, 0.1849558, 
    0.120733, 0.152054, 0.2014581, 0.07010896, 0.01618887, 0.03457034,
  0.006117287, 0.004028312, 0.0001882954, 0.006995122, 0.009935742, 
    0.0002438112, -4.749696e-06, -1.864161e-06, 0, -1.090295e-10, 
    -1.094435e-10, 0.000896254, 0.04254471, 0.08660222, 0.06896493, 
    0.1369726, 0.1043674, 0.124096, 0.1005134, 0.01688444, -4.302613e-05, 
    0.0007400324, 0.000873338, 0.03178234, 0.08299302, 0.08305277, 0.1441511, 
    0.01221518, 0.000117817,
  0.0002553705, 0.001835442, 0.009506101, 0.006319691, -0.0001008813, 
    -1.677285e-08, 0, 0, 0, 0, 0, 0, 0.001096037, 0.008339176, 0.02419878, 
    0.0245687, 0.0172208, 0.07797246, 0.07215928, 0.01591776, 0.0067605, 
    0.003413013, 0.0001773588, 0.01087227, 0.04579046, 0.04272497, 
    0.06015475, 0.04646567, 0.02718939,
  0.01013956, 0.001114965, 0, 0, 0.0001203925, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, -0.0001460297, 0.002580728, 0.005053454, 0.003403256, 0.0003604788, 
    0, 0.006776928, 0.02285867, 0.07391331, 0.03002011, 0.03097033, 0.03153307,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.00178252, -3.465236e-06, 0, -1.634262e-08, -7.514525e-06, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -9.072273e-06, 0.002616292, 
    0.0007390106, -2.952011e-10, 7.310426e-05, 0, -3.626998e-06, 0.003117597, 
    0.003578948, 0, 4.494438e-05, 0, 0,
  0.01349686, 0.01129442, 0.01107241, 0.0006430735, 0.002505741, 0.005408875, 
    0.007748661, 0.01013305, 0.02466453, 0.02184042, 0.004600161, 
    0.005354648, 0.0223894, 0.0234747, 0.006286492, 0.001513086, 0.008750297, 
    0.01131962, 0.01736902, 0.01829854, 0.01872293, 0.004364384, 
    0.0007692752, 5.000504e-05, -2.05857e-05, 0, 0.004013192, 0.006050196, 
    0.01358416,
  0.05302673, 0.05944104, 0.05730886, 0.06035867, 0.1013556, 0.08762532, 
    0.09032536, 0.04728817, 0.08283479, 0.05683761, 0.07491574, 0.1063903, 
    0.09477825, 0.1054373, 0.0541232, 0.04466442, 0.05366822, 0.02680457, 
    0.008423823, 0.01576644, 0.02895934, 0.03188745, 0.02110512, 
    0.0005668062, 0.02127297, 0.05911022, 0.08319589, 0.07101078, 0.0605936,
  0.05847541, 0.03648781, 0.04812347, 0.1194951, 0.1511889, 0.1352128, 
    0.121574, 0.1007921, 0.1088905, 0.115963, 0.1480903, 0.1140277, 
    0.07879575, 0.1150766, 0.05969343, 0.08640768, 0.05374043, 0.03199764, 
    0.07554511, 0.1625246, 0.1362943, 0.1401361, 0.09433262, 0.02686581, 
    0.1475935, 0.1451989, 0.1371308, 0.1188097, 0.1482882,
  0.006373024, 0.02420734, 0.06047114, 0.06817136, 0.09888384, 0.07442166, 
    0.05422228, 0.08862573, 0.09990249, 0.08717826, 0.06100263, 0.08471557, 
    0.05290618, 0.0589279, 0.06688678, 0.0940389, 0.1470369, 0.1747146, 
    0.3280502, 0.1464633, 0.114805, 0.07540171, 0.01046664, 0.002920497, 
    0.07505549, 0.1008569, 0.08725386, 0.07245976, 0.05781408,
  -1.111373e-05, -3.304499e-05, 0.2874764, 0.06487323, 0.03635458, 
    0.07498408, 0.01792129, 0.01422575, 4.230119e-05, 0.05232945, 0.08355428, 
    0.008128363, 0.0008374713, 0.02570108, 0.06060832, 0.09952943, 0.1190347, 
    0.16265, 0.1022126, 0.03084936, 0.000295892, 2.616131e-07, -4.536911e-09, 
    0.0352357, 0.05696344, 0.1325347, 0.1227727, 0.07343149, 0.0122667,
  4.481554e-08, 0.002417525, 0.2605086, 0.06982276, 0.05271034, 0.07798887, 
    0.1097131, 0.06845556, 0.05209331, 0.00473454, 0.000663606, 0.006411043, 
    0.006798691, 0.1314365, 0.1139705, 0.08042601, 0.03200291, 0.0005059493, 
    -1.636272e-06, -1.707257e-08, -4.444375e-11, 3.059035e-08, 2.372207e-06, 
    0.2438587, 0.2072575, 0.3049331, 0.06597167, 0.08322082, 3.327897e-06,
  0.01312585, 0.1009845, 0.3117535, 0.010113, 0.007462893, 0.04363663, 
    0.01456653, 0.006894216, 0.1958946, 0.1583855, 0.07325826, 0.03506427, 
    0.02582036, 0.1194839, 0.02979737, 0.0159119, 0.002802948, 1.325678e-05, 
    0.001376075, -7.139792e-06, 4.550326e-07, 5.075317e-08, 0.00944315, 
    0.3311471, 0.2331669, 0.03686913, 0.02496823, 0.00246095, 0.0001175268,
  3.128001e-07, 0.0001574763, 1.012561e-05, 2.197645e-06, 0.002805551, 
    0.05052007, 0.0416219, 0.08275598, 0.06405061, 0.2063776, 0.1068512, 
    0.07422764, 0.1744219, 0.1315739, 0.05691646, 0.02493578, 0.07471711, 
    0.09885309, 0.06683533, 0.07480904, 0.2100353, 0.03327755, 0.04939712, 
    0.002611958, 0.006097383, 0.03757577, 0.08506035, 0.01228763, 
    -0.0001481986,
  0.03834434, 0.002517017, 2.331427e-07, 1.658603e-05, -2.871932e-08, 
    0.005168491, 0.0877745, 0.01109758, 0.02009386, 0.002187932, 0.07511994, 
    0.04707058, 0.02171066, 0.02898862, 0.003126224, 0.01233322, 0.001871052, 
    0.007486592, 0.0224473, 0.03743071, 0.03416256, 0.102231, 0.0838036, 
    0.03069591, 0.02863461, 0.04705205, 0.05593177, 0.1289055, 0.0718575,
  0.04158679, 0.04052137, 0.03154991, 0.03430473, 0.002553596, 0.02408521, 
    0.09016042, -5.892181e-05, 0.006251445, 0.08075113, 0.02150647, 
    0.0860356, 0.1049625, 0.1394537, 0.1280925, 0.1256242, 0.1516445, 
    0.106832, 0.131411, 0.06162343, 0.04023376, 0.0974107, 0.1748772, 
    0.1157688, 0.1183987, 0.1629394, 0.05342557, 0.0513003, 0.08439407,
  0.02140691, 0.01394266, 0.02739889, 0.01308461, 0.02764263, 0.01878173, 
    0.0007694004, 0.004827631, -4.093432e-05, 4.337597e-05, 0.001967102, 
    0.01358868, 0.05740741, 0.1117725, 0.1046464, 0.164913, 0.1626719, 
    0.2398811, 0.1586628, 0.07860999, 0.002694919, 0.02258568, 0.0405231, 
    0.06594985, 0.1537573, 0.1601765, 0.2586786, 0.1122364, 0.04408746,
  0.02825641, 0.008995084, 0.01821043, 0.01228585, 0.00270542, 0.006211543, 
    -5.303482e-06, -4.132373e-07, 0, 0, 0, 0, 0.004304739, 0.01569987, 
    0.02632095, 0.02738418, 0.05371448, 0.183829, 0.239646, 0.0432295, 
    0.02420789, 0.02184164, 0.01384308, 0.02247762, 0.06797303, 0.06621035, 
    0.1250889, 0.1059339, 0.07109351,
  0.03449697, 0.008972597, -2.864094e-05, 0.0001704117, 0.0009410017, 
    0.001426439, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.00093806, -7.754694e-05, 
    0.005800352, 0.0112627, 0.007691371, 0.0136769, 0.009687318, 
    -0.0002359918, 0.007423669, 0.04753295, 0.1173478, 0.08915057, 
    0.06200158, 0.05611029,
  0, 0, 0, 0, 0, 0, 0.0002064675, 0, 0, 0, 0, 0, 0, 0, 0, -4.35931e-06, 
    2.653058e-06, 0, 0, 0, 0, 0, -0.0002586897, 0.003652444, 9.141336e-05, 0, 
    -5.679619e-08, -9.111867e-05, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  -7.892619e-06, -0.0005108424, 0.009830098, -3.587672e-05, -6.46908e-06, 0, 
    0.0003422015, -0.0001319059, 0, 0, 0, 0, -4.615282e-08, 0.0005973129, 
    0.0004906566, -3.696458e-05, 0.001918807, 0.00437668, 0.004978233, 
    -0.0001863235, -3.329918e-05, -0.0002394845, 0.009885629, 0.01643889, 
    0.02384676, 0.01121042, 0.01047628, 0.0003573072, 0,
  0.03304981, 0.04240259, 0.04679447, 0.04921966, 0.04868448, 0.03751125, 
    0.02918722, 0.04057757, 0.03315749, 0.04302765, 0.02467344, 0.04562014, 
    0.0830193, 0.1120049, 0.09790692, 0.08588923, 0.09534907, 0.07563088, 
    0.05490593, 0.03017087, 0.04075225, 0.04107774, 0.04399638, 0.03341165, 
    0.02402605, 0.01908782, 0.01738594, 0.02823799, 0.0394077,
  0.08447759, 0.0876316, 0.1304538, 0.1432028, 0.147443, 0.1295735, 
    0.1127072, 0.09939063, 0.1765606, 0.1590094, 0.1564372, 0.1906927, 
    0.2139096, 0.1931259, 0.1596734, 0.1183944, 0.09893739, 0.09568539, 
    0.08256858, 0.06582857, 0.07339755, 0.08118024, 0.06058072, 0.02409904, 
    0.09178775, 0.1552256, 0.1308264, 0.1274963, 0.08676156,
  0.06995554, 0.05189441, 0.05133912, 0.09863225, 0.1286232, 0.1333396, 
    0.1322695, 0.1004639, 0.1037561, 0.1129147, 0.1319271, 0.09770522, 
    0.09963949, 0.1324442, 0.08316999, 0.09893356, 0.07659228, 0.03649738, 
    0.08323836, 0.1632202, 0.1345301, 0.1558992, 0.1320612, 0.08973957, 
    0.1377954, 0.1365069, 0.1378925, 0.1308962, 0.1595523,
  -0.0001574619, 0.003016579, 0.04564988, 0.05421738, 0.1085346, 0.05633555, 
    0.0354147, 0.07754568, 0.09304737, 0.06459838, 0.03246157, 0.07660879, 
    0.04133062, 0.06095235, 0.04201703, 0.07970873, 0.09994201, 0.1547817, 
    0.3038807, 0.09719442, 0.08931856, 0.07006169, 0.0139597, 0.000749388, 
    0.06364161, 0.07999834, 0.1002726, 0.06610397, 0.06940973,
  3.088692e-09, -6.589333e-05, 0.284452, 0.08646201, 0.03575466, 0.07670464, 
    0.01380458, 0.004726458, 8.91771e-06, 0.02773839, 0.07059085, 
    0.004836723, 0.0009225212, 0.02157936, 0.04832157, 0.09636484, 0.1155582, 
    0.1341326, 0.08049943, 0.003647903, 0.0003867278, -5.147342e-09, 
    -1.37979e-10, 0.01671127, 0.04255474, 0.1321613, 0.09727899, 0.03399974, 
    0.00593065,
  3.64563e-08, 0.001082582, 0.2183947, 0.05974843, 0.04775841, 0.07661659, 
    0.09615314, 0.05513141, 0.05166372, 0.0039485, 0.00126129, 0.004055062, 
    0.006633011, 0.1001353, 0.08873498, 0.0651511, 0.04273936, 0.000531368, 
    1.892302e-07, -3.29556e-08, 0, 3.109789e-08, 1.029607e-06, 0.1900148, 
    0.1659783, 0.2564289, 0.06870311, 0.05074712, 4.897547e-07,
  0.01689642, 0.07281305, 0.266137, 0.01052015, 0.01448276, 0.03784459, 
    0.01256386, 0.005908403, 0.1551905, 0.1399189, 0.04514739, 0.0261606, 
    0.02106959, 0.09896853, 0.03206777, 0.01764062, 0.002899048, 
    -5.777004e-06, 0.001506483, -2.281728e-05, -5.315784e-07, 2.19215e-07, 
    0.0008325608, 0.2859666, 0.1485849, 0.04630151, 0.0296184, 0.0007349938, 
    0.0001210935,
  -3.0025e-06, 4.115868e-05, 1.950307e-05, -1.688335e-06, 0.00165732, 
    0.04342606, 0.03153418, 0.07605139, 0.07042144, 0.1927637, 0.09978836, 
    0.05980494, 0.1494821, 0.1107308, 0.04279375, 0.02034479, 0.06451146, 
    0.08181094, 0.04980334, 0.06937349, 0.190542, 0.02698606, 0.02674394, 
    0.00312026, 0.007126041, 0.03296196, 0.06717535, 0.00496472, -7.636005e-05,
  0.01483194, 0.0001358239, 1.285383e-06, 2.559991e-05, -8.116708e-09, 
    0.007173707, 0.06100815, 0.005113334, 0.02165849, 0.0001886222, 
    0.0851112, 0.03787654, 0.01726785, 0.01992802, 0.003867469, 0.008730022, 
    0.0003180015, 0.008422597, 0.0123393, 0.04132157, 0.0353854, 0.1158959, 
    0.06702694, 0.0222962, 0.02121643, 0.04336422, 0.0354143, 0.1277205, 
    0.04423133,
  0.02195087, 0.04336431, 0.03658558, 0.03736171, 0.01107593, 0.05411223, 
    0.09469368, 0.0007725556, 0.01092182, 0.0815049, 0.02867473, 0.1281442, 
    0.1011076, 0.1284105, 0.1054199, 0.1104397, 0.116927, 0.09292804, 
    0.1096446, 0.02941801, 0.04757455, 0.07471445, 0.130209, 0.09197572, 
    0.08330097, 0.1347042, 0.03752138, 0.03493019, 0.097619,
  0.07924689, 0.07193, 0.07127202, 0.04824021, 0.1297501, 0.1101274, 
    0.002650505, 0.04324149, 0.01738683, 0.005358694, 0.02626625, 0.04389832, 
    0.0965214, 0.1464842, 0.1340103, 0.1661234, 0.1737485, 0.2429191, 
    0.1451233, 0.1275687, 0.04053028, 0.0616618, 0.1288154, 0.1453488, 
    0.2131393, 0.1606678, 0.2711643, 0.09820449, 0.05420779,
  0.07559486, 0.04751449, 0.03729066, 0.08419912, 0.1286814, 0.07534134, 
    0.001976745, -1.090394e-05, 0, -1.889141e-05, 0.009866571, 0.001675196, 
    0.01216194, 0.03200559, 0.03374033, 0.04802344, 0.08803175, 0.2459907, 
    0.3063144, 0.1440306, 0.07385024, 0.09568462, 0.0393503, 0.03891011, 
    0.1129218, 0.1329434, 0.1464205, 0.1319337, 0.1020842,
  0.08234154, 0.02582994, -0.0001533713, 0.004380743, 0.01047842, 0.02257996, 
    0.004519836, 2.260473e-06, 0.0001373365, 0, 0, 0, 0, -1.702007e-07, 
    -0.0003669443, 0.08572534, 0.009014847, 0.02937358, 0.02474541, 
    0.04190406, 0.03060505, 0.01416789, 0.007118914, 0.01630675, 0.06327779, 
    0.1334715, 0.1363679, 0.1500985, 0.1013558,
  0, -5.74356e-05, -9.172221e-06, 0, 0, 0, 0.003782662, 0, 0, 0, 0, 0, 0, 0, 
    0.02715725, 0.03964036, 0.01492459, 0.03411014, 0.005264825, 2.51435e-05, 
    0, -0.0007456857, 0.01505113, 0.02003514, 0.04072223, -0.0001581514, 
    -3.623958e-05, 0.02475664, -2.022717e-06,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3.918193e-06, 0.001869683, 
    6.21852e-05, 0.002463736, 0.0004954731, -0.0001199565, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  -5.674686e-05, 0.008014745, 0.02856519, 0.01826734, -0.0001520454, 
    -0.0005888753, 0.01333427, -0.0001656139, 0, -8.459041e-05, 
    -5.274783e-07, 0, -0.0006440119, 0.009391468, 0.01780951, 0.03212629, 
    0.03117627, 0.05612569, 0.04439236, 0.04184822, 0.01877985, 0.006583233, 
    0.01195224, 0.03010892, 0.05012307, 0.04739866, 0.03553926, 0.02254797, 
    0.0003518299,
  0.09926231, 0.1138812, 0.07521887, 0.121, 0.1306934, 0.09676436, 
    0.08794773, 0.0794951, 0.04982257, 0.09759466, 0.06639928, 0.09857286, 
    0.1287823, 0.1389377, 0.1480068, 0.1391486, 0.1452644, 0.1489628, 
    0.1231171, 0.1342809, 0.1439849, 0.1682645, 0.164607, 0.1179088, 
    0.08633975, 0.06375992, 0.07961521, 0.1198379, 0.1156109,
  0.09659167, 0.129427, 0.1457135, 0.1604275, 0.1424942, 0.1187777, 
    0.1176391, 0.1177472, 0.1938844, 0.1769329, 0.1877576, 0.184309, 
    0.229179, 0.1668945, 0.155581, 0.1159351, 0.123377, 0.1197063, 0.1123317, 
    0.09222706, 0.1098263, 0.111175, 0.1128743, 0.1057138, 0.1385237, 
    0.1944368, 0.129844, 0.1512891, 0.1272507,
  0.05346339, 0.05555132, 0.04157721, 0.07570361, 0.1112868, 0.1148655, 
    0.1323031, 0.08749726, 0.09252344, 0.1256595, 0.1250323, 0.0932873, 
    0.08156017, 0.1300684, 0.07927009, 0.08111612, 0.06844429, 0.0342598, 
    0.06850971, 0.15105, 0.1406134, 0.1709272, 0.118297, 0.08502563, 
    0.1224928, 0.142875, 0.1303006, 0.1565256, 0.1345906,
  -9.775006e-05, 0.0004108813, 0.03590857, 0.04561349, 0.08817719, 
    0.04647041, 0.04971461, 0.06146379, 0.0759482, 0.05832706, 0.0256496, 
    0.0690084, 0.03772671, 0.06325801, 0.03407597, 0.06207906, 0.0750022, 
    0.1306536, 0.2733037, 0.09215876, 0.06543244, 0.05297507, 0.006768879, 
    0.0002444825, 0.05421855, 0.06056203, 0.1004105, 0.05790256, 0.02607208,
  3.711708e-07, -4.30313e-06, 0.2653553, 0.1070767, 0.03494677, 0.0715323, 
    0.01253911, 0.005422692, 2.199296e-05, 0.007168591, 0.04785446, 
    0.003137928, 0.0007303464, 0.01457699, 0.03839374, 0.09888228, 
    0.07935791, 0.1151218, 0.0668704, 0.0004017341, 1.661053e-05, 
    2.826336e-08, 0, 0.00864108, 0.03020074, 0.1314528, 0.09339622, 
    0.02157241, 0.001911857,
  1.993783e-08, 0.002486639, 0.1710453, 0.03931891, 0.04414093, 0.07732982, 
    0.09025773, 0.05877992, 0.04835686, 0.003427035, 0.001150857, 
    0.002520374, 0.006093576, 0.07150537, 0.05413342, 0.0563943, 0.02364456, 
    0.0003597635, 1.296697e-07, -6.986478e-09, 0, 1.329153e-08, 9.151195e-07, 
    0.1376183, 0.1449104, 0.2109693, 0.06715252, 0.01049991, 1.103641e-07,
  0.02243192, 0.05061164, 0.2153673, 0.006935881, 0.01548054, 0.03335953, 
    0.01375413, 0.009162051, 0.1182106, 0.1229994, 0.03003746, 0.02450325, 
    0.01811899, 0.07110938, 0.03338672, 0.02013945, 0.005589215, 
    -2.397548e-05, 0.0004464486, -2.013728e-05, -8.577517e-08, 5.442418e-08, 
    3.124769e-05, 0.2293746, 0.07754892, 0.06263703, 0.04914639, 
    0.0003863381, 3.437547e-05,
  0.0001596785, 2.085833e-05, 3.102473e-05, -1.129445e-05, 0.002009566, 
    0.03922701, 0.02010216, 0.07285618, 0.07507494, 0.1892142, 0.09572846, 
    0.04740021, 0.1232642, 0.09516522, 0.04202851, 0.01274944, 0.05722785, 
    0.05936666, 0.03148892, 0.08944688, 0.1832748, 0.02255052, 0.01876248, 
    0.002760217, 0.005216217, 0.03521105, 0.06041108, 0.000946202, 
    -0.0002333564,
  0.0321065, 1.895167e-05, 9.45805e-07, 6.632848e-05, -7.052741e-09, 
    0.007837232, 0.04979252, 0.004158575, 0.0268445, -0.000345947, 
    0.08549426, 0.03202305, 0.01181702, 0.01516824, 0.0006312479, 
    0.000753996, -0.0003485955, 0.005547926, 0.005234409, 0.02680941, 
    0.03790133, 0.1255693, 0.0680076, 0.01770662, 0.01407689, 0.03914423, 
    0.02037843, 0.121943, 0.03191247,
  0.02098357, 0.03405415, 0.0390906, 0.044831, 0.02846454, 0.0503113, 
    0.06991462, 0.004728409, 0.04042435, 0.08220706, 0.03417745, 0.1007105, 
    0.09672194, 0.112595, 0.09761545, 0.09360562, 0.0921995, 0.07254596, 
    0.04926131, 0.0238202, 0.02996269, 0.04396532, 0.1051891, 0.06421729, 
    0.0691858, 0.1219558, 0.04610643, 0.02848078, 0.1002826,
  0.0907931, 0.09650216, 0.1251801, 0.1533537, 0.1513631, 0.132731, 
    0.02215178, 0.08074233, 0.03919027, 0.0214376, 0.04439756, 0.0879935, 
    0.1123879, 0.1573104, 0.1468049, 0.180161, 0.1803214, 0.2268908, 
    0.1353914, 0.1252127, 0.08481055, 0.08322102, 0.1447413, 0.1371135, 
    0.2067266, 0.1350239, 0.2899168, 0.07906706, 0.05474074,
  0.1091119, 0.08769866, 0.1350788, 0.2321837, 0.2769288, 0.232079, 
    0.08328465, -0.0003187782, 0.001196307, 0.01927773, 0.03106788, 
    0.01661458, 0.05152483, 0.07698082, 0.07169896, 0.1096302, 0.1405445, 
    0.2960274, 0.3123088, 0.1956098, 0.1086344, 0.1145641, 0.09457696, 
    0.07726388, 0.1614495, 0.1706473, 0.1733553, 0.1507627, 0.1184494,
  0.1071539, 0.06986889, 0.02385349, 0.03056527, 0.07121112, 0.1262304, 
    0.1860344, 0.1814701, 0.06115345, 0.01597679, 0, 0, 0, 0.0002400521, 
    0.07765108, 0.1733688, 0.07077899, 0.05350551, 0.105773, 0.08354387, 
    0.08135707, 0.06610595, 0.06382104, 0.04172414, 0.07940546, 0.1478778, 
    0.1760746, 0.1814003, 0.1258134,
  0.006509838, 0.02523616, 0.004251216, 0.001486227, -0.0004740171, 
    0.01395742, 0.01964634, 0.002449227, 0.0007368917, 0, 0, -5.079111e-07, 
    0, 0.002110511, 0.0604783, 0.07635694, 0.09122036, 0.1000087, 0.04920124, 
    0.01000128, 0.0005335524, 0.01659741, 0.03909488, 0.0360156, 0.04702302, 
    0.00465815, 0.0003112444, 0.09182393, 0.02042543,
  0.006477085, -0.0001905688, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002044789, 
    0.02998308, 0.02956706, 0.03225423, 0.02792385, 0.02053668, 0.0002950632, 
    0, -2.292321e-05, -0.000244273, -0.001811367, 0.001069915, -1.105666e-08, 
    0, -0.00159213, 0.01046652,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3.799187e-06, 0, 0, 0, 0, 
    0, -2.075288e-09, -0.000112781, 0.00114392, -0.003210101, -0.0008072607, 
    0, 0,
  0.05943179, 0.1145319, 0.1070337, 0.06258769, 0.0009141924, 0.002273385, 
    0.02307076, 0.001262497, -0.000182067, -0.0002723373, -4.832536e-05, 
    -2.254807e-05, 0.00256994, 0.04559511, 0.08308709, 0.07196734, 0.1128686, 
    0.1048591, 0.08524744, 0.07977094, 0.07494722, 0.06744418, 0.07521731, 
    0.1133289, 0.1074655, 0.1112944, 0.1210105, 0.1104272, 0.07322051,
  0.1528754, 0.1823187, 0.1110691, 0.1751122, 0.1939418, 0.1847008, 0.137265, 
    0.08679435, 0.07316837, 0.137068, 0.1124141, 0.115611, 0.1343448, 
    0.17083, 0.1982164, 0.2130691, 0.1940945, 0.1912608, 0.1522516, 
    0.1717874, 0.177587, 0.2035878, 0.2097275, 0.2023127, 0.1599343, 
    0.1176154, 0.1286642, 0.1422359, 0.1461168,
  0.0987001, 0.1380901, 0.1501279, 0.1824825, 0.1542565, 0.1305926, 
    0.1250093, 0.1275045, 0.1856633, 0.1871693, 0.1996816, 0.166535, 
    0.2116231, 0.1573918, 0.1568045, 0.107108, 0.1180106, 0.1235918, 
    0.1118306, 0.1042461, 0.131923, 0.1055867, 0.1290112, 0.1483182, 
    0.1429578, 0.1967349, 0.1697157, 0.1502986, 0.1268428,
  0.04600144, 0.06081542, 0.03550551, 0.06951264, 0.09017166, 0.1102845, 
    0.1309395, 0.09179627, 0.0906747, 0.1312324, 0.1117865, 0.08930111, 
    0.06298254, 0.1268074, 0.07893299, 0.08648706, 0.06783137, 0.04077141, 
    0.05655969, 0.1450607, 0.1514265, 0.167271, 0.1409836, 0.08579483, 
    0.1132717, 0.132326, 0.1274688, 0.1571929, 0.1222663,
  0.0006719691, 0.0001894431, 0.02812647, 0.04766101, 0.06753791, 0.06049599, 
    0.03586632, 0.04380478, 0.05826459, 0.03803545, 0.03577097, 0.0732611, 
    0.03642105, 0.06149088, 0.02944738, 0.05083856, 0.04355096, 0.1139377, 
    0.2542818, 0.08082104, 0.04931356, 0.05280299, 0.004042157, 9.444714e-06, 
    0.04393785, 0.05553798, 0.09428339, 0.05995006, 0.01355529,
  2.18073e-07, 0.0008556654, 0.2238076, 0.09112708, 0.02740977, 0.07530124, 
    0.01884438, 0.002160602, 0.0002611716, 0.0004037477, 0.02644383, 
    0.002962813, 0.0006867496, 0.006665501, 0.03744622, 0.09010632, 
    0.06880378, 0.1098589, 0.05353689, 0.000163524, 2.845133e-06, 
    5.012404e-09, 0, 0.009270162, 0.0241031, 0.1257567, 0.09312513, 
    0.0113853, -1.998393e-05,
  -2.378575e-06, 0.002135565, 0.1350259, 0.02989442, 0.04532125, 0.08431175, 
    0.1014689, 0.05626266, 0.03812918, 0.00378145, 0.001353331, 0.001280874, 
    0.004162592, 0.05545568, 0.03312907, 0.05366345, 0.02200722, 
    0.0003721878, 5.331315e-08, 3.645897e-09, 0, 0, 4.445222e-06, 0.08901915, 
    0.1285973, 0.1667492, 0.05726643, 1.641115e-05, 2.256327e-08,
  0.03700088, 0.04599882, 0.1715252, 0.01138256, 0.0117362, 0.03256196, 
    0.009652364, 0.005849361, 0.09112144, 0.134486, 0.02060429, 0.02059931, 
    0.01288444, 0.06414209, 0.03286644, 0.02076501, 0.01205428, 
    -1.988446e-06, 4.669716e-05, 2.02718e-05, -8.288207e-10, 4.758663e-08, 
    0.005715289, 0.1865234, 0.05274501, 0.07294282, 0.07419688, 0.0002207817, 
    2.113098e-05,
  0.002097499, 5.392262e-08, 1.121176e-05, -2.64164e-05, 0.002690817, 
    0.03394499, 0.01158204, 0.07205804, 0.08074912, 0.1914451, 0.09827526, 
    0.04383818, 0.1074826, 0.08412921, 0.03765184, 0.009571484, 0.04830602, 
    0.06016532, 0.02536098, 0.1067385, 0.1919102, 0.01956876, 0.01526857, 
    0.002566452, 0.005277253, 0.03894197, 0.04820976, 0.001035044, 
    -2.490527e-06,
  0.01356021, 7.536901e-07, -5.116319e-08, 6.404971e-05, 3.921316e-08, 
    0.01190076, 0.01782838, 0.00200059, 0.02338327, -0.0005826174, 
    0.08329008, 0.02902254, 0.00773044, 0.008872497, 1.483947e-06, 
    -3.138204e-05, -0.0003705906, 0.005216246, 0.009517098, 0.01563603, 
    0.04040566, 0.1396329, 0.05485806, 0.0142323, 0.008940045, 0.0324313, 
    0.006185832, 0.09255907, 0.03645656,
  0.01165153, 0.02500988, 0.03614122, 0.04727059, 0.03123073, 0.04894236, 
    0.05804256, 0.006346058, 0.05746963, 0.08641519, 0.03251634, 0.0780898, 
    0.1003834, 0.1082592, 0.09079016, 0.08049974, 0.08738311, 0.06500324, 
    0.0177031, 0.01045451, 0.01452735, 0.04092191, 0.09285463, 0.05779968, 
    0.07384694, 0.1148874, 0.04826722, 0.02448514, 0.1006665,
  0.07942171, 0.09037825, 0.113927, 0.2001185, 0.1291424, 0.1307736, 
    0.04822449, 0.1099904, 0.04665085, 0.02304873, 0.05614436, 0.09228729, 
    0.1166541, 0.155208, 0.1680385, 0.1749902, 0.2014032, 0.2173238, 
    0.1459451, 0.1440675, 0.1032447, 0.07851515, 0.1230285, 0.1189215, 
    0.1885502, 0.1258129, 0.2400707, 0.06744733, 0.05211085,
  0.1312951, 0.1731496, 0.2418687, 0.2658554, 0.2673583, 0.207429, 0.1132157, 
    0.005313971, 0.01698955, 0.02947789, 0.06807628, 0.03562759, 0.207409, 
    0.126574, 0.1094875, 0.1550922, 0.1672762, 0.2778428, 0.3014653, 
    0.2278179, 0.1278059, 0.1488526, 0.1760997, 0.1767554, 0.1861887, 
    0.166512, 0.1453717, 0.1594729, 0.1208932,
  0.1452247, 0.1201179, 0.1921678, 0.1715955, 0.2023265, 0.2421625, 
    0.2716133, 0.2820433, 0.1972069, 0.06280546, 0.01867388, -8.7522e-05, 
    0.002426538, 0.04421213, 0.1200818, 0.2541677, 0.1303349, 0.1057992, 
    0.1661894, 0.1230308, 0.1104778, 0.1098757, 0.08061863, 0.06289533, 
    0.1344509, 0.2098919, 0.214555, 0.232875, 0.1742895,
  0.04154954, 0.0296201, 0.0117146, 0.06562625, 0.08024773, 0.09285485, 
    0.1301647, 0.09399075, 0.06124532, 0.07618811, 0.04273145, 0.02401346, 
    0.06202535, 0.1520425, 0.2069435, 0.1644017, 0.1382783, 0.1399495, 
    0.1092037, 0.06228922, 0.02482711, 0.05973157, 0.08731141, 0.05112598, 
    0.05281749, 0.04105488, -0.001286988, 0.1072878, 0.06940623,
  0.03951793, 0.0265006, 0.0234765, 0.02578622, 0.03173189, 0.02659886, 
    0.02163896, -9.256261e-05, 0, 0, 0.0001861686, 0.02067542, 0.02590759, 
    0.03850329, 0.04967674, 0.05443295, 0.06050944, 0.04998093, 0.04774405, 
    0.02925885, 0.013108, 0.0003245925, 0.01046949, 0.008779921, 0.01558568, 
    0.0004872552, -0.001763862, 0.005624364, 0.05763792,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.223541e-05, -0.000119271, 
    0.0003422842, -0.0003578724, -2.020465e-06, 0, 0, 0, 0, 0.001235976, 
    0.03984405, 0.0729559, 0.02893964, 0.02932963, -0.002704331, 0,
  0.1324703, 0.1742687, 0.1532315, 0.1131804, 0.00542783, 0.006902281, 
    0.07624899, 0.004879528, 0.002734063, -0.0009566552, -0.0001393145, 
    -0.001217622, 0.02478591, 0.11428, 0.1504194, 0.1403484, 0.1654758, 
    0.1507604, 0.125124, 0.1064442, 0.1256178, 0.1569271, 0.1545497, 
    0.2383368, 0.1932912, 0.1945963, 0.1716172, 0.1529147, 0.1167966,
  0.1779768, 0.2144243, 0.1586847, 0.1921015, 0.2347091, 0.2421617, 
    0.2060324, 0.179053, 0.1416667, 0.1705479, 0.1443396, 0.1256849, 
    0.1510217, 0.1891408, 0.244964, 0.2255573, 0.1958607, 0.2049707, 
    0.1953105, 0.2148616, 0.2105459, 0.2159078, 0.2197576, 0.2450418, 
    0.1933991, 0.1241849, 0.1289624, 0.1422289, 0.1655175,
  0.1046685, 0.1379008, 0.1460406, 0.1759985, 0.1575324, 0.1279166, 
    0.1225105, 0.1306498, 0.1863393, 0.1796749, 0.1877142, 0.1685741, 
    0.2255497, 0.1724312, 0.1514351, 0.1047948, 0.1157724, 0.1144512, 
    0.1190758, 0.112545, 0.1370602, 0.09860523, 0.1296386, 0.1619174, 
    0.1342568, 0.1984699, 0.1761709, 0.1360985, 0.1184459,
  0.05255746, 0.05929041, 0.02229138, 0.07051422, 0.08764092, 0.109384, 
    0.1281034, 0.09046897, 0.08714887, 0.1190461, 0.1048365, 0.09065754, 
    0.04280718, 0.1151797, 0.07589108, 0.09106519, 0.07497303, 0.05436803, 
    0.04538336, 0.1306476, 0.1461203, 0.1512874, 0.1542742, 0.07395729, 
    0.1171884, 0.1310478, 0.1225389, 0.1628586, 0.1078512,
  2.232196e-05, 0.005637493, 0.02522583, 0.04369782, 0.04642972, 0.03368172, 
    0.02045344, 0.04137456, 0.05483498, 0.03093402, 0.05411028, 0.08139409, 
    0.03168326, 0.06441461, 0.03420211, 0.04313181, 0.03739496, 0.09811905, 
    0.21587, 0.064945, 0.03473517, 0.03833771, 0.005411182, 6.403421e-05, 
    0.05385573, 0.04845291, 0.1026129, 0.04145284, 0.001142212,
  1.805668e-07, 9.102543e-05, 0.1848136, 0.07496777, 0.02530277, 0.0771604, 
    0.03199073, 0.0003307887, 5.053815e-06, 0.0001256639, 0.01536847, 
    0.002411381, 0.0005283362, 0.004199108, 0.046069, 0.07595316, 0.05488799, 
    0.1087406, 0.04477889, 3.878978e-05, 9.647293e-07, 9.039347e-09, 
    -5.392557e-11, 0.004204397, 0.01965453, 0.1329166, 0.1071811, 0.01547403, 
    8.301608e-07,
  -1.383674e-05, 0.003042691, 0.1158661, 0.02974156, 0.0382688, 0.09115451, 
    0.1254221, 0.05467262, 0.02859318, 0.005732756, 0.001419865, 0.001730266, 
    0.003979497, 0.0533162, 0.03323703, 0.05011392, 0.02512968, 0.0003568383, 
    1.521965e-05, 0, 0, 0, 5.026575e-06, 0.0633042, 0.1343231, 0.1536796, 
    0.04061579, -4.966633e-05, 1.20343e-07,
  0.05803273, 0.05699571, 0.1550587, 0.007167985, 0.01635393, 0.04499252, 
    0.006708399, 0.005244238, 0.09228798, 0.1363915, 0.01304243, 0.02172146, 
    0.009703211, 0.05511676, 0.02928525, 0.01853911, 0.001595646, 
    -2.892348e-06, 0.0001638373, 0.002756795, -1.173234e-07, 0.0003046859, 
    0.002276392, 0.1437428, 0.04842309, 0.09503431, 0.0787486, 0.0003319512, 
    -3.750481e-05,
  0.001276663, -4.084341e-06, 8.747901e-06, 3.091077e-05, 0.006556833, 
    0.03099515, 0.008061963, 0.07806141, 0.07991272, 0.1877092, 0.0882856, 
    0.0449171, 0.09218455, 0.07619039, 0.04527275, 0.007938392, 0.039278, 
    0.06422416, 0.02185952, 0.1458267, 0.1995274, 0.02759165, 0.01306405, 
    0.002016795, 0.00600969, 0.04195975, 0.04606375, 0.0020417, 3.077335e-05,
  0.006288652, -5.566972e-09, -8.288493e-09, 6.670118e-05, 2.535343e-07, 
    0.01380176, 0.008582558, 0.0007598608, 0.02669021, 0.0009673637, 
    0.08501533, 0.02957187, 0.006668879, 0.008463503, 6.656447e-08, 
    2.018472e-07, 0.0005392345, 0.003282519, 0.01267517, 0.01517649, 
    0.04078253, 0.149153, 0.04217653, 0.01054139, 0.006626225, 0.02977749, 
    0.001109453, 0.07083098, 0.06316166,
  0.01007505, 0.01362654, 0.02973447, 0.04558798, 0.02636198, 0.04739494, 
    0.04156554, 0.02433095, 0.086587, 0.08847835, 0.0356129, 0.0652329, 
    0.0970532, 0.09425327, 0.08305282, 0.08135147, 0.0706062, 0.06263637, 
    0.0122111, 0.02347943, 0.0127512, 0.02963607, 0.08402213, 0.06037917, 
    0.07696729, 0.1054201, 0.04048561, 0.01992579, 0.09471296,
  0.07202536, 0.08017694, 0.10658, 0.2206816, 0.103553, 0.1049861, 0.1003201, 
    0.1182622, 0.05711509, 0.0367513, 0.07732496, 0.1098563, 0.1235617, 
    0.1503137, 0.1809429, 0.1829313, 0.2143341, 0.2019707, 0.1475604, 
    0.1391025, 0.110372, 0.07915352, 0.09718556, 0.1051582, 0.1990869, 
    0.1105606, 0.2469544, 0.06343389, 0.06043739,
  0.1517268, 0.1682108, 0.2474031, 0.2564623, 0.2469337, 0.1873063, 
    0.1124678, 0.06131003, 0.04979257, 0.07478976, 0.1482299, 0.1048816, 
    0.2308347, 0.1373091, 0.140217, 0.1790418, 0.1865978, 0.2588833, 
    0.2696556, 0.2389228, 0.1350357, 0.1845261, 0.2394169, 0.2017652, 
    0.1912376, 0.1562706, 0.1299671, 0.1676813, 0.1243662,
  0.1437068, 0.1810934, 0.2699512, 0.2505594, 0.2695362, 0.2702385, 
    0.2865923, 0.2907977, 0.2359567, 0.1576894, 0.03749516, 0.02521694, 
    0.09692348, 0.1364391, 0.1758648, 0.2897691, 0.1628544, 0.1616767, 
    0.2342927, 0.1831124, 0.1554554, 0.192502, 0.1203775, 0.1564409, 
    0.248207, 0.2881061, 0.2720658, 0.2926416, 0.2137045,
  0.05911135, 0.09338034, 0.04814219, 0.1679319, 0.2090528, 0.1880769, 
    0.1829393, 0.1654514, 0.1592763, 0.1695441, 0.09228668, 0.1091923, 
    0.1954637, 0.2292531, 0.3260475, 0.1670945, 0.1398122, 0.2073715, 
    0.1746072, 0.08703911, 0.09346818, 0.1018859, 0.0964135, 0.06658576, 
    0.1192454, 0.07294542, 0.0192331, 0.1506469, 0.1081242,
  0.05666532, 0.0406189, 0.03057474, 0.05612914, 0.05983789, 0.06127835, 
    0.04122572, 0.001417899, -0.002388385, 0.03877436, 0.06258982, 
    0.06904197, 0.08605888, 0.08033703, 0.05816085, 0.06033567, 0.05582029, 
    0.05890491, 0.05967679, 0.07001489, 0.05046755, 0.02366719, 0.02081005, 
    0.01029752, 0.02707582, 0.005996521, -0.0007659078, 0.03865881, 0.1211673,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.051009e-05, 0.0101238, 0.01239053, 
    0.01781788, 0.03684637, 0.02546373, 0.005612647, -1.504531e-05, 
    -2.102657e-06, 0, 0.01678877, 0.2342471, 0.2192022, 0.1040272, 0.1060915, 
    0.02523354, 0,
  0.226203, 0.2303934, 0.1611543, 0.130047, 0.02927052, 0.02170956, 
    0.1520239, 0.01497428, 0.009017936, 0.002782491, 0.01112238, 0.01110623, 
    0.06727705, 0.1384896, 0.1634597, 0.15439, 0.1877013, 0.1780393, 
    0.1979734, 0.1763417, 0.2232888, 0.2586544, 0.3017022, 0.3761468, 
    0.237961, 0.2190536, 0.1991968, 0.2318166, 0.199505,
  0.2113589, 0.2202109, 0.1594277, 0.2079045, 0.2597619, 0.2542376, 
    0.2460483, 0.2111989, 0.1706458, 0.216393, 0.1892934, 0.1506989, 
    0.1568712, 0.2106969, 0.2571028, 0.2512118, 0.2007346, 0.2156852, 
    0.2097653, 0.2762245, 0.2159457, 0.2374707, 0.2280621, 0.2432305, 
    0.1857816, 0.1151689, 0.1366698, 0.173714, 0.2113669,
  0.1092879, 0.1313647, 0.1476579, 0.1720152, 0.1550409, 0.1180797, 
    0.1127087, 0.1382471, 0.1861201, 0.1723435, 0.1699801, 0.1631913, 
    0.2271096, 0.1618036, 0.1557622, 0.1060772, 0.1186788, 0.1114972, 
    0.1261325, 0.1251887, 0.1334935, 0.08645416, 0.1376394, 0.1662106, 
    0.1360415, 0.2066453, 0.1747287, 0.1335234, 0.1123108,
  0.06239489, 0.05119378, 0.01661824, 0.06477638, 0.09497903, 0.1070958, 
    0.128774, 0.08123567, 0.07698713, 0.1014633, 0.1053078, 0.08746249, 
    0.03803572, 0.1151072, 0.08343467, 0.0879704, 0.06877539, 0.05312078, 
    0.05107163, 0.1223668, 0.1514468, 0.1475252, 0.1915523, 0.06373134, 
    0.1152619, 0.1239267, 0.1186998, 0.1760492, 0.1112262,
  9.761762e-06, 0.00199335, 0.03019607, 0.03917311, 0.03227224, 0.02301764, 
    0.007319213, 0.03462585, 0.04488062, 0.01535032, 0.06915492, 0.09724185, 
    0.02812245, 0.05448503, 0.03691781, 0.03158342, 0.02652034, 0.08819345, 
    0.2118837, 0.05577613, 0.03082167, 0.04358438, 0.01156853, 0.001829017, 
    0.04605946, 0.05003069, 0.1090186, 0.04682919, 0.0006248073,
  2.623369e-07, 7.532917e-05, 0.1461981, 0.07845798, 0.03463051, 0.07789096, 
    0.03462338, 0.0001681441, 2.577832e-07, 6.600755e-05, 0.01337602, 
    0.005676845, 0.0004480231, 0.007644081, 0.03874507, 0.06411254, 
    0.0465516, 0.08804049, 0.03456702, 4.181448e-05, 2.640926e-07, 
    -7.421875e-10, -1.027836e-11, 0.003821696, 0.01972758, 0.1431334, 
    0.09964281, 0.01240669, -1.366431e-06,
  -3.961138e-05, 0.006363983, 0.1149302, 0.04406368, 0.03341241, 0.1014817, 
    0.1425526, 0.05061403, 0.02312755, 0.007626308, 0.001816733, 0.004341753, 
    0.003695644, 0.0476768, 0.0296548, 0.04128509, 0.0246549, 0.0007103064, 
    7.618312e-05, 0, 0, -1.057374e-10, 3.686656e-06, 0.04332873, 0.127164, 
    0.1507504, 0.01691045, 2.330216e-06, 3.431423e-07,
  0.1130773, 0.07181668, 0.1303641, 0.009812219, 0.009938062, 0.04850838, 
    0.005593674, 0.005201966, 0.09030349, 0.1355146, 0.01361183, 0.01399851, 
    0.008324763, 0.04792283, 0.02684864, 0.03009927, 0.006753075, 
    -1.11088e-05, 0.0004999891, -1.055341e-05, -5.288e-07, 5.499203e-05, 
    0.001372217, 0.125428, 0.05337711, 0.08565481, 0.08702172, 0.0006459769, 
    -0.0003131863,
  0.008520663, -5.125959e-05, -4.317189e-06, 2.997469e-06, 0.0103156, 
    0.02726076, 0.009858198, 0.07353495, 0.07659697, 0.1856036, 0.08086552, 
    0.03822472, 0.0841919, 0.07804763, 0.03439698, 0.01048762, 0.03168266, 
    0.0722062, 0.01855672, 0.17693, 0.1911925, 0.03365801, 0.0111072, 
    0.001790994, 0.006949979, 0.03652951, 0.04372701, 0.001146788, 
    0.0002277788,
  1.454511e-05, -4.102986e-07, -3.434675e-09, 2.977218e-05, 5.295375e-09, 
    0.01432865, 0.004272074, 0.0006937989, 0.05278868, 0.00113192, 
    0.09569073, 0.03851794, 0.005882973, 0.01185772, -3.887272e-06, 
    2.174257e-07, 0.0009408342, 0.0008951401, 0.009406781, 0.01764188, 
    0.04019557, 0.1629859, 0.03946988, 0.008429147, 0.008425059, 0.02763294, 
    0.0002096776, 0.06186153, 0.05490391,
  0.01187614, 0.006165484, 0.02276075, 0.03127957, 0.0207631, 0.04863993, 
    0.03298109, 0.04194965, 0.1290723, 0.1025245, 0.02702905, 0.05612588, 
    0.09378602, 0.08422131, 0.07363191, 0.06741629, 0.06385405, 0.04165063, 
    0.01142612, 0.01387598, 0.01007974, 0.02040159, 0.07240015, 0.05738372, 
    0.07409638, 0.07902823, 0.02443866, 0.01660178, 0.1015702,
  0.06752575, 0.08122916, 0.09741975, 0.2068447, 0.08699236, 0.07680702, 
    0.1395231, 0.1139042, 0.05062938, 0.045509, 0.08561022, 0.1305453, 
    0.1347465, 0.1620262, 0.1914943, 0.1874251, 0.2319757, 0.1778383, 
    0.138651, 0.1421551, 0.08830162, 0.07438279, 0.1000681, 0.09056801, 
    0.2094539, 0.09656664, 0.2061019, 0.05672896, 0.04416891,
  0.1444565, 0.1714762, 0.2229252, 0.2340435, 0.216615, 0.1526378, 0.1008433, 
    0.0955663, 0.1231459, 0.1349894, 0.176314, 0.1762478, 0.2310586, 
    0.1981626, 0.1750965, 0.1861045, 0.2094601, 0.2426233, 0.2496712, 
    0.2446603, 0.1381474, 0.2063441, 0.2415453, 0.2238449, 0.1992186, 
    0.1357018, 0.1264419, 0.1779223, 0.1102911,
  0.1373932, 0.2653837, 0.2673187, 0.2572351, 0.2992722, 0.2823632, 
    0.2706877, 0.3117177, 0.2774757, 0.1655797, 0.1043775, 0.1901519, 
    0.1402597, 0.1299687, 0.1756536, 0.2857141, 0.1724402, 0.1846534, 
    0.2907021, 0.1926821, 0.1897784, 0.2965796, 0.1472957, 0.2046853, 
    0.3333683, 0.4204654, 0.2863922, 0.2894563, 0.23632,
  0.08355992, 0.1218259, 0.1592943, 0.313796, 0.3734655, 0.3685536, 
    0.3328706, 0.3382874, 0.2452287, 0.2371703, 0.1565689, 0.2602374, 
    0.2580145, 0.2632511, 0.345705, 0.1750382, 0.1253705, 0.1722049, 
    0.1956725, 0.173524, 0.1294422, 0.1625723, 0.1733651, 0.1047984, 
    0.2215216, 0.09000333, 0.08152441, 0.1770818, 0.1300901,
  0.1768636, 0.1189324, 0.07410198, 0.102509, 0.1417982, 0.1673879, 
    0.1377015, 0.05425384, 0.08764475, 0.1242575, 0.0977796, 0.1059175, 
    0.1396781, 0.1582427, 0.1661461, 0.1441738, 0.0941965, 0.1234799, 
    0.150287, 0.1286545, 0.08230115, 0.08654632, 0.1048833, 0.03263446, 
    0.05168322, 0.01237803, 0.01998065, 0.08528213, 0.1719871,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.012848e-05, 0.05923627, 0.05422629, 
    0.08671772, 0.1635731, 0.1701253, 0.06311984, 0.0269693, 0.003453705, 
    -0.0008838758, 0.07597828, 0.277349, 0.2448048, 0.150471, 0.1865713, 
    0.1016468, 0.004730424,
  0.2472845, 0.2565383, 0.2115071, 0.2486607, 0.07752275, 0.06409384, 
    0.1871533, 0.03411108, 0.01064573, 0.02064744, 0.0215741, 0.03840102, 
    0.1133278, 0.2065166, 0.2211014, 0.1928014, 0.2204735, 0.255901, 
    0.2496265, 0.2215059, 0.2490629, 0.2823131, 0.3071935, 0.4723425, 
    0.2649499, 0.2193131, 0.1877688, 0.2398867, 0.2519954,
  0.2144936, 0.2422012, 0.1737132, 0.1945458, 0.2340796, 0.2501823, 
    0.2635416, 0.2203002, 0.1992398, 0.2317289, 0.1890674, 0.1711134, 
    0.1632159, 0.209289, 0.2441071, 0.236432, 0.2300274, 0.2437956, 
    0.2197608, 0.3157081, 0.2231391, 0.2549271, 0.2365208, 0.2309558, 
    0.1795628, 0.1086958, 0.1397435, 0.1674119, 0.2074527,
  0.09407219, 0.1305564, 0.1573787, 0.1683342, 0.1538658, 0.1147326, 
    0.1153582, 0.1431433, 0.1965018, 0.185362, 0.1597394, 0.1520234, 
    0.2277233, 0.1915627, 0.1652326, 0.1095192, 0.113104, 0.1189297, 
    0.1289131, 0.1148936, 0.1175106, 0.08560674, 0.1359517, 0.1530979, 
    0.1109625, 0.2122654, 0.1838342, 0.1388464, 0.1036808,
  0.07642827, 0.06652138, 0.01682192, 0.06267659, 0.08217755, 0.1056304, 
    0.1239616, 0.07557134, 0.07561199, 0.07225247, 0.09959929, 0.08795971, 
    0.05361812, 0.1347845, 0.08695558, 0.07206276, 0.05428358, 0.05762224, 
    0.05119117, 0.1251356, 0.1346748, 0.1279824, 0.1589468, 0.05230546, 
    0.1181824, 0.1134827, 0.1071325, 0.1781514, 0.1218276,
  -3.503249e-06, 0.0002313064, 0.05074716, 0.04315241, 0.02453375, 
    0.02045457, 0.005443489, 0.02727404, 0.03585156, 0.01013743, 0.07318032, 
    0.06070641, 0.02198279, 0.05687002, 0.04538262, 0.03900047, 0.02212789, 
    0.08179145, 0.2095786, 0.04847851, 0.03018165, 0.04071275, 0.01847709, 
    0.0008675134, 0.040818, 0.05323035, 0.1170042, 0.05125774, 0.002922454,
  8.95936e-07, 0.001174352, 0.1154345, 0.07200227, 0.03790502, 0.07639331, 
    0.02356532, 0.0002861028, 4.893989e-08, 2.158635e-05, 0.05933066, 
    0.01021005, 0.0005834966, 0.009204041, 0.0421047, 0.05851376, 0.03788589, 
    0.07378034, 0.02940371, 0.0002840238, 6.019736e-08, 1.326095e-09, 
    -2.63292e-09, 0.003020971, 0.02501965, 0.1621113, 0.1205146, 0.005153507, 
    1.693003e-06,
  0.00104982, 0.02030806, 0.09654599, 0.04951914, 0.03079421, 0.1016021, 
    0.143947, 0.04387392, 0.0143433, 0.006815376, 0.001694629, 0.002783624, 
    0.004638077, 0.0474229, 0.03546057, 0.04142385, 0.03389673, 0.001407198, 
    0.0003840466, 3.674699e-10, 3.956091e-10, 1.248218e-08, 6.211386e-06, 
    0.05085719, 0.1556067, 0.1582786, 0.02633244, 1.096562e-06, 3.459322e-05,
  0.1950474, 0.09513779, 0.1170237, 0.01524716, 0.007561954, 0.05163351, 
    0.004425863, 0.00360744, 0.1234259, 0.1523642, 0.01505923, 0.01116959, 
    0.009398855, 0.04146451, 0.02697925, 0.0232247, 0.01025541, 0.0003437088, 
    0.0002060659, -1.03589e-05, -2.716051e-05, 1.410237e-06, 0.003185791, 
    0.1179574, 0.06272813, 0.07313016, 0.1112198, 0.002098008, 0.01908616,
  0.02461913, -2.464333e-05, -2.951248e-06, -3.53106e-06, 0.0108565, 
    0.03443523, 0.01096179, 0.07162471, 0.08289792, 0.1872354, 0.1095567, 
    0.03480895, 0.08291882, 0.0884185, 0.04486197, 0.02207607, 0.02980118, 
    0.0819662, 0.02055638, 0.1811024, 0.196978, 0.03730297, 0.01107253, 
    0.002239982, 0.008287565, 0.02221073, 0.03974217, 0.001439647, 
    0.0003075153,
  2.240369e-06, -1.277664e-05, -5.902562e-09, 4.488554e-05, -7.345255e-09, 
    0.01661978, 0.00284191, 0.0005547185, 0.06175505, 0.007043663, 0.1084438, 
    0.0511552, 0.004561904, 0.01358513, -1.020298e-05, 1.391569e-07, 
    0.004184504, 0.0001351882, 0.006110168, 0.01799087, 0.02539804, 
    0.1754972, 0.03492094, 0.007236229, 0.01345288, 0.03277851, 6.318666e-05, 
    0.06478325, 0.05794906,
  0.009691676, 0.003906102, 0.01684999, 0.009637362, 0.02709374, 0.0505449, 
    0.02870889, 0.09174412, 0.1529283, 0.1050806, 0.01973085, 0.04680525, 
    0.08949788, 0.08035406, 0.05005234, 0.06051446, 0.06321699, 0.03319254, 
    0.01794124, 0.00636644, 0.008450952, 0.01274565, 0.06831139, 0.05504866, 
    0.06010081, 0.07560157, 0.01791152, 0.02595006, 0.1007637,
  0.06213272, 0.08243447, 0.1066815, 0.2038099, 0.07267239, 0.05868222, 
    0.1340303, 0.1021787, 0.04422953, 0.04940337, 0.09260426, 0.1373942, 
    0.1474494, 0.167883, 0.1795778, 0.18123, 0.2161676, 0.1792019, 0.1303845, 
    0.13351, 0.07242002, 0.06150926, 0.09248272, 0.09564549, 0.2125858, 
    0.07917017, 0.2052965, 0.04589279, 0.05584009,
  0.141419, 0.1707307, 0.2059427, 0.2226742, 0.198493, 0.151012, 0.08919806, 
    0.1067719, 0.1437922, 0.1575878, 0.1784908, 0.2251275, 0.2106967, 
    0.1965964, 0.1694164, 0.2041554, 0.2213987, 0.2400613, 0.2442026, 
    0.2494804, 0.1414203, 0.2238915, 0.2612776, 0.246669, 0.2111198, 
    0.1415709, 0.1169486, 0.1650094, 0.09599619,
  0.1515855, 0.2746287, 0.2481685, 0.278628, 0.3205705, 0.2919601, 0.2542982, 
    0.3120256, 0.3344569, 0.1973189, 0.1994788, 0.2454402, 0.163872, 
    0.1220768, 0.1691849, 0.2701986, 0.1790367, 0.2009593, 0.2830618, 
    0.2436363, 0.2000048, 0.3410144, 0.2244035, 0.2643104, 0.3895071, 
    0.442012, 0.2887582, 0.2789316, 0.2317089,
  0.09082569, 0.1269139, 0.1717953, 0.3391674, 0.4515826, 0.4031577, 
    0.3839954, 0.4361472, 0.3608612, 0.2789254, 0.1825805, 0.2888822, 
    0.2689912, 0.2554941, 0.338211, 0.171079, 0.1184803, 0.1624504, 
    0.2328199, 0.1884417, 0.1247319, 0.2302522, 0.2102426, 0.1826372, 
    0.2196066, 0.1372319, 0.1314108, 0.189742, 0.119843,
  0.2287972, 0.2685206, 0.1769208, 0.1155195, 0.1313139, 0.2150546, 
    0.1520457, 0.07063299, 0.1302324, 0.1538754, 0.1442687, 0.1742167, 
    0.218642, 0.2626193, 0.2809497, 0.1618299, 0.1528883, 0.1341535, 
    0.1909899, 0.1977913, 0.1423978, 0.1198059, 0.1322405, 0.06349885, 
    0.08220926, 0.01176178, 0.0263006, 0.0999348, 0.1806786,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  -0.005807792, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001376122, 0.1243018, 
    0.0598544, 0.07737783, 0.1592696, 0.2535512, 0.1748568, 0.07839314, 
    0.03731889, 0.02116097, 0.2307707, 0.2780789, 0.2206713, 0.1470736, 
    0.1840414, 0.2042692, 0.04626048,
  0.2119544, 0.2607968, 0.2080946, 0.3047245, 0.1342201, 0.1225803, 
    0.2213268, 0.08326457, 0.01511346, 0.09019931, 0.08550141, 0.07481556, 
    0.1847972, 0.2269723, 0.2357429, 0.2119036, 0.2385763, 0.2815973, 
    0.2938274, 0.2524769, 0.2369343, 0.2940969, 0.327238, 0.5036107, 
    0.2679534, 0.2180566, 0.1890075, 0.2514431, 0.2416277,
  0.2133574, 0.2344695, 0.1556953, 0.1942468, 0.223722, 0.2660779, 0.279957, 
    0.2464261, 0.21441, 0.2509866, 0.1707484, 0.1792266, 0.1676637, 
    0.2075545, 0.2325601, 0.2299006, 0.2185543, 0.225144, 0.2190714, 
    0.305233, 0.2290792, 0.2715367, 0.2434661, 0.2174595, 0.1468897, 
    0.09855759, 0.129324, 0.1653362, 0.1987837,
  0.09675586, 0.1303878, 0.1620038, 0.1568139, 0.1359396, 0.1181992, 
    0.1209326, 0.1336569, 0.1727686, 0.1778701, 0.1428298, 0.1557394, 
    0.2397519, 0.177751, 0.1563471, 0.110298, 0.1115848, 0.1084725, 
    0.1265988, 0.1131278, 0.1209095, 0.08418882, 0.1372631, 0.1424034, 
    0.1108166, 0.2158858, 0.1532814, 0.1480894, 0.1257194,
  0.09102619, 0.06523391, 0.0156764, 0.06541094, 0.07408289, 0.09695695, 
    0.117496, 0.07304979, 0.06852534, 0.06670517, 0.1035005, 0.06981196, 
    0.06290483, 0.1287345, 0.08995408, 0.07182214, 0.05954535, 0.07224569, 
    0.04679596, 0.1190294, 0.1151836, 0.1369963, 0.1928864, 0.03817254, 
    0.1035405, 0.1033343, 0.1136547, 0.176561, 0.1148713,
  -1.429884e-06, 4.268879e-05, 0.0659663, 0.05214022, 0.01910517, 0.027604, 
    0.001970578, 0.02440557, 0.02136237, 0.01007899, 0.03963097, 0.02405584, 
    0.02991282, 0.06561318, 0.0425048, 0.03466265, 0.03250343, 0.09833899, 
    0.2244144, 0.04213067, 0.03040907, 0.0341671, 0.0201098, -9.288724e-05, 
    0.04647639, 0.0552639, 0.1225998, 0.0668614, 0.002948638,
  2.118398e-06, 0.01903483, 0.1120313, 0.0631977, 0.04526466, 0.1013565, 
    0.01654648, 0.0004526385, 9.763872e-05, 0.0002839626, 0.1133969, 
    0.02841422, 0.003504251, 0.01145886, 0.04254904, 0.05200086, 0.03365692, 
    0.07762886, 0.02948478, 0.001026936, 5.739945e-07, 7.130512e-08, 
    2.345766e-08, 0.002568387, 0.03457021, 0.181346, 0.1099437, 0.003168018, 
    4.480862e-06,
  0.0006569417, 0.0377487, 0.1030699, 0.05468837, 0.0291955, 0.1271023, 
    0.1751172, 0.0495964, 0.01277927, 0.005526908, 0.001767051, 0.01590114, 
    0.006227599, 0.05982535, 0.05760521, 0.03785634, 0.03704308, 0.001958867, 
    0.0002107301, 1.453122e-08, 9.815472e-09, 2.516123e-08, 4.255984e-05, 
    0.08124513, 0.2045075, 0.1677974, 0.01623796, 1.026595e-06, 0.0009595411,
  0.2833691, 0.1394913, 0.1396657, 0.02359991, 0.006737711, 0.05543862, 
    0.005460786, 0.003531558, 0.1454664, 0.1626491, 0.02242964, 0.01665101, 
    0.01477257, 0.04922833, 0.02602826, 0.01491769, 0.01582422, 0.01247453, 
    0.0001642725, -7.078196e-05, 0.0004931707, 4.600517e-07, 0.005245547, 
    0.1391239, 0.09662735, 0.07454841, 0.1080502, 0.003359033, 0.07798306,
  0.003230923, 8.946926e-07, 0.0003808718, 8.142045e-05, 0.01814301, 
    0.04890729, 0.01503572, 0.07939624, 0.09251547, 0.2052411, 0.1283788, 
    0.04372827, 0.09375655, 0.107747, 0.06360967, 0.02748751, 0.03264327, 
    0.08585635, 0.02117023, 0.1730563, 0.2011078, 0.0529885, 0.01128029, 
    0.002759546, 0.008736161, 0.01291593, 0.04219637, 0.0007631464, 
    0.0004773969,
  8.290413e-06, -2.680603e-05, 3.52016e-08, 5.831574e-05, 3.919832e-09, 
    0.01619802, 0.003635308, 0.001833296, 0.04975707, 0.04811065, 0.1569049, 
    0.05616121, 0.008705677, 0.01271645, -1.962566e-05, 8.145436e-07, 
    0.007453855, 0.0001431646, 0.001810071, 0.01982736, 0.02250457, 
    0.1855284, 0.03446703, 0.009448458, 0.01809409, 0.03787912, 0.001876376, 
    0.06415254, 0.0333284,
  0.004623617, 0.002103116, 0.01095247, 0.001929626, 0.03570994, 0.0541721, 
    0.03704726, 0.1175078, 0.1530684, 0.1012745, 0.01402231, 0.04544677, 
    0.08629221, 0.08395082, 0.05632498, 0.05187489, 0.06434674, 0.04997348, 
    0.02085948, 0.02271698, 0.006480039, 0.009827166, 0.06196636, 0.05942282, 
    0.04677134, 0.06746802, 0.01739793, 0.02992305, 0.09080146,
  0.05658352, 0.08949275, 0.1105299, 0.2052497, 0.06842566, 0.04162069, 
    0.125426, 0.08644429, 0.03873425, 0.04784219, 0.095544, 0.1395112, 
    0.1434048, 0.1708676, 0.1650288, 0.1711294, 0.23552, 0.1827933, 
    0.1115039, 0.1230434, 0.05694862, 0.04208196, 0.1039274, 0.0813202, 
    0.1899193, 0.0883997, 0.1864366, 0.04512528, 0.03384038,
  0.1525551, 0.1603467, 0.1992851, 0.2242729, 0.161881, 0.1330423, 
    0.08433408, 0.1102014, 0.1851964, 0.1668626, 0.1571337, 0.210745, 
    0.2050427, 0.2067494, 0.1772931, 0.2143054, 0.2221305, 0.2256191, 
    0.2290901, 0.2435581, 0.1832011, 0.2182475, 0.2648925, 0.2702963, 
    0.2398351, 0.1338635, 0.1162736, 0.1527596, 0.1352438,
  0.1797916, 0.3236171, 0.2367783, 0.3012711, 0.2977606, 0.2953922, 
    0.2435236, 0.3278188, 0.3518808, 0.1992427, 0.239194, 0.2533986, 
    0.1448664, 0.1141682, 0.1812635, 0.2639101, 0.1911051, 0.233061, 
    0.2835811, 0.2638898, 0.1977673, 0.359364, 0.3137884, 0.369881, 
    0.4079836, 0.4715373, 0.3072571, 0.2960941, 0.2631697,
  0.0808105, 0.1648626, 0.2229287, 0.3479874, 0.4915915, 0.4076762, 
    0.4015222, 0.4379451, 0.3957414, 0.2830915, 0.2059875, 0.2883437, 
    0.2674807, 0.2516437, 0.3011944, 0.1628108, 0.09046312, 0.1564531, 
    0.2151073, 0.1804839, 0.1292904, 0.2785038, 0.2761932, 0.2314173, 
    0.2202895, 0.2458546, 0.1875977, 0.1962847, 0.1196327,
  0.2189586, 0.2555628, 0.1992095, 0.0758026, 0.07838713, 0.1813624, 
    0.0926056, 0.04499929, 0.1176898, 0.1553945, 0.1602877, 0.2037369, 
    0.2691494, 0.2606087, 0.2907005, 0.1915665, 0.1783377, 0.1572906, 
    0.1916689, 0.2279793, 0.148382, 0.1240097, 0.1098316, 0.05939413, 
    0.0917026, 0.0315998, 0.02574947, 0.08122953, 0.2109991,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0.04682167, -0.001002102, -1.067726e-05, 0, 0, -9.228343e-06, 0, 0, 0, 0, 
    0, 0, 0.001045502, 0.136447, 0.05876502, 0.06379818, 0.1481079, 
    0.2250102, 0.230802, 0.1797196, 0.1752621, 0.1383318, 0.4354391, 
    0.2714962, 0.2040983, 0.1348781, 0.1783961, 0.2172524, 0.09074817,
  0.1999771, 0.281306, 0.1996977, 0.3246719, 0.1774507, 0.2037148, 0.2267869, 
    0.1296444, 0.05180496, 0.1787736, 0.149441, 0.0944429, 0.228517, 
    0.2238831, 0.2370637, 0.2178183, 0.2608651, 0.2895584, 0.3173545, 
    0.2619422, 0.2416047, 0.3154548, 0.3255976, 0.5123252, 0.2742258, 
    0.2152713, 0.2032056, 0.2595035, 0.2499512,
  0.2138312, 0.2293121, 0.156233, 0.193192, 0.2345917, 0.2660813, 0.280505, 
    0.2856807, 0.2386232, 0.2588772, 0.1698189, 0.1715673, 0.180743, 
    0.2030936, 0.2480481, 0.242578, 0.2304453, 0.2399388, 0.2293243, 
    0.3244029, 0.2650199, 0.246245, 0.2302133, 0.2159626, 0.1436164, 
    0.09730545, 0.1094444, 0.1681794, 0.211275,
  0.09338535, 0.1168801, 0.159307, 0.1588954, 0.1251381, 0.1187534, 
    0.1065206, 0.1487496, 0.1844079, 0.1849734, 0.152226, 0.1520186, 
    0.2674559, 0.1874223, 0.1517609, 0.1074798, 0.1094977, 0.1108728, 
    0.1176103, 0.104171, 0.123577, 0.1083833, 0.1458679, 0.1448641, 
    0.1194525, 0.246892, 0.178903, 0.1301766, 0.1079508,
  0.09533449, 0.06678421, 0.02050965, 0.06375083, 0.07807551, 0.093047, 
    0.122931, 0.09579629, 0.06606827, 0.06801631, 0.0995057, 0.06258789, 
    0.07633228, 0.1197534, 0.1068675, 0.07093886, 0.05432466, 0.06853648, 
    0.05117891, 0.1111529, 0.09637018, 0.1274558, 0.1630795, 0.0310234, 
    0.1060311, 0.1069926, 0.1123097, 0.1643421, 0.1230684,
  0.0002039637, 0.0003964456, 0.06845185, 0.06229116, 0.01894366, 0.02952591, 
    0.005182787, 0.02836027, 0.02537347, 0.009837659, 0.03020115, 0.00414172, 
    0.03715484, 0.07305767, 0.04920938, 0.04764127, 0.02608504, 0.116205, 
    0.24503, 0.05871457, 0.05045878, 0.02279416, 0.0152644, -7.381525e-06, 
    0.08030785, 0.06289007, 0.1527868, 0.06425864, 0.001903748,
  3.288073e-06, 0.01558997, 0.1161925, 0.0578923, 0.06622002, 0.1163669, 
    0.01369527, 0.001007703, 0.001495945, 0.001447564, 0.1059487, 0.05675904, 
    0.005623613, 0.01570066, 0.05010796, 0.04986731, 0.02948324, 0.08557129, 
    0.0335881, 0.002808919, 5.610923e-07, 1.087219e-07, 3.946517e-08, 
    0.0008018837, 0.04791902, 0.203874, 0.07929415, 0.001697569, -1.735959e-05,
  0.00302611, 0.04306173, 0.1378783, 0.06533793, 0.03286638, 0.1488287, 
    0.1979112, 0.05746878, 0.01480178, 0.004717238, 0.001425425, 0.02095679, 
    0.007132404, 0.07841203, 0.06447534, 0.04618674, 0.03584255, 0.002933695, 
    0.0001108024, 3.111855e-08, 1.952596e-08, 1.730808e-08, 0.0001836765, 
    0.1168726, 0.2376854, 0.2003133, 0.009194703, 4.168755e-07, 9.69691e-06,
  0.2566376, 0.1978342, 0.1784527, 0.03774649, 0.005358019, 0.06473415, 
    0.004361329, 0.003675165, 0.1890265, 0.1986039, 0.03024306, 0.02058754, 
    0.01420341, 0.05101654, 0.02763071, 0.02033691, 0.01614694, 0.009444749, 
    -0.000109887, -3.363717e-06, 0.002330007, -8.666153e-05, 0.01034006, 
    0.1867927, 0.1440974, 0.06472839, 0.1148523, 0.005780385, 0.04790483,
  0.0002042658, 3.238926e-06, 0.00318313, 0.003141303, 0.04488477, 
    0.05887592, 0.03978325, 0.08414355, 0.1044705, 0.2167255, 0.1382903, 
    0.0538729, 0.1098915, 0.1215848, 0.08331801, 0.02872534, 0.04373452, 
    0.08669958, 0.02501208, 0.1690943, 0.224366, 0.05389811, 0.01007905, 
    0.003405564, 0.009315267, 0.0112702, 0.03360134, 0.00148883, 0.001050056,
  1.763049e-05, 1.864554e-06, 1.067943e-07, 4.797359e-05, -1.424863e-07, 
    0.01863309, 0.01177933, 0.006306862, 0.03953303, 0.06765933, 0.1941623, 
    0.06193535, 0.01273865, 0.01146986, -4.345581e-05, 2.997891e-06, 
    0.02648133, 0.001530182, 0.01228858, 0.001772209, 0.01425332, 0.1907521, 
    0.04095091, 0.01281356, 0.02163604, 0.04839312, 0.00928867, 0.06941474, 
    0.006424393,
  0.0008168304, 0.002372889, 0.005821939, 0.0009914704, 0.03925864, 
    0.05640268, 0.03158258, 0.129424, 0.1600409, 0.1010209, 0.01781013, 
    0.04824971, 0.08987432, 0.08447972, 0.06541783, 0.05651322, 0.06380812, 
    0.05902585, 0.01788781, 0.004840775, 0.006408575, 0.00395982, 0.05885251, 
    0.06450562, 0.04207343, 0.08593579, 0.02483155, 0.04795671, 0.06488582,
  0.05222664, 0.08941947, 0.1099052, 0.2116054, 0.06800445, 0.02915195, 
    0.1169276, 0.0754616, 0.03014449, 0.04104641, 0.110412, 0.1407321, 
    0.1426962, 0.1742135, 0.1587142, 0.1724767, 0.2250602, 0.1896643, 
    0.09072106, 0.11815, 0.04650486, 0.02975168, 0.09722012, 0.0883226, 
    0.1891723, 0.07831945, 0.1804799, 0.0330263, 0.03637787,
  0.1271477, 0.1656191, 0.2131286, 0.2180501, 0.1608379, 0.1258615, 
    0.0861406, 0.1207466, 0.1673366, 0.182706, 0.1420572, 0.1960759, 
    0.2118583, 0.2148674, 0.1862413, 0.2124528, 0.2322118, 0.2480613, 
    0.2232101, 0.2332069, 0.1815889, 0.2132946, 0.2514871, 0.2809524, 
    0.2468356, 0.1522208, 0.1182433, 0.1627793, 0.127629,
  0.1967896, 0.3485883, 0.2601541, 0.3632646, 0.2968115, 0.2825493, 
    0.2155027, 0.3258179, 0.3556808, 0.1962548, 0.2527124, 0.207932, 
    0.1280014, 0.09644178, 0.1921551, 0.282189, 0.1881987, 0.2344227, 
    0.3246209, 0.2899221, 0.2043461, 0.3745015, 0.2942257, 0.3776501, 
    0.4167823, 0.4807715, 0.3138253, 0.2940805, 0.2809941,
  0.106006, 0.1736628, 0.2107874, 0.3721518, 0.4955387, 0.4242758, 0.3984829, 
    0.4304075, 0.4129878, 0.2685807, 0.2161464, 0.2852505, 0.2661042, 
    0.2563875, 0.2731225, 0.1365392, 0.06685966, 0.1290593, 0.2303484, 
    0.1408555, 0.1254795, 0.3227779, 0.2693158, 0.2451328, 0.2091576, 
    0.3021396, 0.233753, 0.1776381, 0.1366072,
  0.1670657, 0.2149826, 0.1280814, 0.06107707, 0.0716198, 0.1468842, 
    0.07356048, 0.04046048, 0.118473, 0.1598672, 0.1574735, 0.1784595, 
    0.2477173, 0.2880518, 0.292973, 0.2134946, 0.2065704, 0.1523857, 
    0.169799, 0.2200847, 0.1459453, 0.1056828, 0.1137953, 0.06773885, 
    0.08660889, 0.02243353, 0.04522412, 0.06121626, 0.1845028,
  0.002258079, 0.001228736, 0.000199392, -0.0008299515, -0.001859295, 
    -0.002888639, -0.003917982, 0, 0, 0, 0, 0, 0, 0, -0.003436236, 
    -0.002345367, -0.001254499, -0.0001636303, 0.0009272383, 0.002018107, 
    0.003108975, -0.004828497, -0.004890022, -0.004951547, -0.005013072, 
    -0.005074597, -0.005136122, -0.005197647, 0.003081554,
  0.1150018, 0.01118559, 0.01310859, 0.000617214, -0.0002069959, 
    -0.0005898736, 4.995768e-06, 0, 0, 0, -1.892861e-06, 0.0004157126, 
    0.0201257, 0.1365886, 0.04416201, 0.04169358, 0.1449379, 0.1971026, 
    0.2141887, 0.1791275, 0.2721501, 0.3650193, 0.4235972, 0.260433, 0.18099, 
    0.1320685, 0.1674028, 0.2207998, 0.1275752,
  0.2149268, 0.2692688, 0.1944939, 0.3384354, 0.2670592, 0.2601397, 
    0.2228925, 0.1627787, 0.1016603, 0.2488099, 0.2221793, 0.1650718, 
    0.2490691, 0.234453, 0.2716413, 0.2238749, 0.2634302, 0.2935, 0.3125436, 
    0.2673657, 0.2609911, 0.338282, 0.2688003, 0.5245894, 0.268874, 
    0.2109336, 0.2086174, 0.310489, 0.268411,
  0.2493758, 0.2412658, 0.1762357, 0.2199994, 0.2597874, 0.2830327, 0.272085, 
    0.2922471, 0.2345144, 0.3003549, 0.1938114, 0.1808456, 0.1607285, 
    0.1940467, 0.2446584, 0.2512326, 0.2411625, 0.24001, 0.2271354, 
    0.3125669, 0.2835551, 0.2612248, 0.2391298, 0.2062575, 0.12957, 
    0.0755856, 0.09190002, 0.1794279, 0.2318494,
  0.1088004, 0.1144363, 0.1587935, 0.1790216, 0.1289203, 0.1338006, 
    0.1253612, 0.1533612, 0.1870607, 0.1645964, 0.1351872, 0.1656811, 
    0.2150294, 0.1697415, 0.1263361, 0.1036564, 0.1027217, 0.1145616, 
    0.1124653, 0.1059099, 0.1226914, 0.1081234, 0.1497896, 0.155606, 
    0.1264464, 0.2337762, 0.1358338, 0.1186827, 0.1057219,
  0.1093622, 0.07417666, 0.03737146, 0.07399275, 0.08545593, 0.09586331, 
    0.118568, 0.1022885, 0.05964997, 0.07063419, 0.0821883, 0.0560591, 
    0.07061113, 0.1276458, 0.1052419, 0.06456686, 0.04925431, 0.0697186, 
    0.05694807, 0.1243384, 0.09664018, 0.1181673, 0.1508749, 0.03042092, 
    0.09783704, 0.1059845, 0.1079927, 0.1466097, 0.1236703,
  0.00251039, 0.0007353298, 0.06002808, 0.0731856, 0.01971041, 0.03911002, 
    0.01026309, 0.03401814, 0.04347752, 0.01211263, 0.01407041, 0.0008056179, 
    0.04802566, 0.09464069, 0.06238077, 0.06490499, 0.03565215, 0.1180939, 
    0.2519109, 0.06571914, 0.0887102, 0.007108722, 0.009200673, 2.448326e-07, 
    0.09060715, 0.08118748, 0.1620882, 0.07041348, 7.442538e-05,
  2.424375e-06, 0.009036276, 0.1355338, 0.0558406, 0.06124816, 0.1185577, 
    0.006365966, 0.000914216, 1.617486e-05, 0.0008083488, 0.03945686, 
    0.03873643, 0.00418445, 0.01827352, 0.0530561, 0.05999075, 0.03131686, 
    0.08914872, 0.04730082, 0.00169724, 4.762489e-07, 1.682931e-07, 
    7.918116e-08, 0.000200771, 0.05227157, 0.2212411, 0.06664122, 
    -1.297763e-05, 1.075074e-05,
  5.887478e-05, 0.02869694, 0.1674383, 0.06400579, 0.03586197, 0.14746, 
    0.1566864, 0.06334298, 0.0142877, 0.006505647, 0.002959319, 0.008935454, 
    0.007927809, 0.06169514, 0.0626692, 0.05034306, 0.03389214, 0.006673787, 
    0.002144441, 4.323558e-08, 1.592793e-08, 5.090573e-08, 1.879375e-05, 
    0.1285125, 0.2280385, 0.2355355, 0.003088422, 2.019617e-07, -6.996838e-06,
  0.2598746, 0.2768129, 0.2093792, 0.05810486, 0.00792968, 0.06086442, 
    0.00552149, 0.003872799, 0.2206677, 0.2218782, 0.02529142, 0.01155539, 
    0.01095464, 0.04480557, 0.0240074, 0.02023802, 0.01399699, 0.001981446, 
    6.128251e-06, 9.886217e-06, 0.002421146, 0.008134305, 0.03618608, 
    0.2051704, 0.1672968, 0.06198215, 0.1243616, 0.007833875, 0.04352146,
  0.000155487, 1.092825e-05, 0.01098488, 0.01935377, 0.05638584, 0.05417253, 
    0.06292813, 0.07106715, 0.09033515, 0.1830829, 0.1273206, 0.04360082, 
    0.09799373, 0.09751125, 0.08533835, 0.03583001, 0.05907813, 0.0864507, 
    0.03407237, 0.153235, 0.207159, 0.05527218, 0.01110903, 0.004957204, 
    0.01688444, 0.01387435, 0.03294365, 0.003717438, 0.003158468,
  1.342701e-05, 1.531511e-06, 1.798363e-07, 5.736827e-05, -2.904886e-06, 
    0.02220596, 0.0198949, 0.005235357, 0.03781872, 0.09134739, 0.1968201, 
    0.04801526, 0.01170219, 0.01101302, -6.19062e-05, 7.57927e-06, 
    0.03309211, 0.00428435, 0.02386674, 0.0009788263, 0.01710458, 0.1872572, 
    0.04289006, 0.01687208, 0.02611369, 0.05484989, 0.01773139, 0.06590944, 
    0.0008761706,
  0.0001055488, 0.003434402, 0.004031392, 0.005397937, 0.04114128, 0.0677863, 
    0.03727354, 0.1503183, 0.1738679, 0.09971991, 0.01876982, 0.04239576, 
    0.0895938, 0.07908396, 0.07806306, 0.06654427, 0.06677079, 0.05783865, 
    0.01231185, 0.0002321603, 0.01062801, 0.001699885, 0.0584298, 0.06493602, 
    0.04354534, 0.08905438, 0.0354431, 0.05683595, 0.04373299,
  0.05048128, 0.08810167, 0.1173109, 0.2152079, 0.08138508, 0.02587929, 
    0.122981, 0.06488407, 0.02520562, 0.02594617, 0.1205805, 0.1396196, 
    0.1407849, 0.1695853, 0.1669368, 0.1612438, 0.208177, 0.1939642, 
    0.08199709, 0.1077146, 0.04781893, 0.01508974, 0.07502841, 0.09192671, 
    0.1861718, 0.08473797, 0.1662793, 0.03181672, 0.04961114,
  0.135623, 0.1902987, 0.2164242, 0.2076325, 0.1320075, 0.140446, 0.09012077, 
    0.1152715, 0.1472326, 0.1758431, 0.136951, 0.1913226, 0.2199645, 
    0.2407526, 0.2004324, 0.2166618, 0.2127939, 0.2414482, 0.2000363, 
    0.2375341, 0.171915, 0.2076944, 0.259305, 0.2898091, 0.267996, 0.156171, 
    0.1215824, 0.1787488, 0.1381612,
  0.2639281, 0.3893025, 0.3005594, 0.3462526, 0.2462002, 0.299555, 0.2356368, 
    0.3369452, 0.3549029, 0.2300431, 0.2575274, 0.1873974, 0.1178397, 
    0.08379129, 0.2354778, 0.2674178, 0.1780638, 0.3191588, 0.2999732, 
    0.2662702, 0.1983675, 0.424071, 0.3075922, 0.3293757, 0.4111793, 
    0.4776087, 0.3221669, 0.313963, 0.2806035,
  0.1339768, 0.1996643, 0.2503701, 0.3882041, 0.5081886, 0.4857143, 
    0.3542834, 0.4481574, 0.4422896, 0.2961277, 0.1965065, 0.300267, 
    0.2683766, 0.2464295, 0.2785922, 0.1216668, 0.04412363, 0.1283761, 
    0.2261693, 0.1487327, 0.1013999, 0.3501223, 0.2658912, 0.2444024, 
    0.1498195, 0.319509, 0.2977979, 0.2047965, 0.1928776,
  0.1438888, 0.178111, 0.0877572, 0.04942925, 0.08474731, 0.103325, 
    0.04669231, 0.03011525, 0.1116134, 0.1506058, 0.1586652, 0.245815, 
    0.3177605, 0.2923595, 0.3213282, 0.2605847, 0.1585018, 0.1524866, 
    0.1961884, 0.2375086, 0.1579322, 0.1088659, 0.08304308, 0.06647819, 
    0.07403915, 0.03746343, 0.05317342, 0.04816094, 0.1659452,
  0.08450992, 0.07685507, 0.06920023, 0.06154538, 0.05389053, 0.04623568, 
    0.03858084, 0.03566435, 0.03446647, 0.03326858, 0.0320707, 0.03087281, 
    0.02967492, 0.02847704, 0.0261016, 0.03476835, 0.0434351, 0.05210186, 
    0.06076861, 0.06943537, 0.07810212, 0.09715174, 0.09733772, 0.0975237, 
    0.09770968, 0.09789565, 0.09808163, 0.09826761, 0.0906338,
  0.1499721, 0.04051647, 0.01841679, 0.01617742, 0.007311963, 0.0003118131, 
    -2.00108e-05, -3.116575e-06, 0, 0, 0.004811373, 0.02658708, 0.05608157, 
    0.1317863, 0.02357394, 0.02286299, 0.1335853, 0.1747068, 0.1843554, 
    0.1758976, 0.2851612, 0.4932566, 0.4048173, 0.2468368, 0.1608488, 
    0.1323329, 0.1634384, 0.2222202, 0.1458171,
  0.2183622, 0.2420221, 0.1871201, 0.3476649, 0.3556248, 0.2739117, 
    0.2294963, 0.1865532, 0.1946235, 0.2674305, 0.2652759, 0.1737883, 
    0.265727, 0.2776479, 0.2772828, 0.2695393, 0.2999875, 0.3428089, 
    0.3227955, 0.2846608, 0.3082169, 0.3419658, 0.3165823, 0.5742831, 
    0.2539759, 0.2167476, 0.2728025, 0.3620413, 0.2637802,
  0.2419251, 0.2713962, 0.1654178, 0.2698061, 0.2904548, 0.3710948, 
    0.3179195, 0.3393489, 0.3220618, 0.3491381, 0.2405286, 0.2048686, 
    0.1622922, 0.2061483, 0.239775, 0.2488943, 0.2452636, 0.253577, 
    0.2465134, 0.3270195, 0.2914893, 0.2616928, 0.2310863, 0.1912206, 
    0.1340058, 0.1016718, 0.1044124, 0.1941482, 0.2372192,
  0.1084211, 0.1268145, 0.1781902, 0.1732013, 0.134198, 0.130216, 0.1244674, 
    0.1419761, 0.18198, 0.18278, 0.1466977, 0.1637116, 0.1832829, 0.155294, 
    0.1289913, 0.1149297, 0.1152221, 0.1211811, 0.1242937, 0.1184154, 
    0.112628, 0.121201, 0.168957, 0.168042, 0.1552308, 0.2279612, 0.153738, 
    0.1390091, 0.1145484,
  0.1246921, 0.07947037, 0.05737844, 0.09717724, 0.1032696, 0.09612899, 
    0.1222858, 0.1035051, 0.06395822, 0.0818584, 0.05401621, 0.03447982, 
    0.07088348, 0.137246, 0.09887457, 0.07547864, 0.05305012, 0.07010091, 
    0.05914536, 0.1307984, 0.1035746, 0.1223137, 0.1612579, 0.03682105, 
    0.08295465, 0.1156046, 0.1046887, 0.1522886, 0.1244897,
  0.004746923, 0.0007396901, 0.06270363, 0.08186664, 0.01828555, 0.0387, 
    0.01335421, 0.04127478, 0.05565673, 0.009683714, 0.005570503, 
    3.058043e-05, 0.04320359, 0.1212257, 0.08222148, 0.06612993, 0.05548512, 
    0.1258537, 0.2702879, 0.05238442, 0.1002306, 0.004034916, 0.01186628, 
    2.643272e-08, 0.04288289, 0.07553078, 0.144354, 0.07346187, 0.0007588746,
  1.206272e-06, 0.0004045317, 0.1360562, 0.03585356, 0.05578915, 0.1048781, 
    0.003082221, 0.001572775, 6.648598e-06, 9.691696e-05, 0.01022217, 
    0.009030983, 0.01395067, 0.01793021, 0.05988918, 0.05621582, 0.03182809, 
    0.09061143, 0.05186337, 0.0103436, 3.093129e-07, 1.833391e-07, 
    9.313752e-08, 1.711236e-05, 0.05189427, 0.2338354, 0.06092384, 
    -1.592234e-05, 6.921902e-06,
  -5.574379e-06, 0.009878762, 0.1485005, 0.05812164, 0.03947521, 0.142975, 
    0.1326509, 0.05579133, 0.01270601, 0.005573733, 0.003894384, 0.006866984, 
    0.006441937, 0.04955417, 0.06260935, 0.0491616, 0.036583, 0.01063507, 
    0.002965337, 5.291228e-08, 8.783428e-09, 6.195556e-08, 6.863266e-06, 
    0.08749288, 0.183489, 0.188813, 0.003059332, 1.681357e-07, -4.370996e-07,
  0.1881884, 0.2873304, 0.1508344, 0.0695218, 0.00795753, 0.06091049, 
    0.007661765, 0.00383048, 0.1961227, 0.2121542, 0.02433165, 0.009379805, 
    0.01070343, 0.03705172, 0.01855473, 0.01763028, 0.006271465, 
    2.132774e-05, 1.187299e-05, 4.908076e-06, 0.0007699293, 0.01020236, 
    0.04055331, 0.1490705, 0.1627866, 0.05405582, 0.1413717, 0.01754482, 
    0.04941315,
  4.307522e-05, 0.0001336466, 0.01308938, 0.1229591, 0.0716716, 0.04895018, 
    0.0777191, 0.06288871, 0.07670256, 0.1605327, 0.1192784, 0.03464158, 
    0.08243669, 0.08159497, 0.0885516, 0.04229651, 0.06352318, 0.07854852, 
    0.04500233, 0.150005, 0.1941443, 0.04605177, 0.02355525, 0.006280897, 
    0.01756811, 0.01145367, 0.02890214, 0.0007523923, 0.002100305,
  7.344171e-06, 6.547057e-07, 3.614686e-07, 1.817898e-05, 3.400711e-05, 
    0.02607, 0.03156745, 0.004449754, 0.04067802, 0.08745827, 0.1607658, 
    0.04407641, 0.01211128, 0.01198296, 6.224421e-06, 0.0002891074, 
    0.03642913, 0.002997692, 0.02676737, 0.0006108622, 0.01197909, 0.1966321, 
    0.0429311, 0.01881413, 0.02453936, 0.06050331, 0.01630335, 0.05521786, 
    2.998501e-05,
  -2.386963e-05, 0.006569932, 0.003705804, 0.01014133, 0.04159498, 
    0.05266779, 0.05521067, 0.1657607, 0.191848, 0.09591084, 0.01889841, 
    0.04543998, 0.08606102, 0.08496982, 0.09890708, 0.07240709, 0.07579201, 
    0.06017286, 0.01962054, 1.196628e-05, 0.01976158, 0.001637864, 
    0.06174346, 0.05514347, 0.04558175, 0.08808535, 0.04822999, 0.07016211, 
    0.02096201,
  0.04755593, 0.08759965, 0.1299101, 0.2248113, 0.07026611, 0.02374686, 
    0.1298746, 0.05561967, 0.01902174, 0.02072765, 0.1096036, 0.13463, 
    0.14894, 0.1689848, 0.1678305, 0.1553122, 0.2206367, 0.1897939, 
    0.08205152, 0.1051508, 0.04764117, 0.01308463, 0.06836821, 0.08911358, 
    0.189019, 0.1056116, 0.1775672, 0.03504482, 0.05295167,
  0.1389509, 0.2349033, 0.2134914, 0.1887037, 0.1288877, 0.1272554, 
    0.08321116, 0.1045096, 0.1403541, 0.1687603, 0.1312358, 0.1901939, 
    0.2437553, 0.2583089, 0.1949336, 0.2302462, 0.2066821, 0.2503641, 
    0.2077767, 0.2433988, 0.1892926, 0.2020235, 0.2733633, 0.2863143, 
    0.2316847, 0.150456, 0.1284598, 0.2019978, 0.1379886,
  0.2587414, 0.404697, 0.3246391, 0.3356045, 0.2285721, 0.2875266, 0.2165017, 
    0.3348001, 0.3584752, 0.257947, 0.2337744, 0.1398363, 0.1489833, 
    0.08324251, 0.23623, 0.2288275, 0.2069195, 0.3243597, 0.2930334, 
    0.3016157, 0.2459865, 0.4195898, 0.3764919, 0.3368164, 0.391383, 
    0.5210718, 0.3215233, 0.2969284, 0.2996864,
  0.1748793, 0.2481994, 0.285698, 0.4167968, 0.5743945, 0.531566, 0.4365415, 
    0.5437875, 0.461284, 0.3197688, 0.2121782, 0.2549274, 0.2661649, 
    0.265651, 0.2722096, 0.1188367, 0.0939761, 0.1639923, 0.2145275, 
    0.1751646, 0.1489397, 0.3963031, 0.3203963, 0.3370635, 0.146373, 
    0.339552, 0.3526372, 0.2111494, 0.1970428,
  0.1483313, 0.1925723, 0.1086521, 0.06299654, 0.08780296, 0.05627069, 
    0.03044059, 0.02458298, 0.1065999, 0.1434793, 0.1740351, 0.2423688, 
    0.3282336, 0.2917467, 0.3554199, 0.3060883, 0.2033811, 0.1674114, 
    0.2581647, 0.2298489, 0.1646372, 0.1596243, 0.08735353, 0.04459435, 
    0.0578513, 0.04488757, 0.04510431, 0.04935395, 0.1575373,
  0.1784922, 0.1723485, 0.1662048, 0.1600611, 0.1539174, 0.1477737, 
    0.1416301, 0.1535149, 0.1515606, 0.1496063, 0.147652, 0.1456977, 
    0.1437434, 0.1417891, 0.1281496, 0.1383034, 0.1484573, 0.1586111, 
    0.168765, 0.1789188, 0.1890727, 0.2026021, 0.2005463, 0.1984904, 
    0.1964346, 0.1943787, 0.1923228, 0.190267, 0.1834071,
  0.1824355, 0.07230795, 0.01855004, 0.02151709, 0.0196365, 0.01428925, 
    0.00571099, -0.0005908213, -2.724046e-05, 0.001260161, 0.06193144, 
    0.04788537, 0.116056, 0.1352767, 0.02197598, 0.007623529, 0.1105025, 
    0.1436072, 0.1771749, 0.1643015, 0.261862, 0.5191927, 0.4000694, 
    0.2627842, 0.1671714, 0.1199893, 0.1492395, 0.2270409, 0.1649539,
  0.2137443, 0.2580569, 0.1893859, 0.3611669, 0.3699479, 0.2780909, 
    0.2507285, 0.1763038, 0.2163165, 0.2650436, 0.2793459, 0.1956869, 
    0.313024, 0.2532673, 0.2464577, 0.2875223, 0.3014362, 0.3316671, 
    0.3582359, 0.2793627, 0.3251118, 0.3116094, 0.3495205, 0.5974295, 
    0.2105125, 0.1986909, 0.2563655, 0.3366561, 0.2278552,
  0.277523, 0.2573245, 0.1987789, 0.2837235, 0.2990255, 0.3613953, 0.3365465, 
    0.3196227, 0.2889339, 0.3677951, 0.2764816, 0.2071026, 0.2080201, 
    0.2290154, 0.2665921, 0.2886434, 0.286361, 0.2813237, 0.2979274, 
    0.3389046, 0.2766416, 0.2692633, 0.2395315, 0.2174296, 0.1444365, 
    0.09854028, 0.1080073, 0.2093398, 0.2607607,
  0.1240651, 0.1518397, 0.1885431, 0.1614529, 0.1352783, 0.126129, 0.1146012, 
    0.1341069, 0.2089681, 0.2011539, 0.1455378, 0.1735259, 0.1758005, 
    0.1506383, 0.1099704, 0.1135206, 0.1372899, 0.1469161, 0.137644, 
    0.1111045, 0.1417002, 0.1374098, 0.172084, 0.1854435, 0.1779546, 
    0.2032171, 0.1555387, 0.1338066, 0.1340044,
  0.1396486, 0.08463793, 0.07663009, 0.1223483, 0.111765, 0.106686, 
    0.1283294, 0.1042958, 0.07227463, 0.0828978, 0.05505411, 0.03021393, 
    0.07507172, 0.1518145, 0.113596, 0.07329074, 0.07614409, 0.07160175, 
    0.06639195, 0.1353054, 0.1290059, 0.140049, 0.1810734, 0.04200686, 
    0.07804094, 0.1181121, 0.1001306, 0.1560955, 0.1204474,
  0.005152781, 0.001295251, 0.07485307, 0.06962691, 0.01734067, 0.03523247, 
    0.01939536, 0.06049449, 0.07049502, 0.003811633, 0.0005811334, 
    7.084541e-06, 0.03664077, 0.1348233, 0.1068439, 0.0725241, 0.07753111, 
    0.1185154, 0.2581519, 0.04779989, 0.1024059, 0.005129679, 0.03909343, 
    1.009669e-07, 0.0288359, 0.07892325, 0.1198723, 0.0619139, 0.006272985,
  9.575747e-07, -0.0003389089, 0.05712689, 0.02553734, 0.05812359, 0.106222, 
    0.002418796, 0.01335047, 2.871999e-06, -9.63979e-07, 0.003397348, 
    0.001921939, 0.006144308, 0.01486643, 0.05701595, 0.04827638, 0.02887253, 
    0.08821154, 0.05462895, 0.03533287, 9.762178e-07, 2.121727e-07, 
    1.235929e-07, 2.112873e-05, 0.05878395, 0.238757, 0.06377389, 
    0.001636742, 3.08942e-06,
  4.205367e-07, 0.002147347, 0.0958509, 0.05694238, 0.04552781, 0.1280767, 
    0.1238191, 0.05193511, 0.01527907, 0.006161697, 0.00314486, 0.002564632, 
    0.008116685, 0.04326554, 0.05827222, 0.0491741, 0.03638323, 0.01538335, 
    0.01064352, 4.245913e-06, 1.138264e-08, 5.991769e-08, 1.614695e-06, 
    0.07229935, 0.1672268, 0.1489707, 0.003589835, 3.765683e-07, 1.444373e-07,
  0.1362441, 0.2265566, 0.1259951, 0.0808771, 0.012038, 0.05999327, 
    0.01126531, 0.004368505, 0.2042709, 0.2187043, 0.02605053, 0.009876816, 
    0.01474405, 0.03254688, 0.01448396, 0.01754131, 0.006743899, 
    0.0001374912, 3.257572e-05, 9.42646e-05, 0.0006836544, 0.01583778, 
    0.04129668, 0.1404887, 0.1717417, 0.03963703, 0.1498159, 0.0309507, 
    0.05680378,
  1.19579e-05, 3.527187e-05, 0.003203947, 0.1205242, 0.07993697, 0.0439488, 
    0.0819495, 0.06223961, 0.07462011, 0.1497648, 0.1128456, 0.03106819, 
    0.07580402, 0.07848684, 0.08626374, 0.04866881, 0.06964844, 0.0730136, 
    0.04248461, 0.1708751, 0.1579336, 0.04739526, 0.03613218, 0.009864867, 
    0.02103597, 0.01329435, 0.01989921, 0.000680094, 0.0005318538,
  2.939553e-06, 3.193261e-07, -2.322701e-07, 1.867729e-05, 7.677083e-08, 
    0.02139282, 0.03640769, 0.007699165, 0.03833795, 0.05651663, 0.1439588, 
    0.05741409, 0.01722493, 0.01365658, 0.000937769, 0.001986758, 0.04157299, 
    0.004092517, 0.01890449, 0.000623999, 0.00165014, 0.2083006, 0.042438, 
    0.0204221, 0.02900338, 0.06333688, 0.017541, 0.01898129, 1.885062e-05,
  -8.910611e-05, 0.0152415, 0.01623019, 0.01862847, 0.04380229, 0.04973246, 
    0.05371347, 0.1679956, 0.1852871, 0.09321914, 0.01651989, 0.05202384, 
    0.08425407, 0.09299059, 0.09220161, 0.07610871, 0.07989806, 0.06372975, 
    0.05081951, 2.407174e-05, 0.02215572, 0.01345737, 0.061799, 0.04519407, 
    0.04586185, 0.08359673, 0.04663571, 0.06991229, 0.01253457,
  0.04914607, 0.09510485, 0.1461928, 0.2274499, 0.07829459, 0.01657431, 
    0.1330942, 0.04816755, 0.01372832, 0.0218204, 0.1015487, 0.157889, 
    0.172527, 0.1677052, 0.1768606, 0.1586745, 0.2173392, 0.1986816, 
    0.09288159, 0.1177937, 0.04142501, 0.0111416, 0.07345445, 0.1101836, 
    0.2027351, 0.1259106, 0.1875828, 0.04977383, 0.05530076,
  0.148243, 0.2486202, 0.2578262, 0.2198774, 0.1680882, 0.1179434, 
    0.08022848, 0.1117948, 0.1351452, 0.1648699, 0.1272521, 0.2103347, 
    0.2924702, 0.2788345, 0.2103617, 0.2263611, 0.2264192, 0.2625273, 
    0.2160197, 0.2531694, 0.1496364, 0.1624659, 0.2811207, 0.3249224, 
    0.21645, 0.1467174, 0.1512767, 0.2299334, 0.1541805,
  0.2782463, 0.3965451, 0.4631102, 0.3469552, 0.2945456, 0.3306219, 
    0.2627915, 0.3361399, 0.3047868, 0.2748967, 0.2647786, 0.1158863, 
    0.2009354, 0.1174499, 0.1998245, 0.2378844, 0.1891598, 0.340361, 
    0.2973464, 0.2769464, 0.2159243, 0.4056641, 0.3968679, 0.3319691, 
    0.4217553, 0.5592895, 0.3197226, 0.3131101, 0.2942621,
  0.2582023, 0.3184314, 0.3163348, 0.4431402, 0.5606124, 0.5500625, 
    0.4125835, 0.5677402, 0.4873284, 0.3074116, 0.1971453, 0.2475165, 
    0.2488978, 0.2555698, 0.2736624, 0.1312756, 0.1561441, 0.1948092, 
    0.1757154, 0.1611212, 0.1093654, 0.3022678, 0.2292921, 0.3332075, 
    0.1699826, 0.385464, 0.3540665, 0.2203862, 0.2606852,
  0.1664248, 0.2187071, 0.1074891, 0.05360487, 0.06523585, 0.02617597, 
    0.02372428, 0.02346673, 0.09160405, 0.1279167, 0.2053268, 0.2404604, 
    0.3003333, 0.3131271, 0.3375686, 0.3169355, 0.2523769, 0.1945295, 
    0.2005955, 0.2353318, 0.1333171, 0.1876266, 0.08119618, 0.01789838, 
    0.04403878, 0.04422449, 0.05112687, 0.05288976, 0.1803615,
  0.238776, 0.2337206, 0.2286652, 0.2236098, 0.2185544, 0.2134991, 0.2084437, 
    0.2298099, 0.2294468, 0.2290837, 0.2287206, 0.2283575, 0.2279944, 
    0.2276313, 0.211704, 0.2210875, 0.230471, 0.2398545, 0.249238, 0.2586215, 
    0.268005, 0.2699816, 0.2660165, 0.2620515, 0.2580865, 0.2541215, 
    0.2501564, 0.2461914, 0.2428203,
  0.216827, 0.1110514, 0.06367097, 0.02421629, 0.03800539, 0.0365846, 
    0.03514581, 0.0136164, 0.02204084, 0.103753, 0.1168663, 0.09984481, 
    0.1767212, 0.1665749, 0.03457789, 0.01087816, 0.08654231, 0.1203316, 
    0.1666342, 0.1456665, 0.2744735, 0.533072, 0.4007272, 0.2327475, 
    0.1614954, 0.1276675, 0.1297847, 0.2163564, 0.1945633,
  0.206843, 0.2373919, 0.1754251, 0.3509207, 0.3549431, 0.2861145, 0.2621978, 
    0.1625846, 0.2244307, 0.2807855, 0.2706858, 0.2027539, 0.2853851, 
    0.1916714, 0.2429254, 0.2877229, 0.3394526, 0.3061652, 0.3333643, 
    0.2390152, 0.2928748, 0.3442659, 0.2962984, 0.6063978, 0.1636451, 
    0.1818538, 0.2618543, 0.3177317, 0.2059437,
  0.2234956, 0.2381596, 0.2049674, 0.2682719, 0.3510031, 0.3803745, 0.340539, 
    0.3240945, 0.3000705, 0.3760136, 0.3007351, 0.2432547, 0.2264172, 
    0.2593638, 0.2894518, 0.2967175, 0.2950922, 0.2828062, 0.3095035, 
    0.3389068, 0.2983407, 0.2746603, 0.2718869, 0.2308758, 0.1443943, 
    0.1145878, 0.1068807, 0.1540185, 0.2143041,
  0.1346181, 0.1551816, 0.2077234, 0.1680896, 0.1406864, 0.1189019, 
    0.1060848, 0.1577395, 0.2468701, 0.2146232, 0.1730358, 0.208747, 
    0.1772045, 0.1685148, 0.1178192, 0.1349908, 0.1500818, 0.1544651, 
    0.152721, 0.1214277, 0.1508893, 0.1754909, 0.2061959, 0.2018062, 
    0.1713726, 0.2269749, 0.1598752, 0.1363249, 0.1379962,
  0.1404373, 0.09617266, 0.1106358, 0.1512904, 0.1292028, 0.1116593, 
    0.1434824, 0.1047821, 0.1031733, 0.07322105, 0.05426113, 0.03190435, 
    0.07873224, 0.176672, 0.1281859, 0.07971922, 0.09524969, 0.08198515, 
    0.06727798, 0.1329137, 0.1273094, 0.1494811, 0.2038409, 0.05310285, 
    0.05714243, 0.09801757, 0.1087327, 0.1597914, 0.1403523,
  0.004546256, 0.002003811, 0.05321098, 0.04744566, 0.02378642, 0.03261844, 
    0.02216902, 0.05733922, 0.07206209, 0.002490397, 1.729886e-05, 
    2.762482e-06, 0.03353605, 0.1114067, 0.1286844, 0.07102293, 0.06623009, 
    0.1092843, 0.233019, 0.05250249, 0.09869228, 0.01671899, 0.03158931, 
    3.033727e-07, 0.03058713, 0.05608961, 0.1026418, 0.05496036, 0.02114029,
  8.122963e-07, -6.089978e-05, 0.03672333, 0.02111289, 0.05725869, 0.1164711, 
    0.01070829, 0.02375838, -2.206465e-05, 3.11499e-07, 0.001676397, 
    0.0002759671, 0.006303079, 0.0112238, 0.05682591, 0.04979229, 0.02985709, 
    0.08823086, 0.0512928, 0.05585615, 0.00164875, 2.081291e-05, 
    4.557996e-08, 1.172304e-05, 0.05072311, 0.2330215, 0.06197054, 
    0.006576332, 0.000526692,
  2.368118e-07, -0.0006693276, 0.0860525, 0.0598523, 0.05392076, 0.1075227, 
    0.1279557, 0.06033408, 0.02240159, 0.006762241, 0.002073052, 0.002453177, 
    0.013659, 0.03978214, 0.05185842, 0.05410368, 0.03180173, 0.0316502, 
    0.02638093, 0.001265189, 1.237293e-07, 4.091077e-08, 9.341341e-07, 
    0.05972281, 0.1496945, 0.120301, 0.008230158, 8.629931e-07, 2.06017e-07,
  0.1094506, 0.1618127, 0.1146735, 0.1014729, 0.01747542, 0.0564268, 
    0.01308665, 0.005813059, 0.2002044, 0.2282065, 0.0275178, 0.01208627, 
    0.01904166, 0.03110108, 0.01512357, 0.01880603, 0.007163638, 
    0.0003378874, 0.002729412, 0.0003401053, 0.01671868, 0.02243443, 
    0.02493559, 0.122449, 0.1634484, 0.02818142, 0.1612997, 0.05012435, 
    0.08824725,
  1.389882e-05, 1.046703e-05, 0.0002046277, 0.08029848, 0.09098116, 
    0.04257346, 0.08516329, 0.06409597, 0.0838399, 0.1448645, 0.1132383, 
    0.03401888, 0.07171159, 0.07881138, 0.08911058, 0.05678393, 0.07137241, 
    0.07697085, 0.04328929, 0.1921524, 0.1438188, 0.04830582, 0.05559976, 
    0.01260988, 0.02257689, 0.01907402, 0.01935684, 0.0009108426, 0.0004886435,
  9.411292e-07, 1.248123e-07, 5.814857e-08, -4.905243e-06, 3.837929e-08, 
    0.02061189, 0.05852963, 0.01508334, 0.03579953, 0.06045289, 0.1151889, 
    0.07055157, 0.02249223, 0.02467438, 0.01171757, 0.009836578, 0.04433644, 
    0.01504372, 0.01957471, 0.01276413, 0.005270857, 0.218612, 0.04211759, 
    0.03065644, 0.03819527, 0.06822653, 0.03201732, 0.001081775, 1.196947e-05,
  0.001999045, 0.02449226, 0.01948016, 0.02776423, 0.0443654, 0.04802378, 
    0.02513013, 0.1382755, 0.1468583, 0.08977098, 0.02063937, 0.05787577, 
    0.08940426, 0.1055843, 0.09339595, 0.07826551, 0.08904231, 0.06787141, 
    0.05791538, 0.00064201, 0.01499685, 0.01215821, 0.06872664, 0.04499732, 
    0.05773356, 0.08297744, 0.05367715, 0.05434812, 0.01289229,
  0.04860613, 0.1088658, 0.1565386, 0.2208073, 0.08455181, 0.02703987, 
    0.1385403, 0.04086932, 0.007721876, 0.02701968, 0.1006289, 0.1906871, 
    0.1882158, 0.1827486, 0.2013816, 0.1688253, 0.2458341, 0.2087048, 
    0.1005154, 0.1362656, 0.04371062, 0.007597957, 0.0872362, 0.1078012, 
    0.2110674, 0.1187658, 0.189531, 0.05806319, 0.0740094,
  0.178496, 0.2810337, 0.2871062, 0.2153925, 0.1458413, 0.1556741, 
    0.07228554, 0.1228122, 0.1202698, 0.1848888, 0.1490568, 0.2212134, 
    0.3095289, 0.3162749, 0.1982681, 0.2277882, 0.2601082, 0.3017577, 
    0.224328, 0.2753997, 0.1135675, 0.1717934, 0.2917899, 0.3302523, 
    0.2064218, 0.1699666, 0.1684263, 0.2405103, 0.1849096,
  0.2783032, 0.3835564, 0.4308232, 0.3983082, 0.3129161, 0.2954827, 
    0.2403477, 0.3431118, 0.3314945, 0.3800913, 0.3491104, 0.0910396, 
    0.2172355, 0.09135947, 0.2200849, 0.2763045, 0.145588, 0.3495087, 
    0.2585793, 0.2463222, 0.1818919, 0.3436989, 0.4324034, 0.3201966, 
    0.4546984, 0.5588269, 0.3514862, 0.3097328, 0.3127629,
  0.2620521, 0.2921444, 0.2659811, 0.4705095, 0.5872929, 0.5202999, 0.472494, 
    0.5571879, 0.4498733, 0.2786609, 0.1753875, 0.226362, 0.2268759, 
    0.2409721, 0.2563691, 0.1302791, 0.1000403, 0.1941581, 0.1954326, 
    0.1329861, 0.09371918, 0.2627997, 0.238578, 0.3040385, 0.1833291, 
    0.4237547, 0.3406443, 0.2346408, 0.2442411,
  0.220967, 0.1811437, 0.08735251, 0.03911525, 0.03778593, 0.0191403, 
    0.01943972, 0.02723536, 0.1049106, 0.1655198, 0.2378935, 0.3237918, 
    0.3354371, 0.2603608, 0.2896131, 0.2467226, 0.213345, 0.1838332, 
    0.1203485, 0.2058989, 0.1370445, 0.1476544, 0.05908861, 0.003137587, 
    0.04055543, 0.04433061, 0.05326535, 0.08033343, 0.1902144,
  0.2799259, 0.2782658, 0.2766058, 0.2749457, 0.2732857, 0.2716257, 
    0.2699656, 0.2779865, 0.279418, 0.2808494, 0.2822809, 0.2837123, 
    0.2851438, 0.2865752, 0.2855409, 0.2931437, 0.3007464, 0.3083492, 
    0.315952, 0.3235548, 0.3311575, 0.305636, 0.2982618, 0.2908876, 
    0.2835135, 0.2761393, 0.2687651, 0.2613909, 0.2812539,
  0.2196311, 0.1588986, 0.1110747, 0.03414405, 0.04276517, 0.05207299, 
    0.050586, 0.02800262, 0.09316595, 0.1292991, 0.1426818, 0.1257566, 
    0.1889838, 0.1358131, 0.01702016, 0.007555188, 0.09004191, 0.09510099, 
    0.1828697, 0.1416211, 0.2972434, 0.5440888, 0.390305, 0.219271, 0.146505, 
    0.1003362, 0.1152316, 0.2042263, 0.1919225,
  0.2094136, 0.2580153, 0.2148557, 0.3462369, 0.3607455, 0.3173844, 
    0.2652335, 0.1656065, 0.2320551, 0.2727112, 0.2774148, 0.2050354, 
    0.2581275, 0.1974849, 0.2212264, 0.267594, 0.3128641, 0.2817009, 
    0.3024444, 0.2607794, 0.2732137, 0.3363821, 0.3021104, 0.594831, 
    0.1191774, 0.1473226, 0.2510693, 0.3425604, 0.288576,
  0.2143448, 0.2257403, 0.1990512, 0.2695597, 0.3786442, 0.3548964, 
    0.3129118, 0.3558953, 0.2860486, 0.3638096, 0.3012799, 0.2217331, 
    0.2146206, 0.2603368, 0.2922697, 0.3027409, 0.2997258, 0.2925709, 
    0.3053387, 0.3295652, 0.3115759, 0.265214, 0.2403589, 0.2334394, 
    0.1540736, 0.142601, 0.1221282, 0.1400045, 0.1945508,
  0.1549264, 0.1674796, 0.2035917, 0.1787077, 0.1482139, 0.1086613, 
    0.1298359, 0.1994692, 0.2842693, 0.2167081, 0.232062, 0.2160813, 
    0.2013377, 0.1650872, 0.1031244, 0.1313301, 0.1560352, 0.178801, 
    0.1691395, 0.1437235, 0.1650541, 0.1969974, 0.2181856, 0.217807, 
    0.1292006, 0.222618, 0.178154, 0.1537881, 0.1527779,
  0.1459338, 0.09833367, 0.1451155, 0.1649019, 0.1170255, 0.136445, 
    0.1565406, 0.1221432, 0.1216219, 0.06405886, 0.05737029, 0.03029423, 
    0.07123405, 0.1758416, 0.1477035, 0.08225252, 0.1009991, 0.1062855, 
    0.1180012, 0.1288879, 0.1276799, 0.1700242, 0.2118276, 0.06526564, 
    0.04201851, 0.08610721, 0.1296096, 0.1676769, 0.1484899,
  0.01080274, 0.004124617, 0.039051, 0.04181043, 0.03520929, 0.0372539, 
    0.03316291, 0.05947652, 0.07753123, 0.006638533, 5.664295e-06, 
    1.374542e-06, 0.022175, 0.1058852, 0.1267245, 0.0681416, 0.07534286, 
    0.1030844, 0.2112706, 0.06399571, 0.1060602, 0.06246479, 0.01808632, 
    4.675047e-07, 0.02414107, 0.0459751, 0.1080198, 0.05502278, 0.0419879,
  -2.628354e-06, 4.303786e-05, 0.03447745, 0.01482642, 0.05519403, 0.1250627, 
    0.02197709, 0.03697955, 0.001307172, 1.511977e-07, 0.0008356523, 
    7.923541e-05, 0.005354417, 0.01137882, 0.05701178, 0.04672927, 
    0.03083626, 0.08679202, 0.05382186, 0.07370211, 0.04395203, 0.003298675, 
    3.476452e-07, 2.143776e-05, 0.04831979, 0.202713, 0.05714907, 0.01433908, 
    0.001682259,
  3.301948e-07, 0.001618441, 0.08565591, 0.06884972, 0.06682193, 0.09666416, 
    0.1182681, 0.06872047, 0.02435791, 0.006132662, 0.002821104, 0.00232385, 
    0.01662106, 0.03146137, 0.04191658, 0.0452163, 0.0299735, 0.02583685, 
    0.03620778, 0.03529884, 9.865516e-05, 7.431399e-08, 2.969212e-07, 
    0.04993003, 0.137184, 0.1030775, 0.03202942, 7.137689e-05, 1.060378e-06,
  0.1187477, 0.1325401, 0.1057916, 0.1333252, 0.02568768, 0.06787854, 
    0.01512361, 0.007145638, 0.1884331, 0.2438375, 0.02916372, 0.01143698, 
    0.0186453, 0.02934973, 0.01495582, 0.02047068, 0.0061782, 0.001768988, 
    0.004172997, 0.003527673, 0.02380689, 0.01523632, 0.02107397, 0.1054712, 
    0.1387536, 0.01978623, 0.157143, 0.08784352, 0.09572947,
  9.442791e-06, 1.219272e-06, -4.595732e-06, 0.03545624, 0.103822, 
    0.03687346, 0.08387373, 0.07109135, 0.08880672, 0.1289279, 0.0992799, 
    0.03136246, 0.06001369, 0.07423414, 0.08282191, 0.05474605, 0.07257372, 
    0.07064366, 0.05170729, 0.1929734, 0.136654, 0.04908746, 0.06652751, 
    0.01974374, 0.02308085, 0.02687072, 0.02110777, 0.001367005, -0.0001053716,
  2.50441e-07, 4.265186e-08, 3.513976e-08, 0.0007447887, 2.065222e-09, 
    0.02227841, 0.04417826, 0.01762463, 0.05915255, 0.05149241, 0.09669172, 
    0.07599004, 0.03026205, 0.02840169, 0.03089544, 0.02644092, 0.06275581, 
    0.02546161, 0.0218865, 0.03338114, 0.006445272, 0.2322696, 0.04632951, 
    0.03693052, 0.03254999, 0.05736681, 0.03723083, 3.566028e-05, 6.402722e-06,
  0.004245649, 0.05397263, 0.01764982, 0.03154644, 0.04634185, 0.05128329, 
    0.007159628, 0.09532078, 0.112784, 0.07704523, 0.05060381, 0.08074556, 
    0.1137994, 0.1090775, 0.1108526, 0.09194925, 0.1102126, 0.07413465, 
    0.03707474, 0.0009489257, 0.00754983, 0.01163208, 0.05619255, 0.06098573, 
    0.07542133, 0.07960715, 0.05362776, 0.05774858, 0.01551096,
  0.04386771, 0.1236834, 0.1637756, 0.2308778, 0.07212882, 0.03493561, 
    0.1368641, 0.03593774, 0.006832013, 0.04220228, 0.1012229, 0.2522004, 
    0.2181097, 0.2185205, 0.2151294, 0.1737258, 0.2639156, 0.1947066, 
    0.1134127, 0.1339654, 0.04180821, 0.007744138, 0.1071804, 0.09936196, 
    0.2356911, 0.1122493, 0.1673503, 0.06168317, 0.07789276,
  0.1778848, 0.298687, 0.2577289, 0.2463387, 0.1327823, 0.1469142, 0.1108556, 
    0.1307551, 0.1092553, 0.2018855, 0.184868, 0.251116, 0.3267443, 
    0.3607634, 0.2514439, 0.2539078, 0.2457345, 0.3161918, 0.2428143, 
    0.3120712, 0.103819, 0.1704842, 0.2906195, 0.3042482, 0.231509, 
    0.1956328, 0.1736698, 0.2429182, 0.1958832,
  0.2816315, 0.3678039, 0.3637899, 0.3971061, 0.2443876, 0.2649802, 
    0.1817974, 0.2977363, 0.3679949, 0.4379589, 0.3791537, 0.0824247, 
    0.2473063, 0.1112227, 0.2550758, 0.292144, 0.1600157, 0.3376453, 
    0.2324549, 0.263957, 0.2088746, 0.3667815, 0.4498098, 0.3289257, 
    0.4682727, 0.5131908, 0.3332399, 0.3065615, 0.3291681,
  0.2160427, 0.3112304, 0.2858987, 0.4642521, 0.5121025, 0.5182029, 
    0.4192274, 0.5325633, 0.4222651, 0.3067134, 0.1782849, 0.2212286, 
    0.2020025, 0.2844985, 0.226617, 0.1162512, 0.09078342, 0.1966145, 
    0.1691651, 0.171755, 0.1956785, 0.277139, 0.3026139, 0.291478, 0.1846336, 
    0.42823, 0.3706837, 0.2477083, 0.2262315,
  0.2548214, 0.1372358, 0.07625704, 0.02898012, 0.02480992, 0.02973029, 
    0.01983728, 0.04806924, 0.1321807, 0.1884516, 0.2203715, 0.2790443, 
    0.2999685, 0.2427039, 0.2388961, 0.2321278, 0.1621322, 0.1106967, 
    0.1494432, 0.1880647, 0.117739, 0.1193002, 0.03121204, 0.007194948, 
    0.0442368, 0.05625632, 0.02386296, 0.1244015, 0.2469674,
  0.3002201, 0.297475, 0.2947299, 0.2919848, 0.2892396, 0.2864945, 0.2837494, 
    0.2755067, 0.279977, 0.2844473, 0.2889175, 0.2933879, 0.2978581, 
    0.3023284, 0.3232751, 0.327723, 0.3321709, 0.3366189, 0.3410668, 
    0.3455148, 0.3499627, 0.3358151, 0.329642, 0.3234688, 0.3172957, 
    0.3111226, 0.3049495, 0.2987764, 0.3024162,
  0.2242833, 0.1812991, 0.155789, 0.1081714, 0.05082795, 0.07882443, 
    0.08161075, 0.0413211, 0.1507375, 0.1580151, 0.1671498, 0.1282603, 
    0.2200072, 0.1425995, 0.103468, 0.07353716, 0.08323833, 0.09289877, 
    0.1613488, 0.1247969, 0.3553009, 0.5834666, 0.428441, 0.1728671, 
    0.111754, 0.1111349, 0.1803343, 0.1766436, 0.1920945,
  0.2158034, 0.2554327, 0.1917272, 0.3074841, 0.3432729, 0.3496343, 
    0.2703676, 0.175089, 0.2375271, 0.2969337, 0.2908529, 0.2004971, 
    0.2431786, 0.1757815, 0.2269439, 0.2241321, 0.2800503, 0.2917673, 
    0.2460509, 0.2582866, 0.26301, 0.3269045, 0.3416784, 0.6170096, 
    0.08998509, 0.1595892, 0.2844102, 0.3687057, 0.3244004,
  0.240738, 0.2713662, 0.2621478, 0.3148957, 0.4082867, 0.3620516, 0.3999369, 
    0.3449588, 0.3042274, 0.3712592, 0.270828, 0.2043025, 0.2534681, 
    0.2606817, 0.3031789, 0.2979125, 0.305619, 0.30116, 0.3341242, 0.3621743, 
    0.3179831, 0.2898514, 0.2533277, 0.2502275, 0.1340654, 0.1448153, 
    0.1330011, 0.2322834, 0.2601409,
  0.1800469, 0.2069401, 0.2047021, 0.2058385, 0.1830186, 0.1099196, 
    0.1578168, 0.2754411, 0.2758892, 0.2386225, 0.3198993, 0.2401795, 
    0.223869, 0.1622147, 0.09110907, 0.1663995, 0.1784401, 0.206614, 
    0.1969599, 0.1732042, 0.1799811, 0.2433536, 0.286505, 0.2387439, 
    0.1020632, 0.2286187, 0.2022377, 0.1999651, 0.191195,
  0.2280711, 0.1698481, 0.1811946, 0.1699266, 0.1224566, 0.1702533, 
    0.1617357, 0.1610404, 0.1393649, 0.09236857, 0.07108497, 0.05778781, 
    0.08090288, 0.1654608, 0.1698619, 0.09624089, 0.1250501, 0.164792, 
    0.1435489, 0.1378248, 0.1708449, 0.19886, 0.2466621, 0.07168029, 
    0.03216152, 0.09924725, 0.1531978, 0.1877826, 0.1484494,
  0.03431361, 0.01246734, 0.03395765, 0.05077984, 0.05417419, 0.04678089, 
    0.04052604, 0.08948219, 0.08791828, 0.01389775, -2.968123e-05, 
    7.938661e-07, 0.04599534, 0.1092945, 0.143871, 0.08648416, 0.09066084, 
    0.1109349, 0.2165284, 0.0772741, 0.1092656, 0.09997641, 0.03143959, 
    6.632153e-07, 0.0138462, 0.04566956, 0.1247341, 0.06316467, 0.06097182,
  0.0004433902, -3.650293e-07, 0.03275611, 0.01239767, 0.04557004, 
    0.09721576, 0.04382632, 0.04834066, 0.007896648, 8.36403e-08, 
    0.0002550467, 1.467843e-05, 0.00548714, 0.0163748, 0.06269598, 0.0445405, 
    0.02705377, 0.08208735, 0.05519477, 0.09082814, 0.08915809, 0.02573279, 
    3.426624e-06, 6.595918e-05, 0.06047234, 0.1883269, 0.06111886, 
    0.06458557, 0.01217861,
  3.982619e-06, 0.001471694, 0.08496891, 0.07399724, 0.07224968, 0.0928157, 
    0.1054819, 0.06947006, 0.02831082, 0.008273935, 0.003843232, 0.003100126, 
    0.02423207, 0.02821792, 0.0327875, 0.04022859, 0.02683173, 0.02328184, 
    0.02558155, 0.0405975, 0.009021296, 2.656826e-07, 5.73299e-07, 
    0.04298434, 0.1283106, 0.09724052, 0.05191386, 0.005134105, 6.535219e-05,
  0.111945, 0.1344318, 0.09771161, 0.1602913, 0.02607746, 0.06446973, 
    0.01597504, 0.007423652, 0.1766331, 0.2514728, 0.02771306, 0.01242498, 
    0.01884721, 0.02853505, 0.01442802, 0.02113056, 0.007318628, 0.002081532, 
    0.003343455, 0.0004083508, 0.007783585, 0.008867257, 0.01969672, 
    0.08793464, 0.1067286, 0.019981, 0.1466008, 0.08607298, 0.10022,
  8.088842e-06, 1.773123e-07, -6.587815e-07, 0.01551434, 0.1029139, 
    0.03301524, 0.07979947, 0.06060212, 0.08256734, 0.1144445, 0.08233139, 
    0.0311719, 0.04752206, 0.06056752, 0.06912922, 0.048971, 0.0758765, 
    0.06454329, 0.05965214, 0.1715306, 0.1287999, 0.04339262, 0.05863708, 
    0.02796697, 0.02528386, 0.02931482, 0.019244, 0.001186798, 4.093269e-05,
  8.682039e-08, 1.961766e-08, 2.681485e-08, 0.02199969, -3.043783e-06, 
    0.01784358, 0.03856092, 0.01619706, 0.07424956, 0.06806794, 0.1199499, 
    0.09335475, 0.04201193, 0.02929189, 0.04130606, 0.05274298, 0.08318433, 
    0.03787192, 0.01634217, 0.02520976, 0.01076357, 0.2489056, 0.05310735, 
    0.04216188, 0.02708399, 0.04098027, 0.03547838, 0.0007408942, 2.574247e-06,
  0.000165828, 0.04463462, 0.0238311, 0.03888037, 0.04883726, 0.054162, 
    0.001654139, 0.05946723, 0.1071464, 0.05597453, 0.1393882, 0.1498259, 
    0.1492135, 0.1473849, 0.1488511, 0.1166595, 0.1255008, 0.07788626, 
    0.06628017, 0.001151349, 0.005166751, 0.02494477, 0.04183004, 0.06740414, 
    0.08899539, 0.07336641, 0.04478928, 0.06445482, 0.01628241,
  0.0342121, 0.1535422, 0.1741877, 0.2209317, 0.05475976, 0.01822264, 
    0.1336126, 0.02861254, 0.003621378, 0.03991875, 0.1058468, 0.3045707, 
    0.2742888, 0.2288561, 0.2245214, 0.1983921, 0.2856047, 0.220345, 
    0.1153872, 0.1287491, 0.03374561, 0.00782928, 0.1040575, 0.1231811, 
    0.2802833, 0.1435076, 0.1925731, 0.08249265, 0.09143325,
  0.1776412, 0.3289686, 0.2902806, 0.31097, 0.1427574, 0.1280811, 0.09067998, 
    0.1272122, 0.09701061, 0.216093, 0.2514254, 0.2775103, 0.3753411, 
    0.3726523, 0.3140223, 0.313871, 0.3458099, 0.3647216, 0.3281399, 
    0.3322881, 0.1253246, 0.1936033, 0.319714, 0.3190289, 0.2522407, 
    0.2580868, 0.2111916, 0.2710469, 0.1908648,
  0.2921241, 0.3939612, 0.3503697, 0.4304473, 0.2292611, 0.2283162, 
    0.2362988, 0.3820596, 0.3898681, 0.4604919, 0.3714634, 0.09099388, 
    0.2343103, 0.174365, 0.2616125, 0.3266154, 0.1847599, 0.3634951, 
    0.2372613, 0.3157005, 0.2250475, 0.3643238, 0.4833423, 0.2574982, 
    0.4830345, 0.4598669, 0.3150345, 0.2932715, 0.3423865,
  0.2177562, 0.2666396, 0.2897947, 0.4383181, 0.4722683, 0.5016301, 
    0.3895317, 0.525404, 0.4223046, 0.3383639, 0.1919834, 0.2342574, 
    0.2068946, 0.2910675, 0.2138292, 0.09376567, 0.1670576, 0.2127177, 
    0.1196281, 0.1893312, 0.2311039, 0.2860866, 0.2343231, 0.2815642, 
    0.1846712, 0.4213295, 0.3335723, 0.265894, 0.2411815,
  0.2247702, 0.1181207, 0.08128463, 0.04750244, 0.02029029, 0.04147005, 
    0.02649109, 0.04904909, 0.1178596, 0.1699667, 0.2664792, 0.2780031, 
    0.3279032, 0.2164389, 0.1972635, 0.2185714, 0.158304, 0.1675783, 
    0.1457005, 0.2007238, 0.1057472, 0.1378609, 0.0351005, 0.04720331, 
    0.06803488, 0.08195901, 0.01341986, 0.1598622, 0.3000725,
  0.3265011, 0.3241398, 0.3217785, 0.3194172, 0.3170559, 0.3146946, 
    0.3123334, 0.3143168, 0.3196486, 0.3249804, 0.3303123, 0.3356441, 
    0.3409759, 0.3463077, 0.3529425, 0.3568991, 0.3608556, 0.3648121, 
    0.3687686, 0.3727251, 0.3766817, 0.3605694, 0.3536423, 0.3467153, 
    0.3397883, 0.3328612, 0.3259342, 0.3190071, 0.3283902,
  0.2296282, 0.2018863, 0.2011246, 0.1289493, 0.07698777, 0.1166365, 
    0.1326552, 0.08564242, 0.1578404, 0.1650173, 0.1541775, 0.1355216, 
    0.2408399, 0.1193925, 0.1834621, 0.1647054, 0.07144677, 0.1008392, 
    0.1226891, 0.1287081, 0.3999272, 0.6019851, 0.5024782, 0.1861239, 
    0.1101698, 0.1423036, 0.1508683, 0.1543528, 0.2007756,
  0.2685463, 0.2414003, 0.2094575, 0.280715, 0.314158, 0.3630994, 0.2335793, 
    0.1891196, 0.2437022, 0.3092245, 0.2935859, 0.1872412, 0.2380297, 
    0.1770124, 0.2486709, 0.3134781, 0.3297932, 0.2939467, 0.3088499, 
    0.2862389, 0.3248363, 0.3192328, 0.3521187, 0.6398117, 0.07398371, 
    0.159278, 0.370011, 0.4417082, 0.3052603,
  0.3404077, 0.3320656, 0.3216844, 0.3930191, 0.4376056, 0.41673, 0.4511429, 
    0.3676433, 0.3788199, 0.3376021, 0.2716697, 0.2775344, 0.2711243, 
    0.3027773, 0.3117956, 0.2950829, 0.312053, 0.3178868, 0.3035167, 
    0.359367, 0.3268988, 0.3133869, 0.2767166, 0.2606348, 0.1646844, 
    0.1806277, 0.202502, 0.2247845, 0.3015781,
  0.2726045, 0.2893857, 0.2866417, 0.2666468, 0.1939226, 0.1472084, 
    0.2273357, 0.3449082, 0.3206107, 0.322064, 0.323667, 0.2993747, 
    0.2615263, 0.2042944, 0.1367734, 0.1886965, 0.2006909, 0.1914997, 
    0.2112866, 0.2266348, 0.2745805, 0.3248299, 0.3253209, 0.2052408, 
    0.08406287, 0.2452693, 0.2403476, 0.2233138, 0.2501392,
  0.3063675, 0.2376614, 0.1931616, 0.212194, 0.166733, 0.1674516, 0.2164617, 
    0.22381, 0.2257176, 0.150295, 0.09852125, 0.1263366, 0.1024973, 
    0.1891297, 0.1729983, 0.1103745, 0.1442777, 0.1765033, 0.1796536, 
    0.1980714, 0.2319056, 0.2451786, 0.3058996, 0.07841879, 0.02730305, 
    0.1472351, 0.2086324, 0.236467, 0.2117836,
  0.07840996, 0.05298163, 0.028781, 0.08766069, 0.1298757, 0.1101572, 
    0.1230072, 0.1246545, 0.1282602, 0.03048727, -5.125563e-05, 5.4656e-07, 
    0.0589465, 0.1384896, 0.1458191, 0.09348018, 0.09071007, 0.1363041, 
    0.2051338, 0.1085345, 0.1524934, 0.1273001, 0.06774653, 1.575834e-06, 
    0.0086729, 0.06456917, 0.1342809, 0.09577354, 0.09911255,
  0.03338996, 1.814956e-07, 0.0245474, 0.01472481, 0.04421682, 0.07103297, 
    0.05779851, 0.0785785, 0.01807619, 4.458313e-08, 0.0001131949, 
    2.678431e-07, 0.01191574, 0.02574509, 0.0620084, 0.04209514, 0.02858709, 
    0.08354545, 0.05306624, 0.07191217, 0.1255803, 0.1857647, 0.0009203461, 
    0.00010789, 0.05842727, 0.2106293, 0.05295191, 0.1529892, 0.1110836,
  0.0007144026, 0.001653237, 0.06961942, 0.08499165, 0.07467658, 0.09028546, 
    0.08898279, 0.06148309, 0.03283265, 0.0107703, 0.004678006, 0.005226631, 
    0.02999889, 0.0280046, 0.0275983, 0.03970286, 0.02937227, 0.02568472, 
    0.02632226, 0.03509992, 0.04392169, 3.736107e-05, 5.525092e-06, 
    0.03877232, 0.1116003, 0.07643053, 0.06545575, 0.04454434, 0.007070832,
  0.09724628, 0.1233215, 0.09276112, 0.1651729, 0.02293667, 0.05258187, 
    0.01888239, 0.01103977, 0.1886315, 0.2664768, 0.02651335, 0.01575294, 
    0.02491157, 0.0265988, 0.01649313, 0.02381628, 0.008568793, 0.004174277, 
    0.01034541, 0.005576606, 0.0001470051, 0.003127192, 0.01661754, 
    0.07409793, 0.08548116, 0.02580081, 0.1235914, 0.08599469, 0.1129997,
  3.835584e-06, 6.023196e-08, -6.721539e-07, 0.00449551, 0.08863059, 
    0.03166836, 0.06297314, 0.05095817, 0.0855602, 0.1044643, 0.07372057, 
    0.02912815, 0.03898029, 0.05103865, 0.05865584, 0.04337616, 0.07525485, 
    0.06423157, 0.06384362, 0.1440691, 0.1185476, 0.03766565, 0.05670661, 
    0.03037175, 0.03147841, 0.03573543, 0.02844761, 0.0011365, 2.87032e-05,
  1.846999e-08, 8.724352e-09, 1.732188e-08, 0.04193367, -6.955962e-07, 
    0.04347067, 0.03478943, 0.02154966, 0.09123895, 0.1341676, 0.1729524, 
    0.1210404, 0.05651055, 0.03200543, 0.05116933, 0.06578742, 0.1100385, 
    0.08103545, 0.02605654, 0.02874032, 0.009990295, 0.2595444, 0.06548818, 
    0.05088848, 0.02900423, 0.04078386, 0.04880317, 0.02665265, 9.203926e-07,
  5.411433e-06, 0.02681766, 0.007386079, 0.03916267, 0.04668114, 0.04608874, 
    -0.001209972, 0.0310697, 0.1106346, 0.04979385, 0.2383011, 0.1896507, 
    0.2112952, 0.172237, 0.1500212, 0.1210056, 0.1505887, 0.07060996, 
    0.1598319, 0.01691631, 0.0022471, 0.03312246, 0.04372744, 0.1274088, 
    0.09439387, 0.08540643, 0.04656439, 0.1083387, 0.02293221,
  0.01720836, 0.1094228, 0.1669491, 0.2174744, 0.05345159, 0.05253666, 
    0.117923, 0.01708829, 0.001722915, 0.03499156, 0.1084708, 0.3618161, 
    0.2393483, 0.1863167, 0.171887, 0.1856463, 0.2936649, 0.2355621, 
    0.1630624, 0.1394951, 0.02733151, 0.01897273, 0.1501283, 0.1600674, 
    0.3144384, 0.1746026, 0.206351, 0.1350912, 0.1328793,
  0.1780026, 0.3591994, 0.3827405, 0.3395103, 0.1423888, 0.1640862, 
    0.1249041, 0.1443201, 0.1051446, 0.2969443, 0.224985, 0.2787981, 
    0.4365661, 0.4195354, 0.2586996, 0.3746186, 0.3638302, 0.4223993, 
    0.4061563, 0.3276653, 0.1306082, 0.2250767, 0.3583937, 0.3259266, 
    0.261647, 0.2825796, 0.2772537, 0.3016399, 0.2062376,
  0.2782756, 0.3895093, 0.4108357, 0.4984843, 0.282845, 0.2405387, 0.2792867, 
    0.4307847, 0.4172789, 0.4560916, 0.3882648, 0.09886468, 0.2398991, 
    0.2178822, 0.3629684, 0.3818573, 0.2138118, 0.3693625, 0.2610526, 
    0.3660922, 0.2501282, 0.3971847, 0.5134906, 0.2943874, 0.4777439, 
    0.397337, 0.3021536, 0.3055117, 0.3297872,
  0.2378523, 0.2518153, 0.2863632, 0.4206396, 0.4808342, 0.5187066, 
    0.4049958, 0.5540336, 0.4559388, 0.4071112, 0.2540008, 0.25846, 
    0.2083668, 0.3223987, 0.276533, 0.09861933, 0.1818827, 0.2524225, 
    0.1179283, 0.2352891, 0.2558812, 0.2577314, 0.2625284, 0.360177, 
    0.2163499, 0.4032405, 0.347143, 0.3074046, 0.3283578,
  0.1992295, 0.1296505, 0.106952, 0.03758689, 0.04921017, 0.07711119, 
    0.09097972, 0.07479001, 0.1083795, 0.1994218, 0.3129733, 0.2903113, 
    0.30862, 0.2878205, 0.2402744, 0.2191187, 0.1802434, 0.2154437, 
    0.2301841, 0.1563963, 0.1239331, 0.1247753, 0.05715666, 0.03740116, 
    0.07553879, 0.09028907, 0.01835212, 0.2043024, 0.2848717,
  0.3487751, 0.3470336, 0.3452922, 0.3435507, 0.3418093, 0.3400678, 
    0.3383264, 0.3334206, 0.339563, 0.3457054, 0.3518478, 0.3579901, 
    0.3641325, 0.3702749, 0.4079563, 0.4117905, 0.4156246, 0.4194587, 
    0.4232929, 0.427127, 0.4309612, 0.3959899, 0.3877548, 0.3795197, 
    0.3712847, 0.3630496, 0.3548145, 0.3465794, 0.3501683,
  0.2373523, 0.2307075, 0.215307, 0.1553158, 0.1112101, 0.1658173, 0.1549346, 
    0.1179588, 0.1535485, 0.1918374, 0.1866677, 0.1654411, 0.2490765, 
    0.0625893, 0.1238789, 0.1377732, 0.07021675, 0.08869102, 0.08268399, 
    0.1206034, 0.4366778, 0.6349097, 0.4886394, 0.1865206, 0.1797855, 
    0.1839847, 0.1338823, 0.1432238, 0.1973358,
  0.2514178, 0.204985, 0.2182841, 0.221697, 0.280117, 0.356667, 0.1874113, 
    0.1983391, 0.2727555, 0.3206498, 0.288189, 0.1777274, 0.2412175, 
    0.1569297, 0.2485604, 0.3235557, 0.3842477, 0.3284727, 0.36449, 
    0.3141251, 0.4084127, 0.3738701, 0.3824099, 0.657306, 0.06560449, 
    0.176866, 0.3505149, 0.4340667, 0.318052,
  0.4384153, 0.3947096, 0.3449329, 0.3831822, 0.4299451, 0.4575267, 0.397805, 
    0.4107115, 0.3938603, 0.3245614, 0.2565255, 0.2593198, 0.2706701, 
    0.3090184, 0.3050613, 0.3429433, 0.3343056, 0.4194051, 0.320102, 
    0.3454065, 0.3147812, 0.3542427, 0.2848921, 0.2625055, 0.2011437, 
    0.2337409, 0.280832, 0.2748909, 0.3423981,
  0.3988892, 0.3201223, 0.3300817, 0.297423, 0.2401894, 0.191169, 0.2937592, 
    0.3317278, 0.3223483, 0.3345265, 0.2970101, 0.2775598, 0.2565871, 
    0.3077396, 0.2187466, 0.208967, 0.2052093, 0.200706, 0.2292733, 
    0.2521081, 0.4071704, 0.3321621, 0.370042, 0.1909263, 0.07752112, 
    0.2910691, 0.3085901, 0.3920816, 0.3068714,
  0.3349266, 0.3087668, 0.172721, 0.2520317, 0.2263511, 0.3203216, 0.4152144, 
    0.3780879, 0.2352235, 0.2236487, 0.1668105, 0.1610205, 0.1414556, 
    0.2284691, 0.2015108, 0.1655872, 0.1781324, 0.215353, 0.2581488, 
    0.2404577, 0.2778592, 0.3142045, 0.387786, 0.08426499, 0.0414543, 
    0.1861826, 0.1914372, 0.2545065, 0.2867921,
  0.1364347, 0.09513837, 0.02447919, 0.1247416, 0.1147097, 0.1691334, 
    0.1662275, 0.1345944, 0.2624019, 0.0248919, -6.585631e-05, 4.053025e-07, 
    0.02437682, 0.1936254, 0.1730392, 0.1241181, 0.1168061, 0.2419903, 
    0.2618837, 0.1568987, 0.2048258, 0.1541227, 0.1986746, 1.939037e-05, 
    0.00669238, 0.157744, 0.1653366, 0.1647234, 0.1424498,
  0.2295284, -0.0002378577, 0.0203957, 0.03723278, 0.05981129, 0.06656873, 
    0.08075139, 0.1084804, 0.1078728, -1.432672e-07, 4.753714e-05, 
    -1.594038e-07, 0.04997142, 0.06466561, 0.09820102, 0.06408158, 
    0.06929088, 0.09374401, 0.05624001, 0.07706348, 0.1464712, 0.3669382, 
    0.09219672, 0.0003027056, 0.04264035, 0.2209973, 0.06192804, 0.2100456, 
    0.2925759,
  0.02362456, 0.01282894, 0.04885761, 0.08872402, 0.07784104, 0.08983926, 
    0.09481268, 0.08147412, 0.05572394, 0.02245184, 0.009449276, 0.01946825, 
    0.04695027, 0.03570927, 0.0616059, 0.06290732, 0.04588882, 0.04218905, 
    0.04491644, 0.07693435, 0.168823, 0.02706853, 0.0004612484, 0.03837706, 
    0.08495193, 0.05706985, 0.1093565, 0.1471192, 0.06451782,
  0.08983628, 0.1006907, 0.08442819, 0.1589339, 0.03964599, 0.05036335, 
    0.02956179, 0.01750274, 0.1740132, 0.2504241, 0.02788542, 0.03132044, 
    0.05786728, 0.02943902, 0.06788167, 0.05109588, 0.03722795, 0.008998559, 
    0.01701159, 0.04243709, 0.006833378, 0.0137272, 0.008267542, 0.05632399, 
    0.05779078, 0.03581997, 0.09993957, 0.08144164, 0.1051359,
  1.792029e-06, 2.981428e-08, -4.454384e-07, 0.002577039, 0.07382828, 
    0.08709069, 0.03180745, 0.07652445, 0.1272016, 0.1051283, 0.06805416, 
    0.03394384, 0.04064865, 0.05881649, 0.08103341, 0.04883516, 0.08300164, 
    0.08825133, 0.07112243, 0.124238, 0.1137152, 0.03654909, 0.04818252, 
    0.03658073, 0.06519782, 0.09284317, 0.1157782, 0.002183042, 4.756781e-06,
  4.802598e-09, 2.998938e-09, 8.950714e-09, 0.0234916, -8.913992e-09, 
    0.04812555, 0.02594546, 0.05562473, 0.1008932, 0.2179159, 0.186702, 
    0.2095581, 0.07264926, 0.04240542, 0.05039592, 0.1071457, 0.107137, 
    0.08186141, 0.1063623, 0.0398504, 0.008208239, 0.2601135, 0.1435638, 
    0.05460518, 0.03968235, 0.05008909, 0.08460191, 0.009878078, 2.731912e-07,
  9.858687e-07, 0.03327117, 0.005742205, 0.04654802, 0.04725349, 0.04756737, 
    -0.002368652, 0.01299031, 0.0822662, 0.03807278, 0.1996502, 0.1134067, 
    0.1448621, 0.1307176, 0.1417988, 0.1167054, 0.1945799, 0.08725474, 
    0.246531, 0.01417704, 0.0004938289, 0.04771542, 0.08006462, 0.122427, 
    0.1145492, 0.1043218, 0.0543212, 0.1237743, 0.02208504,
  0.009557331, 0.06213331, 0.1640843, 0.2214611, 0.08423596, 0.02841842, 
    0.1138439, 0.009181486, 0.0002058842, 0.02692676, 0.1415161, 0.2611041, 
    0.165086, 0.1305988, 0.1561349, 0.1608576, 0.2442819, 0.2636831, 
    0.184969, 0.1569008, 0.03209557, 0.04017773, 0.2543805, 0.1889406, 
    0.2838005, 0.2306665, 0.2130395, 0.1572658, 0.160062,
  0.2430077, 0.442136, 0.3810373, 0.2971965, 0.2127068, 0.1933986, 0.1772373, 
    0.1638675, 0.09248384, 0.3780733, 0.1866124, 0.3497281, 0.4048347, 
    0.4020935, 0.283457, 0.3772061, 0.3445943, 0.3649008, 0.3712701, 
    0.3375765, 0.1492835, 0.2489528, 0.3681319, 0.4062417, 0.2536256, 
    0.2650596, 0.2570044, 0.2882438, 0.2537462,
  0.2350669, 0.3671689, 0.4408885, 0.5311267, 0.3578849, 0.3126883, 
    0.3630331, 0.436258, 0.4519546, 0.5733973, 0.3830121, 0.1106398, 
    0.2417929, 0.22241, 0.5935179, 0.4158402, 0.1961265, 0.358172, 0.3385651, 
    0.3684261, 0.3030217, 0.3759396, 0.3500496, 0.3113603, 0.4206252, 
    0.3259324, 0.3133855, 0.2995506, 0.2888226,
  0.1365264, 0.2005373, 0.3397655, 0.3743221, 0.4543199, 0.4904582, 
    0.4571727, 0.6153082, 0.4804761, 0.3981484, 0.3034882, 0.3013019, 
    0.2466656, 0.3970237, 0.3921919, 0.1206889, 0.1608079, 0.2911701, 
    0.1957968, 0.3315306, 0.2568693, 0.2300854, 0.2720664, 0.3659936, 
    0.2287516, 0.4036536, 0.3445257, 0.2971929, 0.3972816,
  0.1509271, 0.1276117, 0.1693013, 0.08021913, 0.1467267, 0.1823134, 
    0.1716772, 0.1132154, 0.1557463, 0.2718264, 0.3454629, 0.3679946, 
    0.2794281, 0.3556401, 0.2799913, 0.2768231, 0.2547616, 0.2561086, 
    0.2466785, 0.1933331, 0.1834458, 0.1429967, 0.08432326, 0.05384383, 
    0.1005765, 0.1416004, 0.05426599, 0.2247167, 0.247425,
  0.3528084, 0.3508893, 0.3489702, 0.3470512, 0.3451321, 0.3432131, 0.341294, 
    0.3701447, 0.376804, 0.3834634, 0.3901227, 0.396782, 0.4034414, 
    0.4101008, 0.4226991, 0.4277496, 0.4328001, 0.4378507, 0.4429012, 
    0.4479517, 0.4530022, 0.4440689, 0.4342781, 0.4244873, 0.4146965, 
    0.4049056, 0.3951148, 0.385324, 0.3543436,
  0.241697, 0.2572981, 0.233934, 0.1736216, 0.1500542, 0.2004659, 0.2085096, 
    0.1454747, 0.1662514, 0.2004639, 0.2029775, 0.1998732, 0.2517026, 
    0.04003625, 0.093169, 0.130722, 0.1758368, 0.1023867, 0.0785798, 
    0.09587947, 0.4350463, 0.6396369, 0.446343, 0.1872319, 0.1410559, 
    0.1906533, 0.09796525, 0.1082674, 0.1911793,
  0.2374586, 0.2088809, 0.2288851, 0.181173, 0.2413724, 0.3425265, 0.1555856, 
    0.2054793, 0.2737256, 0.3057368, 0.2686813, 0.1580618, 0.2511982, 
    0.1524331, 0.2407704, 0.3452699, 0.3434896, 0.3264166, 0.3700546, 
    0.3628337, 0.4289984, 0.4353926, 0.4177834, 0.6912379, 0.060817, 
    0.204394, 0.3625543, 0.4269533, 0.3030866,
  0.4295866, 0.4393576, 0.4142347, 0.4086854, 0.4471327, 0.4366165, 
    0.3925984, 0.3771354, 0.385562, 0.3278862, 0.2812878, 0.21245, 0.3008402, 
    0.3071461, 0.3054732, 0.407106, 0.3607709, 0.4032846, 0.3358706, 
    0.3208021, 0.3333907, 0.3589998, 0.3480175, 0.3520839, 0.2704021, 
    0.2972058, 0.2773195, 0.375124, 0.388162,
  0.374528, 0.3689116, 0.3451553, 0.3436258, 0.3496975, 0.3027535, 0.3431551, 
    0.3068208, 0.3288903, 0.3500691, 0.2879106, 0.2831059, 0.2834404, 
    0.3686474, 0.2556442, 0.2243795, 0.2530178, 0.2270221, 0.2642941, 
    0.3066252, 0.3820159, 0.3408761, 0.3905986, 0.1880264, 0.07666907, 
    0.3153294, 0.3817213, 0.3085654, 0.3000121,
  0.3186954, 0.2193328, 0.1743073, 0.2458239, 0.2255593, 0.263785, 0.3154837, 
    0.3773333, 0.3330212, 0.2428784, 0.2417599, 0.1223927, 0.1476454, 
    0.2906064, 0.2112433, 0.3059936, 0.2879206, 0.1830184, 0.230723, 
    0.2503644, 0.2819534, 0.2537465, 0.3411457, 0.1019133, 0.0253242, 
    0.1812033, 0.2464256, 0.2736112, 0.3166603,
  0.2969942, 0.1576173, 0.02288772, 0.08037878, 0.1147845, 0.1295797, 
    0.1152552, 0.183462, 0.3030471, 0.04613997, -0.0002050593, 3.211267e-07, 
    0.009439958, 0.1549808, 0.1823617, 0.1607486, 0.1476506, 0.1958552, 
    0.335365, 0.2794807, 0.2829274, 0.1211476, 0.353685, 0.0004798417, 
    0.004351796, 0.08738589, 0.1705821, 0.1283, 0.2130455,
  0.5646813, 0.001086883, 0.0312002, 0.0705463, 0.1086144, 0.06809165, 
    0.09919825, 0.0811696, 0.1318758, -0.0004204952, 5.822482e-05, 
    -8.703608e-09, 0.1234775, 0.08189824, 0.1199682, 0.1339476, 0.1561479, 
    0.1373563, 0.08257024, 0.09513919, 0.110264, 0.2380917, 0.521879, 
    0.001451643, 0.0403538, 0.2162114, 0.06510771, 0.1223054, 0.3703571,
  0.2092967, 0.07256975, 0.03027388, 0.1010358, 0.1014967, 0.09016286, 
    0.1095344, 0.1026478, 0.1594841, 0.07916899, 0.01837418, 0.07860309, 
    0.09196538, 0.05403185, 0.07727144, 0.06244227, 0.06469683, 0.1160989, 
    0.0537328, 0.0413007, 0.1524382, 0.4780381, 0.08306145, 0.01522982, 
    0.05530877, 0.04441427, 0.1250451, 0.1458776, 0.4069812,
  0.08480413, 0.08251277, 0.0696339, 0.1561785, 0.1022214, 0.1113471, 
    0.1363821, 0.08808079, 0.141403, 0.2010037, 0.07117475, 0.05075675, 
    0.1274076, 0.1073053, 0.108845, 0.08983909, 0.1263635, 0.06487754, 
    0.1033734, 0.1079017, 0.1105653, 0.04895968, 0.04765091, 0.03387792, 
    0.03104081, 0.05057722, 0.09553087, 0.08357627, 0.1031456,
  2.983566e-07, 2.010967e-08, -2.035895e-07, -0.0007459425, 0.08584457, 
    0.06450718, 0.01722428, 0.0745166, 0.1747823, 0.1059972, 0.06975839, 
    0.06467463, 0.07074564, 0.08292546, 0.05260238, 0.07328654, 0.08231716, 
    0.1501854, 0.142148, 0.1182319, 0.1488066, 0.04939337, 0.06345349, 
    0.04692396, 0.05250588, 0.06573585, 0.1071304, 0.03365314, 4.617661e-06,
  2.91067e-09, 1.182248e-09, 2.651317e-09, 0.01163948, -4.282109e-09, 
    0.02172337, 0.01196748, 0.03904991, 0.05139648, 0.1694122, 0.1357172, 
    0.1477136, 0.09786589, 0.1147542, 0.1241776, 0.09645206, 0.1431173, 
    0.09043156, 0.3006399, 0.1250428, 0.008562973, 0.2961304, 0.08659387, 
    0.04339753, 0.06433991, 0.04711469, 0.06243985, 0.001753493, 7.523161e-08,
  6.719522e-07, 0.03260841, 0.002477188, 0.07572118, 0.04434847, 0.02863067, 
    -0.002571198, 0.005009756, 0.07572576, 0.02180789, 0.09459641, 
    0.05141971, 0.1001784, 0.1010612, 0.1139785, 0.1070487, 0.1524714, 
    0.06906819, 0.2713258, 0.03599871, 0.0001212442, 0.05997091, 0.08796983, 
    0.08482207, 0.1252583, 0.1157046, 0.06003567, 0.07818603, 0.01908233,
  0.008365502, 0.04156525, 0.1343871, 0.2285434, 0.05948006, 0.008935364, 
    0.1273178, 0.004806481, 6.499869e-05, 0.02386325, 0.1713052, 0.1255905, 
    0.1016157, 0.09793702, 0.1363504, 0.1597808, 0.199844, 0.2703706, 
    0.2323357, 0.1833199, 0.04067811, 0.08188724, 0.3351821, 0.1507682, 
    0.2190654, 0.2668373, 0.2504531, 0.2095005, 0.1454442,
  0.239257, 0.482482, 0.381231, 0.3342612, 0.2806258, 0.1930888, 0.1691366, 
    0.1720838, 0.09836943, 0.3774082, 0.1621718, 0.3476379, 0.2852589, 
    0.3189727, 0.288861, 0.3192121, 0.3663604, 0.3529661, 0.3529193, 
    0.3990017, 0.2027256, 0.305741, 0.338259, 0.5509151, 0.2588233, 0.265929, 
    0.2370681, 0.2853172, 0.228885,
  0.1958985, 0.3803841, 0.5177699, 0.6104738, 0.4375604, 0.325594, 0.4771502, 
    0.4889381, 0.5112813, 0.6134061, 0.4392711, 0.1346947, 0.2211536, 
    0.1391685, 0.7520478, 0.4570915, 0.2219549, 0.3537197, 0.3523246, 
    0.3781172, 0.3819354, 0.3061612, 0.2051396, 0.2595185, 0.286206, 
    0.2541039, 0.2690226, 0.2574095, 0.2563689,
  0.08549732, 0.1064781, 0.2634456, 0.28573, 0.4093304, 0.4921038, 0.5160317, 
    0.6404365, 0.4867639, 0.4284617, 0.3437058, 0.3256964, 0.2813855, 
    0.4701522, 0.4668725, 0.2385215, 0.1906305, 0.2999054, 0.295192, 
    0.4136325, 0.2494711, 0.2731532, 0.2814874, 0.408407, 0.2774012, 
    0.4065171, 0.3459142, 0.2719934, 0.2441272,
  0.207693, 0.1526639, 0.22727, 0.1678331, 0.199119, 0.2528466, 0.2018692, 
    0.1778988, 0.2085339, 0.417744, 0.4261245, 0.451775, 0.3797808, 
    0.4004576, 0.3234645, 0.3001841, 0.3019164, 0.301336, 0.2606693, 
    0.2325064, 0.2901488, 0.2124567, 0.1189532, 0.07419796, 0.1259391, 
    0.1962058, 0.105516, 0.2518778, 0.2951458,
  0.3925946, 0.3916629, 0.3907312, 0.3897996, 0.3888679, 0.3879362, 
    0.3870046, 0.3780113, 0.3841177, 0.3902241, 0.3963305, 0.402437, 
    0.4085434, 0.4146498, 0.4702191, 0.4747642, 0.4793093, 0.4838544, 
    0.4883994, 0.4929445, 0.4974896, 0.4537285, 0.4440086, 0.4342888, 
    0.424569, 0.4148491, 0.4051293, 0.3954094, 0.3933399,
  0.2417884, 0.2529759, 0.2418908, 0.2079934, 0.2061332, 0.2637531, 
    0.2390663, 0.1654162, 0.2044969, 0.2148577, 0.2296527, 0.2107368, 
    0.2733827, 0.03175469, 0.1326971, 0.2755226, 0.2929194, 0.1578376, 
    0.09120903, 0.09592162, 0.4187474, 0.6588048, 0.3784597, 0.1693027, 
    0.1092989, 0.1651726, 0.08354927, 0.08653015, 0.2264883,
  0.2004783, 0.1732479, 0.2168192, 0.1497542, 0.1960888, 0.3279902, 
    0.1176911, 0.201129, 0.2476311, 0.2889951, 0.2308631, 0.1394293, 
    0.1918326, 0.1534603, 0.2660082, 0.3463479, 0.3421409, 0.3051873, 
    0.3734316, 0.4079461, 0.4048788, 0.4506597, 0.4001617, 0.6732029, 
    0.05292336, 0.2557484, 0.4238188, 0.4853258, 0.3400519,
  0.4005255, 0.4466655, 0.4485905, 0.3840031, 0.4408697, 0.4476056, 0.373493, 
    0.325452, 0.3829225, 0.3301539, 0.254698, 0.200805, 0.2975722, 0.3014596, 
    0.3166318, 0.4063306, 0.3755155, 0.3825199, 0.3306653, 0.3217517, 
    0.3359974, 0.3253264, 0.320776, 0.4039045, 0.3156112, 0.3912392, 
    0.2657522, 0.4319252, 0.4355637,
  0.3671325, 0.4023826, 0.3708625, 0.3198042, 0.3102382, 0.2998153, 0.318059, 
    0.3046627, 0.3295221, 0.3327582, 0.2574929, 0.2841015, 0.2375242, 
    0.3286864, 0.2211184, 0.2254231, 0.2581988, 0.3041261, 0.282265, 
    0.3358624, 0.3377191, 0.3905903, 0.3671555, 0.168573, 0.07387206, 
    0.3079186, 0.4442589, 0.3102044, 0.3419777,
  0.257008, 0.2117694, 0.1241946, 0.2039184, 0.1799211, 0.1883478, 0.2525998, 
    0.2743362, 0.3332587, 0.2230771, 0.2095365, 0.1136832, 0.1127117, 
    0.2316221, 0.208295, 0.3600324, 0.2570952, 0.1207852, 0.1756193, 
    0.2034478, 0.2788325, 0.2205811, 0.2704924, 0.1227549, 0.01649215, 
    0.1065859, 0.2244615, 0.2878102, 0.2617336,
  0.1487625, 0.1283748, 0.02062326, 0.05373172, 0.07706052, 0.0739721, 
    0.04952573, 0.1535845, 0.1966237, 0.05316622, -0.0001776086, 
    4.965226e-07, 0.002757151, 0.09062844, 0.1676752, 0.09766483, 0.0799145, 
    0.1362746, 0.278552, 0.1722165, 0.2165609, 0.08128311, 0.2804814, 
    0.01722093, 0.003826956, 0.08967807, 0.1517605, 0.07473783, 0.1163457,
  0.3758602, 0.001166103, 0.03912519, 0.07126876, 0.05451402, 0.03917765, 
    0.05598587, 0.07857022, 0.1895443, -0.0002623455, 3.432162e-05, 
    -3.704132e-06, 0.1263553, 0.02849737, 0.0794612, 0.06527691, 0.04440654, 
    0.162202, 0.08490381, 0.03555099, 0.02894588, 0.06624805, 0.4399548, 
    0.05309252, 0.02386503, 0.1967312, 0.04290201, 0.02162881, 0.1602892,
  0.5039593, 0.2186609, 0.01720283, 0.1432061, 0.1616999, 0.09812683, 
    0.06497125, 0.05139584, 0.07886315, 0.04253851, 0.01066419, 0.04703233, 
    0.06283073, 0.04258853, 0.04355836, 0.02862494, 0.02272034, 0.03152305, 
    0.01141568, 0.009495031, 0.03254568, 0.3951373, 0.5681424, 0.005828731, 
    0.03926067, 0.03449839, 0.02818724, 0.04743212, 0.2470227,
  0.07298742, 0.06333435, 0.04716022, 0.1295308, 0.1751833, 0.07556224, 
    0.1065434, 0.2215972, 0.1033038, 0.1405196, 0.02148259, 0.1033684, 
    0.01581514, 0.02497256, 0.01746898, 0.0410852, 0.05703981, 0.0995629, 
    0.1111499, 0.140193, 0.307619, 0.4163755, 0.08605798, 0.02396455, 
    0.01263748, 0.04070432, 0.0801972, 0.08982565, 0.1001987,
  1.114148e-07, 1.585189e-08, -1.417719e-08, -0.001320505, 0.09478257, 
    0.0719672, 0.01193677, 0.03888589, 0.05021043, 0.08784018, 0.06677877, 
    0.04553333, 0.04500549, 0.03449495, 0.02343752, 0.03408353, 0.04845877, 
    0.07301301, 0.1077148, 0.1047888, 0.09495705, 0.04863808, 0.2440766, 
    0.04503566, 0.01199171, 0.01195161, 0.03764278, 0.006917488, -1.121596e-06,
  2.516547e-09, 6.176095e-10, 8.076916e-10, 0.001643145, -5.127521e-10, 
    0.006881605, 0.007508402, 0.006944099, 0.03281133, 0.06669221, 
    0.06774931, 0.06415732, 0.07061449, 0.03575466, 0.04186007, 0.02221215, 
    0.06987665, 0.09722687, 0.1843417, 0.1476881, 0.03605242, 0.2371047, 
    0.02839205, 0.02048484, 0.06666376, 0.01349524, 0.01113519, 0.0003393161, 
    2.57371e-08,
  4.208507e-07, 0.0225941, 0.008183738, 0.05611863, 0.03930558, 0.02645442, 
    -0.002569659, 0.001641105, 0.07723622, 0.0136583, 0.03961305, 0.03359793, 
    0.07399329, 0.07624095, 0.0941689, 0.07904743, 0.1069544, 0.03585541, 
    0.2595544, 0.04433128, 5.23477e-05, 0.08539527, 0.09401383, 0.03136575, 
    0.06740513, 0.09254019, 0.0146175, 0.02124248, 0.01683987,
  0.005866395, 0.01669283, 0.109947, 0.2182371, 0.03586846, 0.004799365, 
    0.1362397, 0.006408378, 0.0001403738, 0.01765626, 0.1754996, 0.06756088, 
    0.05895733, 0.08360153, 0.119429, 0.1464916, 0.1905144, 0.2598078, 
    0.2308271, 0.2104748, 0.0250209, 0.1220652, 0.3021405, 0.09297691, 
    0.1729088, 0.3095692, 0.2369263, 0.1496008, 0.1251415,
  0.1985848, 0.500821, 0.3781482, 0.3604828, 0.2822872, 0.210696, 0.1508936, 
    0.1587669, 0.09580457, 0.3850892, 0.1246418, 0.3776503, 0.2016278, 
    0.2336, 0.2573345, 0.2825967, 0.3738765, 0.3328898, 0.3094505, 0.441461, 
    0.2008331, 0.2792791, 0.3231614, 0.6232092, 0.2458279, 0.2382345, 
    0.2040362, 0.2922969, 0.2091221,
  0.1672533, 0.422608, 0.509423, 0.6462103, 0.5709016, 0.3754598, 0.5758657, 
    0.6067555, 0.5731904, 0.6588436, 0.5551934, 0.1864847, 0.2115873, 
    0.1344364, 0.5941789, 0.4119997, 0.3274828, 0.3297708, 0.3538833, 
    0.4376219, 0.416214, 0.2797304, 0.128434, 0.2197633, 0.2016908, 
    0.2041512, 0.2460123, 0.2046676, 0.2216035,
  0.06217832, 0.05161676, 0.2130806, 0.1809281, 0.3272478, 0.4575067, 
    0.6227208, 0.6583067, 0.4822389, 0.4952489, 0.424481, 0.313875, 
    0.3213147, 0.5292385, 0.4881753, 0.3697295, 0.2030302, 0.3014867, 
    0.3327699, 0.4782234, 0.3556536, 0.3853613, 0.2856946, 0.3694651, 
    0.1547586, 0.3988174, 0.3439511, 0.2336642, 0.1755417,
  0.1582295, 0.1409416, 0.2621906, 0.1875229, 0.2371575, 0.2892303, 
    0.2964745, 0.2478523, 0.2838351, 0.5408683, 0.5008314, 0.515286, 
    0.4485627, 0.4682244, 0.4129561, 0.424189, 0.3851025, 0.3982913, 
    0.2842446, 0.3308378, 0.3499264, 0.2391822, 0.1631224, 0.09151495, 
    0.1544831, 0.2213119, 0.130028, 0.2911748, 0.3207626,
  0.4333732, 0.435076, 0.4367788, 0.4384816, 0.4401844, 0.4418872, 0.44359, 
    0.4145422, 0.4208896, 0.427237, 0.4335844, 0.4399318, 0.4462792, 
    0.4526266, 0.499061, 0.4992815, 0.499502, 0.4997225, 0.499943, 0.5001635, 
    0.500384, 0.4572372, 0.4489665, 0.4406959, 0.4324251, 0.4241544, 
    0.4158837, 0.407613, 0.4320109,
  0.2514358, 0.2597913, 0.2437338, 0.2205036, 0.231166, 0.3169013, 0.256489, 
    0.1779823, 0.2146095, 0.2253228, 0.2111084, 0.1746459, 0.302775, 
    0.02369971, 0.2184153, 0.2970193, 0.2854543, 0.2249688, 0.1027801, 
    0.08722968, 0.3819547, 0.6240716, 0.341585, 0.1512742, 0.1069684, 
    0.1451609, 0.08287814, 0.09335953, 0.2240234,
  0.1741207, 0.1450321, 0.1773643, 0.1263374, 0.1520932, 0.2972583, 
    0.07727543, 0.1599795, 0.1918993, 0.2443395, 0.1824322, 0.1125633, 
    0.1378272, 0.1298535, 0.274302, 0.3594199, 0.3773324, 0.2839356, 
    0.3785906, 0.3579307, 0.3474522, 0.3803676, 0.3939779, 0.624407, 
    0.04513298, 0.2733725, 0.4294754, 0.4813458, 0.3281667,
  0.3663739, 0.4245587, 0.4292384, 0.3766957, 0.3878835, 0.3980708, 0.359645, 
    0.2873755, 0.3621161, 0.3175999, 0.2143541, 0.1668305, 0.2768728, 
    0.2844571, 0.2910868, 0.3731546, 0.370941, 0.3903156, 0.3354188, 
    0.3200364, 0.3199807, 0.3082495, 0.2659774, 0.3193185, 0.2927455, 
    0.3895265, 0.2917213, 0.4374284, 0.4457068,
  0.3437895, 0.3564337, 0.3643091, 0.2656081, 0.2547832, 0.2667444, 
    0.2816472, 0.2675592, 0.3046066, 0.30942, 0.2221998, 0.2704786, 
    0.1829661, 0.2724061, 0.1882052, 0.2449025, 0.242138, 0.300927, 
    0.2534065, 0.3016441, 0.3068078, 0.3748021, 0.3022381, 0.1538355, 
    0.09968212, 0.3133181, 0.4477554, 0.3155723, 0.3430733,
  0.2357523, 0.1445764, 0.07782627, 0.1802933, 0.1814205, 0.1814432, 
    0.2128164, 0.2168721, 0.2764768, 0.2046771, 0.1570138, 0.06016341, 
    0.05309829, 0.1789082, 0.2089316, 0.2497394, 0.2109807, 0.07415145, 
    0.1203266, 0.2009189, 0.2318279, 0.2092253, 0.2193618, 0.1288242, 
    0.01585083, 0.08201449, 0.1790259, 0.1950648, 0.2472159,
  0.04837506, 0.06896824, 0.01679623, 0.06777896, 0.06040903, 0.03600731, 
    0.02935104, 0.08075235, 0.1129974, 0.02737557, -7.846447e-05, 
    2.043837e-07, 0.002434486, 0.05378914, 0.1212169, 0.07407858, 0.03241757, 
    0.09933279, 0.2422892, 0.1053203, 0.1289623, 0.03093546, 0.130237, 
    0.01982447, 0.004548541, 0.09724125, 0.1423922, 0.02922806, 0.03473894,
  0.1319478, 0.01868955, 0.03025758, 0.03153473, 0.02239813, 0.03402105, 
    0.03693876, 0.03941047, 0.1318749, -5.979488e-05, 1.055424e-05, 
    -3.30189e-06, 0.03738712, 0.0127726, 0.0319121, 0.02602983, 0.01745378, 
    0.07241054, 0.04132502, 0.01399101, 0.006702692, 0.01855647, 0.1801816, 
    0.09671045, 0.01404656, 0.1958602, 0.02088797, 0.004455809, 0.05162995,
  0.2210751, 0.1396365, 0.01008765, 0.2194704, 0.02876602, 0.04981863, 
    0.0280233, 0.01127832, 0.0255152, 0.008249404, 0.006217889, 0.006637427, 
    0.02392725, 0.007492269, 0.01207187, 0.005660768, 0.002023063, 
    0.00579378, 0.0007909412, 0.001764174, 0.009622145, 0.1372666, 0.337906, 
    0.001676638, 0.03637775, 0.03072764, 0.0005812528, 0.00916316, 0.08027099,
  0.0925165, 0.05087318, 0.03403468, 0.1170667, 0.02444755, 0.01932892, 
    0.01298083, 0.02805839, 0.08762959, 0.09386028, 0.007896842, 0.00934619, 
    0.002831128, 0.01018355, 0.005012912, 0.009885991, 0.008957976, 
    0.02442169, 0.02684471, 0.04318218, 0.1287628, 0.4001737, 0.4165929, 
    0.009560987, 0.009204907, 0.008864624, 0.05453546, 0.03856704, 0.1758405,
  -1.189292e-07, 1.453543e-08, 6.855674e-08, -0.0007563547, 0.08126781, 
    0.01181155, 0.007158991, 0.0177198, 0.01132164, 0.06441353, 0.03974426, 
    0.009726592, 0.02118037, 0.0212514, 0.007043356, 0.01098402, 0.02359855, 
    0.03294984, 0.0595888, 0.06524549, 0.06987662, 0.03467782, 0.3321676, 
    0.05248727, 0.0009952575, 0.002018578, 0.01420695, 0.002148638, 
    -3.279766e-07,
  2.388389e-09, 4.914755e-10, 3.023618e-10, -1.209827e-05, 4.732185e-10, 
    0.001914222, 0.005414686, 0.001808068, 0.02784611, 0.01838783, 
    0.03345216, 0.02433109, 0.01488981, 0.007571999, 0.007831955, 
    0.005831091, 0.03526234, 0.0402444, 0.1005136, 0.07771342, 0.007689847, 
    0.1797372, 0.006629094, -0.0001629862, 0.01098717, 0.001694806, 
    0.003100638, 0.0003310697, 1.788469e-08,
  -8.881186e-07, 0.01480324, 0.003745384, 0.04807319, 0.04242856, 0.04232688, 
    -0.002521576, 0.0003562099, 0.07080313, 0.01240043, 0.01891875, 
    0.02794243, 0.05150421, 0.06754407, 0.07451836, 0.04324005, 0.05825857, 
    0.0126067, 0.1870567, 0.06934969, 7.912775e-06, 0.07448985, 0.07218037, 
    0.01811466, 0.03842934, 0.04998171, 0.00234554, 0.008822694, 0.01830008,
  0.002294663, 0.00687594, 0.08050394, 0.2125013, 0.01339579, 0.003995712, 
    0.1452323, 0.005454885, 3.06292e-06, 0.0171447, 0.1660428, 0.0417651, 
    0.04078347, 0.06608734, 0.09874921, 0.1280515, 0.1838487, 0.2337482, 
    0.190037, 0.2149709, 0.01631981, 0.1127063, 0.2478766, 0.06481625, 
    0.1265305, 0.2481187, 0.2045289, 0.07788169, 0.08676367,
  0.1606913, 0.509755, 0.3915536, 0.3699178, 0.2270176, 0.1721312, 0.1370345, 
    0.1495847, 0.07137244, 0.3140504, 0.1096815, 0.4183024, 0.1329571, 
    0.1795318, 0.2171918, 0.2860324, 0.3327771, 0.2922028, 0.2793618, 
    0.4643943, 0.1931027, 0.2446633, 0.3456683, 0.6079284, 0.2047642, 
    0.1941124, 0.1993434, 0.2811337, 0.179529,
  0.1332573, 0.4580454, 0.5095323, 0.7250981, 0.7206861, 0.4182003, 
    0.6531048, 0.6475674, 0.5850128, 0.6734039, 0.7016773, 0.2642148, 
    0.211966, 0.1521169, 0.464803, 0.3418219, 0.3947826, 0.297717, 0.3840744, 
    0.5135575, 0.4418081, 0.216544, 0.08762763, 0.2074113, 0.141599, 
    0.1556412, 0.2216576, 0.1560625, 0.1728713,
  0.03861246, 0.04351377, 0.2280077, 0.1117181, 0.2362592, 0.3865562, 
    0.6240483, 0.6519572, 0.4446628, 0.5023544, 0.4733598, 0.3041815, 
    0.3725414, 0.5732768, 0.5088584, 0.397818, 0.2802386, 0.3176848, 
    0.3707031, 0.4932708, 0.3825227, 0.4923053, 0.2696538, 0.3750874, 
    0.1096466, 0.3979076, 0.3519319, 0.193811, 0.1363489,
  0.198898, 0.2859898, 0.2560771, 0.2501737, 0.2822528, 0.3217539, 0.3583892, 
    0.3469423, 0.4186627, 0.5868359, 0.5919453, 0.5667806, 0.5158936, 
    0.5895329, 0.5256585, 0.4965684, 0.4459285, 0.4388153, 0.4063303, 
    0.4610694, 0.4521732, 0.2338033, 0.201018, 0.1918736, 0.1653682, 
    0.2335409, 0.1324129, 0.3134584, 0.3615485,
  0.42853, 0.4325115, 0.436493, 0.4404745, 0.4444561, 0.4484376, 0.4524191, 
    0.4247464, 0.4330027, 0.4412591, 0.4495155, 0.4577718, 0.4660282, 
    0.4742846, 0.5301347, 0.5240018, 0.5178688, 0.5117359, 0.5056029, 
    0.4994699, 0.493337, 0.4590708, 0.4529659, 0.4468609, 0.440756, 
    0.4346511, 0.4285462, 0.4224413, 0.4253448,
  0.2448828, 0.2613389, 0.2436763, 0.2189588, 0.2272468, 0.286204, 0.2538947, 
    0.1777334, 0.2004431, 0.2081873, 0.1746054, 0.1200662, 0.2355821, 
    0.01220322, 0.2030937, 0.2612, 0.2611914, 0.2513995, 0.1103561, 
    0.07537241, 0.3295403, 0.5354527, 0.294786, 0.1265118, 0.08301089, 
    0.1413025, 0.05701394, 0.09644828, 0.1951326,
  0.1703331, 0.1141518, 0.1485256, 0.09741321, 0.1050257, 0.2629467, 
    0.05054145, 0.1086731, 0.1401581, 0.2034638, 0.1306279, 0.08290596, 
    0.1024584, 0.107595, 0.2529227, 0.3513811, 0.3038005, 0.2693846, 
    0.3178436, 0.2785957, 0.2847609, 0.307846, 0.3507892, 0.5678833, 
    0.03814954, 0.2937672, 0.4104928, 0.4382154, 0.2964832,
  0.323549, 0.3626741, 0.3602288, 0.3169654, 0.3314413, 0.3288823, 0.2930083, 
    0.2389957, 0.293868, 0.2874243, 0.1984551, 0.1545118, 0.2565927, 
    0.2564549, 0.2496573, 0.3491749, 0.3273328, 0.3580758, 0.2973678, 
    0.2897524, 0.305464, 0.2639022, 0.2265659, 0.2534826, 0.2376199, 
    0.3443506, 0.3368826, 0.3941691, 0.3913909,
  0.3114451, 0.2803105, 0.3215148, 0.2324886, 0.2283981, 0.2165156, 
    0.2340538, 0.2102139, 0.273827, 0.2958359, 0.1980177, 0.2385878, 
    0.1345274, 0.2089042, 0.1740065, 0.222688, 0.1884352, 0.2063232, 
    0.1978309, 0.2139486, 0.2601862, 0.3170322, 0.25739, 0.1362432, 
    0.1069372, 0.2964391, 0.4112179, 0.3090347, 0.3264875,
  0.2043548, 0.07676321, 0.04451391, 0.1670846, 0.1565844, 0.1299154, 
    0.1590954, 0.1838382, 0.2199825, 0.1341663, 0.09873927, 0.02613809, 
    0.03215696, 0.1445362, 0.1941365, 0.1763561, 0.1715251, 0.06093305, 
    0.09184427, 0.1850656, 0.2086199, 0.2086771, 0.1856487, 0.1228955, 
    0.01393604, 0.06918866, 0.1310635, 0.1362593, 0.1972757,
  0.01931357, 0.03357694, 0.01427611, 0.07950684, 0.03601369, 0.01954149, 
    0.009405627, 0.04190674, 0.07493901, 0.07077405, -3.088168e-05, 
    1.374938e-07, 0.005145294, 0.02950788, 0.06297024, 0.04870317, 
    0.01586817, 0.06559024, 0.2226644, 0.08258975, 0.0809877, 0.008153956, 
    0.05753893, 0.03787535, 0.002932892, 0.07793276, 0.07973613, 0.01578169, 
    0.01301579,
  0.04929464, 0.02792577, 0.0153032, 0.007670495, 0.0003304522, 0.009398114, 
    0.01931498, 0.03362844, 0.06361987, -3.23408e-05, 6.874626e-07, 
    -1.551229e-06, 0.0119414, 0.00752876, 0.01172451, 0.01235384, 0.00670777, 
    0.03392106, 0.02078957, 0.00701283, 0.002434146, 0.007429564, 0.07302187, 
    0.05138989, 0.0106107, 0.1775519, 0.009464351, 0.001820847, 0.01683269,
  0.09895983, 0.05227622, 0.007887835, 0.2115089, 0.007853388, 0.01832165, 
    0.01080875, 0.002451021, 0.005556176, 0.001703741, 0.002146442, 
    0.002265018, 0.006518136, 0.0006561953, 0.002283665, 0.001093413, 
    4.263052e-05, 0.001942115, 0.0002790279, 0.0007691034, 0.004247221, 
    0.05663588, 0.1244322, 0.0006432925, 0.03436301, 0.03029876, 
    -0.0006292053, 0.003055971, 0.03000087,
  0.01931446, 0.05250202, 0.03059099, 0.1028831, 0.007697219, 0.008301613, 
    0.003663019, 0.009764723, 0.06368058, 0.06763232, 0.0007416282, 
    0.002347445, 0.001081299, 0.00416791, 0.002832753, 0.003956828, 
    0.003045466, 0.007883932, 0.008667747, 0.01251073, 0.03546165, 0.1402694, 
    0.1773345, 0.0083667, 0.003304534, 0.001102569, 0.03600126, 0.006603315, 
    0.05994035,
  -3.895192e-08, 1.42281e-08, 1.080657e-07, 0.0008082183, 0.05610488, 
    0.003310751, 0.001058866, 0.006641835, 0.002836039, 0.03095352, 
    0.01889413, 0.003060563, 0.008276075, 0.01055885, 0.0016211, 0.00147996, 
    0.01321588, 0.01230558, 0.01506174, 0.03104847, 0.03940419, 0.008084041, 
    0.2612039, 0.04757019, 0.0001300037, 0.0007435707, 0.00560136, 
    0.000989896, -5.959142e-07,
  2.339618e-09, 4.522732e-10, 1.75611e-10, -5.05948e-05, 4.714171e-10, 
    0.0006436962, 0.005499543, 0.0008730981, 0.02461558, 0.006470035, 
    0.01158068, 0.01061367, 0.003073824, 0.001960967, 0.002633674, 
    0.00261622, 0.01796561, 0.01750476, 0.03593565, 0.02028804, 0.001298712, 
    0.1463008, 0.002036839, -0.001103042, 0.004148854, 0.0001649661, 
    0.001359286, 0.0002111154, 1.649645e-08,
  -1.164727e-05, 0.006835156, 0.0004146276, 0.03999339, 0.03076922, 
    0.02450661, -0.002411692, -0.0002063385, 0.05965478, 0.02288541, 
    0.01090516, 0.01886185, 0.02899454, 0.05200683, 0.05022437, 0.02240509, 
    0.02855422, 0.004941582, 0.1205689, 0.05543095, 3.079837e-07, 0.06010853, 
    0.05192144, 0.009354752, 0.02094672, 0.03319098, 0.0009625164, 
    0.004078244, 0.01536055,
  0.001732468, 0.003986608, 0.05750415, 0.2041066, 0.004803929, 0.002985168, 
    0.1394125, 0.00368442, -0.0001050813, 0.01318327, 0.1501472, 0.02760769, 
    0.02951308, 0.04982381, 0.08080424, 0.1077632, 0.1713404, 0.1907534, 
    0.1253699, 0.2159621, 0.01003112, 0.1009657, 0.2075183, 0.04670457, 
    0.08947209, 0.1858568, 0.1833679, 0.03986439, 0.05281927,
  0.1060638, 0.4903232, 0.3831761, 0.3185098, 0.2246083, 0.1265077, 
    0.1128812, 0.1447555, 0.04562623, 0.2322908, 0.09720167, 0.4189672, 
    0.09609748, 0.1333433, 0.1675337, 0.2669264, 0.2891814, 0.2599498, 
    0.264796, 0.4661608, 0.1696316, 0.1935842, 0.283317, 0.5905146, 0.163002, 
    0.1715521, 0.1887502, 0.2768445, 0.1263983,
  0.1017804, 0.4901361, 0.4932744, 0.7491496, 0.6969321, 0.4250432, 
    0.6325284, 0.6323951, 0.5711485, 0.6013245, 0.6707497, 0.3332277, 
    0.2146092, 0.1826139, 0.3726513, 0.3096648, 0.398425, 0.2534183, 
    0.3740395, 0.5139278, 0.4801286, 0.1523198, 0.06469446, 0.1927644, 
    0.1014544, 0.1239896, 0.1793818, 0.1167291, 0.1378955,
  0.02358435, 0.03021229, 0.2147712, 0.07102003, 0.1708782, 0.3218745, 
    0.611321, 0.5366241, 0.4296468, 0.5136128, 0.5130088, 0.3196774, 
    0.4700543, 0.5698441, 0.539257, 0.4446353, 0.2989902, 0.3609577, 
    0.3913536, 0.4995718, 0.4302588, 0.5558775, 0.3436351, 0.4372693, 
    0.06486575, 0.3644278, 0.3651306, 0.1580739, 0.1041144,
  0.3075882, 0.3736488, 0.3322835, 0.3318104, 0.2605966, 0.4298922, 0.460425, 
    0.4772289, 0.535695, 0.6586843, 0.6438273, 0.6377575, 0.6140726, 
    0.6157522, 0.6267096, 0.5470589, 0.5364431, 0.5674938, 0.5942606, 
    0.4819578, 0.4681084, 0.2807662, 0.24542, 0.2970956, 0.2042596, 
    0.2630489, 0.143005, 0.3371067, 0.4881953,
  0.4127883, 0.414814, 0.4168397, 0.4188654, 0.4208911, 0.4229168, 0.4249425, 
    0.4016849, 0.4076956, 0.4137062, 0.4197169, 0.4257275, 0.4317382, 
    0.4377488, 0.4873905, 0.4823048, 0.4772191, 0.4721334, 0.4670476, 
    0.4619619, 0.4568762, 0.4587326, 0.455782, 0.4528313, 0.4498807, 0.44693, 
    0.4439794, 0.4410287, 0.4111677,
  0.2140058, 0.246437, 0.2259909, 0.1804231, 0.1971028, 0.2449581, 0.235091, 
    0.1716662, 0.1502536, 0.1468701, 0.1173892, 0.05743364, 0.1389379, 
    0.009327427, 0.1922057, 0.2756603, 0.2249177, 0.2344522, 0.1071596, 
    0.0685021, 0.2616222, 0.4631797, 0.2472521, 0.09800259, 0.059439, 
    0.13591, 0.04878904, 0.08383307, 0.1594933,
  0.1434044, 0.0884128, 0.114399, 0.07797365, 0.07419007, 0.2191636, 
    0.03748062, 0.07172877, 0.1075049, 0.1546649, 0.09792683, 0.06658691, 
    0.07586969, 0.08775714, 0.2213757, 0.3098991, 0.2415899, 0.2315165, 
    0.2677978, 0.217482, 0.2221571, 0.236754, 0.2892423, 0.495542, 0.0333971, 
    0.2942344, 0.3510537, 0.36798, 0.2776776,
  0.2787281, 0.2690485, 0.2817356, 0.2353678, 0.2610521, 0.2531181, 
    0.1948641, 0.1732876, 0.2232275, 0.2283027, 0.163645, 0.1335233, 
    0.2258959, 0.2097564, 0.1945267, 0.3059871, 0.2838161, 0.2932709, 
    0.2514552, 0.2642478, 0.2469268, 0.209112, 0.1754209, 0.1882799, 
    0.1970633, 0.3181189, 0.3434457, 0.3282299, 0.3084913,
  0.2712441, 0.2144227, 0.2444283, 0.1855851, 0.1806262, 0.1563962, 
    0.1918238, 0.1561546, 0.2249536, 0.2422262, 0.1612461, 0.199428, 
    0.08470345, 0.1558098, 0.166424, 0.1842518, 0.1246654, 0.1347645, 
    0.1423682, 0.1443186, 0.1842092, 0.2472347, 0.1963056, 0.1149712, 
    0.1102192, 0.2558643, 0.3544438, 0.2826194, 0.2999406,
  0.1601362, 0.04031239, 0.02686129, 0.141847, 0.1073365, 0.08480684, 
    0.1173338, 0.1392336, 0.160493, 0.08776867, 0.0617155, 0.01267801, 
    0.02157054, 0.1175134, 0.1636135, 0.1325152, 0.1342068, 0.04810959, 
    0.07066362, 0.1621031, 0.1773509, 0.1993548, 0.1391169, 0.1128797, 
    0.01686264, 0.06049817, 0.08502349, 0.100988, 0.14931,
  0.01120001, 0.01692363, 0.01431508, 0.04069874, 0.01406113, 0.009930032, 
    0.003515576, 0.02072681, 0.05576116, 0.04603102, -1.139475e-05, 
    1.247839e-07, 0.002955504, 0.01032505, 0.02892027, 0.03437053, 
    0.006165409, 0.03480492, 0.1561734, 0.06391059, 0.05525043, 0.003235301, 
    0.02720645, 0.03695155, 0.001327181, 0.03487327, 0.03678882, 0.005596324, 
    0.007530579,
  0.02357411, 0.0207553, 0.008792541, 0.00276688, -0.00224762, 0.002742548, 
    0.003805981, 0.007822151, 0.03135165, -2.049941e-05, 1.155484e-07, 
    -1.852931e-06, 0.005894318, 0.002510237, 0.003321, 0.006161028, 
    0.003256522, 0.01527414, 0.01091897, 0.006139997, 0.001265775, 
    0.003983439, 0.03679096, 0.02435665, 0.007529662, 0.1482594, 0.004419796, 
    0.00101777, 0.007350643,
  0.05466407, 0.02261104, 0.007135509, 0.1554541, 0.002907058, 0.006733575, 
    0.003783539, 0.0008490367, 0.002475307, 0.0009322412, 0.0006383684, 
    0.001149716, 0.001399548, 0.0001859232, 0.0008427455, 0.0003543544, 
    3.767353e-05, 0.001082959, 0.000142841, 0.0004415055, 0.002425641, 
    0.03059033, 0.06307516, 0.0002405526, 0.02939852, 0.02720601, 
    7.705991e-05, 0.001511384, 0.01526364,
  0.007926373, 0.05286001, 0.03068757, 0.08948504, 0.003928654, 0.004244463, 
    0.001857411, 0.00517462, 0.05085385, 0.06608209, 0.0002016249, 
    0.001108685, 0.0006050077, 0.001438541, 0.00180128, 0.001708754, 
    0.001604523, 0.003931042, 0.004186143, 0.005455745, 0.01450298, 
    0.06343291, 0.08941454, 0.01068249, 0.002371134, 0.0003693244, 0.0231439, 
    0.001884654, 0.03733729,
  2.597581e-09, 1.424294e-08, 1.215e-07, 0.0007078568, 0.03576827, 
    0.001335216, -0.0008161263, 0.001979896, 0.001020395, 0.01184518, 
    0.01026647, 0.001363686, 0.00316118, 0.004897934, 0.0004043194, 
    0.0003799591, 0.00801188, 0.004946533, 0.004258054, 0.01411001, 
    0.01691943, 0.002191062, 0.1777567, 0.04121268, 9.443087e-05, 
    0.0004261088, 0.002681102, 0.0006401737, -7.456889e-07,
  2.31868e-09, 4.425796e-10, 1.53116e-10, -3.322809e-06, 2.454618e-10, 
    0.0003363953, 0.004512944, 0.0005276615, 0.01859105, 0.003303637, 
    0.003752586, 0.004167844, 0.001143625, 0.0008935914, 0.001346909, 
    0.001589116, 0.006610657, 0.003741269, 0.01650537, 0.009445418, 
    0.0006734704, 0.1075132, 0.00102292, -0.000879339, 0.002221707, 
    8.748622e-05, 0.0008156027, 0.0001114617, 1.596374e-08,
  -2.391952e-05, 0.002043154, 9.695371e-05, 0.02754644, 0.01958708, 
    0.0152715, -0.002047626, 0.0002499162, 0.05188802, 0.02399503, 0.0072509, 
    0.01116385, 0.01538911, 0.03159122, 0.02623925, 0.009182957, 0.01316191, 
    0.002092089, 0.07146745, 0.03512431, 8.786442e-05, 0.05272321, 
    0.04100783, 0.004327061, 0.007721161, 0.01737298, 0.0005820098, 
    0.002359605, 0.01523432,
  0.001523828, 0.00234383, 0.03792952, 0.2004529, 0.001698921, 0.002264272, 
    0.1347755, 0.002058894, -8.948908e-05, 0.009026524, 0.1362133, 
    0.02086687, 0.02111527, 0.034232, 0.05889655, 0.08925734, 0.1449864, 
    0.1340296, 0.06988649, 0.204244, 0.00568722, 0.08574435, 0.1772477, 
    0.03783934, 0.05796393, 0.1370112, 0.1460132, 0.02121918, 0.03742182,
  0.062114, 0.4375241, 0.3303588, 0.2866333, 0.2173448, 0.0971083, 0.0910839, 
    0.1291133, 0.03135115, 0.1819918, 0.08612322, 0.3914265, 0.07276201, 
    0.09408729, 0.1268529, 0.2244545, 0.2284316, 0.2142717, 0.2202164, 
    0.4526323, 0.1522341, 0.1484471, 0.2111991, 0.5321671, 0.1348862, 
    0.145126, 0.1613846, 0.2256862, 0.09056941,
  0.06785385, 0.4935292, 0.4309605, 0.7234359, 0.6328428, 0.4347438, 
    0.5658559, 0.5443452, 0.5463917, 0.5051931, 0.5972292, 0.3425935, 
    0.222115, 0.2079368, 0.3176639, 0.2652479, 0.3972183, 0.1996963, 
    0.3160067, 0.4578656, 0.4831883, 0.1539973, 0.04683051, 0.2766177, 
    0.07521521, 0.09746422, 0.1367882, 0.08342993, 0.1038624,
  0.01458973, 0.01619884, 0.2082052, 0.04871381, 0.1246141, 0.2644872, 
    0.5149181, 0.3823171, 0.381653, 0.5005724, 0.5908694, 0.3006121, 
    0.6091806, 0.4766137, 0.5006526, 0.4315272, 0.2641059, 0.3198583, 
    0.3788939, 0.4261814, 0.4013315, 0.5705905, 0.3217459, 0.5019408, 
    0.04352728, 0.3035935, 0.3891034, 0.1204221, 0.08152425,
  0.4132145, 0.3558432, 0.4110469, 0.3897379, 0.3386411, 0.4910962, 
    0.5743687, 0.6305922, 0.6520711, 0.7719043, 0.7752227, 0.7319165, 
    0.6912385, 0.6518243, 0.6441029, 0.5506772, 0.5678463, 0.6965006, 
    0.6371536, 0.578675, 0.6337523, 0.3357648, 0.3103237, 0.4608861, 
    0.1711249, 0.2565235, 0.1227776, 0.3298752, 0.5316507,
  0.3317362, 0.3338371, 0.3359379, 0.3380388, 0.3401396, 0.3422405, 
    0.3443413, 0.3222352, 0.3242894, 0.3263436, 0.3283977, 0.3304519, 
    0.3325061, 0.3345602, 0.3757909, 0.3750784, 0.3743659, 0.3736534, 
    0.372941, 0.3722285, 0.371516, 0.373624, 0.3701814, 0.3667389, 0.3632964, 
    0.3598538, 0.3564112, 0.3529687, 0.3300555,
  0.1811901, 0.2120274, 0.1849269, 0.1444577, 0.1490198, 0.2069603, 
    0.1945575, 0.1664332, 0.1086778, 0.09932268, 0.06495006, 0.02988788, 
    0.08877642, 0.007097545, 0.1822261, 0.2684184, 0.164248, 0.2041895, 
    0.08686376, 0.06847474, 0.1973357, 0.4023497, 0.2125222, 0.07282231, 
    0.04811464, 0.1237062, 0.03221113, 0.06852052, 0.1488611,
  0.1220047, 0.07342387, 0.09398966, 0.06422576, 0.0520571, 0.1838402, 
    0.0304527, 0.05311061, 0.0835318, 0.1104748, 0.08128544, 0.04794316, 
    0.05777468, 0.0786055, 0.1964472, 0.2590971, 0.1884999, 0.1873961, 
    0.199924, 0.1576307, 0.1617021, 0.1812382, 0.2307855, 0.4122415, 
    0.02925472, 0.2500883, 0.2814398, 0.2757672, 0.2453832,
  0.2087282, 0.1898852, 0.2050371, 0.1768205, 0.1981985, 0.1860026, 
    0.1380264, 0.1216766, 0.1612806, 0.1725648, 0.1252676, 0.1068202, 
    0.1908892, 0.1618722, 0.1454088, 0.2502393, 0.2396284, 0.237237, 
    0.2078747, 0.2170499, 0.1857041, 0.1490314, 0.1219334, 0.1268333, 
    0.1639124, 0.2603096, 0.2971797, 0.2473302, 0.2322675,
  0.2203585, 0.1627029, 0.1885779, 0.1381796, 0.13623, 0.1173129, 0.1426535, 
    0.1093147, 0.1635088, 0.1797121, 0.1109072, 0.1370138, 0.04965702, 
    0.1162091, 0.1403665, 0.1293943, 0.07077524, 0.08977742, 0.1083149, 
    0.09451848, 0.1208966, 0.1738492, 0.1272839, 0.09454156, 0.1035427, 
    0.2030031, 0.2955379, 0.2320923, 0.2410497,
  0.1091744, 0.0219832, 0.01580788, 0.1012924, 0.07162191, 0.05616877, 
    0.07691374, 0.09586732, 0.101374, 0.05168164, 0.03969165, 0.008613749, 
    0.01684026, 0.09165565, 0.1340511, 0.07956904, 0.1042949, 0.03145353, 
    0.04656125, 0.1309225, 0.1303197, 0.1650413, 0.08167251, 0.1060399, 
    0.03378261, 0.0484807, 0.05217548, 0.06651738, 0.1046017,
  0.007815037, 0.00956579, 0.01022184, 0.01662805, 0.007548553, 0.005707663, 
    0.002201453, 0.01072341, 0.03466439, 0.03486323, -6.35701e-06, 
    1.21585e-07, 0.00152882, 0.004138004, 0.01297369, 0.02410479, 
    0.002585423, 0.01795522, 0.09440561, 0.04433909, 0.03455496, 0.00185197, 
    0.01475375, 0.03153628, 0.0006989131, 0.01493005, 0.01699873, 
    0.002915483, 0.005199483,
  0.01419819, 0.02508267, 0.005204364, 0.001601918, -0.001744806, 
    0.001167257, 0.001426114, 0.003483733, 0.01854024, -1.461452e-05, 
    9.729509e-08, -4.176077e-06, 0.003750941, 0.0008570042, 0.001098245, 
    0.002995997, 0.001790888, 0.006661356, 0.003660391, 0.004038022, 
    0.0007942562, 0.002545319, 0.02270026, 0.01551995, 0.004335137, 
    0.1131705, 0.001674213, 0.0006687153, 0.00416371,
  0.03544973, 0.01362001, 0.006074222, 0.1186035, 0.001634275, 0.002621628, 
    0.001474571, 0.0004302745, 0.001523373, 0.000684838, 0.0003412381, 
    0.0007061495, 0.0005189959, 0.0001163732, 0.0005097452, 0.0001945054, 
    5.973927e-05, 0.0007264625, 9.111212e-05, 0.0002948873, 0.001621415, 
    0.01996451, 0.03979694, 0.0002502216, 0.02223168, 0.02328855, 
    0.0002456192, 0.000922601, 0.009708356,
  0.003126702, 0.05090528, 0.0280803, 0.07413003, 0.002470881, 0.001778566, 
    0.001148943, 0.003311533, 0.04622107, 0.06892436, 0.0001058088, 
    0.0006523953, 0.0003998791, 0.0005049008, 0.0009495192, 0.0008519444, 
    0.001030296, 0.002513414, 0.002585596, 0.003120987, 0.008338938, 
    0.03736425, 0.05385488, 0.01207083, 0.003080563, 0.0001590586, 
    0.01056447, 0.0006453387, 0.01499211,
  -2.442463e-09, 1.391216e-08, 1.215609e-07, 0.0009911669, 0.02209075, 
    0.0007435183, -0.0005025406, 0.0006749653, 0.000648439, 0.004243977, 
    0.004494517, 0.0005829836, 0.001274172, 0.00196806, 0.0001424661, 
    0.0002261341, 0.004179541, 0.001813483, 0.001981952, 0.005706262, 
    0.006430158, 0.0009198869, 0.1161521, 0.03890975, 6.944803e-05, 
    0.0002866317, 0.00133765, 0.0004646813, -3.58511e-06,
  2.330673e-09, 4.39712e-10, 1.502775e-10, 7.675319e-06, 7.484262e-11, 
    0.0002153494, 0.002554063, 0.0003568213, 0.01477132, 0.002091719, 
    0.001463192, 0.00180242, 0.0006847776, 0.0005701149, 0.00085299, 
    0.001110076, 0.003290387, 0.001687195, 0.009799848, 0.005461418, 
    0.0004185534, 0.078638, 0.0006599686, -0.0007254923, 0.001444292, 
    5.574408e-05, 0.0005629887, 4.986719e-05, 1.604054e-08,
  -2.840689e-05, 0.00107936, 5.723722e-05, 0.01861803, 0.01423549, 
    0.01052734, -0.001445618, 0.00159473, 0.04346035, 0.01554215, 
    0.005467241, 0.006011356, 0.007462247, 0.01214906, 0.01169283, 
    0.003728736, 0.005566779, 0.001148499, 0.03550798, 0.02486576, 
    4.208795e-05, 0.04742836, 0.03707266, 0.00236587, 0.003041924, 
    0.008178106, 0.0004072285, 0.001693661, 0.01127198,
  3.400003e-05, 0.001474924, 0.0235546, 0.1874285, 0.0005815231, 0.001554573, 
    0.1089797, 0.001301875, -6.051507e-05, 0.007024362, 0.119396, 0.01611614, 
    0.01324808, 0.01872634, 0.0410648, 0.06754721, 0.1064415, 0.08794883, 
    0.03572475, 0.1891567, 0.003651903, 0.07814383, 0.1517299, 0.02983191, 
    0.03305884, 0.08439438, 0.09588452, 0.01286426, 0.02559941,
  0.04036857, 0.3728012, 0.2692954, 0.2279382, 0.1858898, 0.0851266, 
    0.07273404, 0.1098437, 0.0255674, 0.1532087, 0.0738226, 0.357989, 
    0.05656045, 0.066771, 0.09568033, 0.1643606, 0.1633608, 0.1574567, 
    0.1565278, 0.4329779, 0.1279986, 0.1130377, 0.1554543, 0.4506243, 
    0.1168911, 0.1225263, 0.1237329, 0.1565592, 0.06036049,
  0.04415944, 0.4809608, 0.3756512, 0.6676672, 0.5829822, 0.4143124, 
    0.5037671, 0.4561059, 0.4802217, 0.4010018, 0.4783987, 0.361016, 
    0.2597158, 0.1964076, 0.2722749, 0.19504, 0.4011025, 0.1556393, 
    0.2705441, 0.4030527, 0.4834015, 0.1437615, 0.03686491, 0.3672974, 
    0.05954757, 0.07552028, 0.09310447, 0.05704212, 0.0715974,
  0.009141282, 0.009809709, 0.2499427, 0.03500849, 0.09494963, 0.2220268, 
    0.4117711, 0.297027, 0.3397084, 0.4581837, 0.564373, 0.2634797, 
    0.6113234, 0.3438965, 0.4177392, 0.3826371, 0.2563945, 0.2251493, 
    0.3362407, 0.2892691, 0.2489286, 0.5678121, 0.2823124, 0.5505467, 
    0.03266223, 0.258879, 0.4223728, 0.09894332, 0.06267633,
  0.4669666, 0.3534895, 0.4178936, 0.4169466, 0.3997028, 0.4376409, 
    0.5086269, 0.6170336, 0.6065075, 0.6520078, 0.7538911, 0.6830527, 
    0.6028914, 0.5635337, 0.4956677, 0.579951, 0.4992922, 0.6004237, 
    0.545476, 0.6303423, 0.6760437, 0.4068555, 0.3852399, 0.5654306, 
    0.1478294, 0.2462625, 0.1135895, 0.3261948, 0.5880356,
  0.2489596, 0.2506604, 0.2523612, 0.254062, 0.2557628, 0.2574637, 0.2591645, 
    0.1996907, 0.2018568, 0.2040229, 0.2061889, 0.208355, 0.2105211, 
    0.2126871, 0.2813494, 0.2801784, 0.2790075, 0.2778365, 0.2766656, 
    0.2754947, 0.2743237, 0.261058, 0.2583621, 0.2556661, 0.2529702, 
    0.2502742, 0.2475783, 0.2448824, 0.2475989,
  0.1539144, 0.1544172, 0.1326471, 0.1172955, 0.1237794, 0.173463, 0.1418875, 
    0.1231891, 0.0691141, 0.06111557, 0.04226924, 0.01983159, 0.06388848, 
    0.005785978, 0.1847758, 0.2381821, 0.1502228, 0.1834436, 0.07222874, 
    0.0688851, 0.1619631, 0.3456391, 0.178805, 0.06402224, 0.07335512, 
    0.1271794, 0.02566146, 0.05625438, 0.1394448,
  0.1285983, 0.07038135, 0.09504692, 0.05653654, 0.04184255, 0.1576501, 
    0.02511447, 0.04232109, 0.06920491, 0.08282632, 0.06909844, 0.03966836, 
    0.04716026, 0.07045451, 0.1751366, 0.2132774, 0.1498966, 0.1625073, 
    0.1596316, 0.1266736, 0.1257629, 0.1408838, 0.1856661, 0.3440416, 
    0.02141116, 0.202811, 0.237445, 0.219412, 0.2054087,
  0.1649601, 0.1491921, 0.1621951, 0.1419945, 0.1582251, 0.1477244, 
    0.1075349, 0.09294504, 0.1248724, 0.1383907, 0.1037652, 0.08615552, 
    0.1642104, 0.1309491, 0.113958, 0.2094213, 0.2109629, 0.2070462, 
    0.1760645, 0.1755998, 0.1453886, 0.1145043, 0.08687355, 0.09114884, 
    0.1336307, 0.2075147, 0.251079, 0.1947215, 0.180325,
  0.1833108, 0.1289553, 0.1501157, 0.1096608, 0.1081424, 0.09835371, 
    0.1081783, 0.08208673, 0.1223877, 0.1388387, 0.08183777, 0.09446114, 
    0.03224682, 0.08383925, 0.1043156, 0.09169386, 0.04772945, 0.06091061, 
    0.07599609, 0.064191, 0.0839391, 0.1307674, 0.08501166, 0.08202973, 
    0.07488639, 0.1591166, 0.2457871, 0.1819878, 0.1955725,
  0.07286772, 0.01440184, 0.009656932, 0.06373968, 0.04425314, 0.03680794, 
    0.04762743, 0.06753242, 0.06961811, 0.03061231, 0.02461855, 0.006502766, 
    0.01240788, 0.06279389, 0.1167718, 0.05097032, 0.08625552, 0.0170856, 
    0.02518014, 0.1072172, 0.09278627, 0.1210998, 0.05208841, 0.09214462, 
    0.03873559, 0.03522099, 0.03407518, 0.0476534, 0.07387426,
  0.006085237, 0.006862352, 0.007423424, 0.00898893, 0.00403291, 0.003717601, 
    0.001711764, 0.006620709, 0.02543543, 0.02790362, -4.087125e-06, 
    1.201131e-07, 0.000990079, 0.002253019, 0.00642035, 0.01405859, 
    0.001604621, 0.009947934, 0.0575651, 0.02667268, 0.01861976, 0.001372516, 
    0.009878031, 0.02668343, 0.000336987, 0.008420452, 0.008955187, 
    0.002060033, 0.00402552,
  0.01000494, 0.0189436, 0.002773868, 0.001131186, -0.001352568, 
    0.0005493365, 0.0009425912, 0.00241339, 0.01316873, -1.146689e-05, 
    9.244697e-08, -7.42278e-07, 0.002757803, 0.000501933, 0.000618365, 
    0.001491242, 0.001121421, 0.003360432, 0.001879408, 0.001904173, 
    0.0005732007, 0.001861054, 0.01610013, 0.01157966, 0.003032183, 
    0.08636276, 0.0009481774, 0.000498968, 0.002809224,
  0.02631986, 0.009899369, 0.008066613, 0.1068855, 0.001127952, 0.001113792, 
    0.0006561285, 0.0003018278, 0.001089604, 0.0005208849, 0.0002402908, 
    0.000490209, 0.000397071, 9.242454e-05, 0.000376322, 0.0001463345, 
    5.776671e-05, 0.0005477958, 6.702007e-05, 0.0002209104, 0.001221607, 
    0.01480228, 0.02888278, 0.001275515, 0.01763798, 0.01766313, 
    0.0002448242, 0.0006614884, 0.007111808,
  0.001381556, 0.04306282, 0.01766477, 0.0621331, 0.001777389, 0.001022074, 
    0.0008190499, 0.002407548, 0.05141039, 0.07409551, 7.235947e-05, 
    0.0004546155, 0.0002950621, 0.0003041939, 0.0006355855, 0.0005357549, 
    0.0007547629, 0.001838985, 0.001858095, 0.002124569, 0.005699448, 
    0.02620856, 0.03804896, 0.009418686, 0.003553767, 0.0001005691, 
    0.004822998, 0.0002758232, 0.00573687,
  -1.572225e-07, 1.317056e-08, 1.202342e-07, 0.001360362, 0.01428162, 
    0.0005276703, -3.216953e-05, 0.0003240805, 0.0004493249, 0.001764202, 
    0.002034268, 0.0003332336, 0.0006262471, 0.001018888, 9.799487e-05, 
    0.0001588731, 0.002051815, 0.0009742034, 0.001268709, 0.002403946, 
    0.002783121, 0.0004978416, 0.08113284, 0.03433961, 5.415573e-05, 
    0.0002163312, 0.0008446035, 0.0003689684, -3.987687e-05,
  2.339359e-09, 4.378146e-10, 1.524752e-10, 9.770441e-06, 9.9205e-11, 
    0.0001641172, 0.001484608, 0.0002712492, 0.01228397, 0.001524896, 
    0.0007833514, 0.001068969, 0.0004865652, 0.0004193992, 0.000619388, 
    0.0008568455, 0.001848079, 0.001082562, 0.006930317, 0.00399043, 
    0.0003076049, 0.06639048, 0.0005032998, -0.0006781846, 0.001063251, 
    4.051224e-05, 0.0004312519, 3.585303e-05, 1.611939e-08,
  -2.388995e-05, 0.0007113132, 4.118556e-05, 0.0161809, 0.01090466, 
    0.006559799, -0.001358028, 0.002641437, 0.04417255, 0.0123157, 
    0.004532157, 0.003670075, 0.00422495, 0.00567262, 0.004928783, 
    0.001955811, 0.003068018, 0.0006851924, 0.01855562, 0.01755504, 
    2.487373e-05, 0.04690025, 0.03578707, 0.001797982, 0.001678045, 
    0.003883619, 0.0003158036, 0.001342369, 0.008822392,
  -0.0006034427, 0.0009572448, 0.01531484, 0.1718848, 0.0002152802, 
    0.001060282, 0.1020183, 0.0009682994, -3.997116e-05, 0.005378088, 
    0.1118319, 0.01381594, 0.00719609, 0.01133254, 0.02586892, 0.04638734, 
    0.07611898, 0.05389514, 0.02072774, 0.1716828, 0.002435167, 0.0738057, 
    0.1341617, 0.0239492, 0.01953506, 0.04934634, 0.04974141, 0.008830547, 
    0.01939169,
  0.02889084, 0.3247288, 0.234508, 0.1879313, 0.15991, 0.07467377, 
    0.06441922, 0.1024068, 0.0289464, 0.1336551, 0.0677, 0.3469793, 
    0.04718477, 0.05318579, 0.07346266, 0.118849, 0.1178601, 0.1083376, 
    0.1123585, 0.417657, 0.1103914, 0.0874367, 0.1319844, 0.3925728, 
    0.1010657, 0.1101653, 0.09836097, 0.1079044, 0.04038014,
  0.03170525, 0.4436163, 0.3395086, 0.5975829, 0.5486578, 0.3845714, 
    0.4581301, 0.4044352, 0.4319187, 0.3219519, 0.3824996, 0.3925282, 
    0.2916677, 0.19999, 0.2331314, 0.1514033, 0.3947722, 0.1333901, 
    0.2391674, 0.3601149, 0.440478, 0.1326617, 0.03095961, 0.4420975, 
    0.04958474, 0.06261083, 0.070648, 0.04059928, 0.05251424,
  0.006337594, 0.007231047, 0.313353, 0.02714957, 0.07740255, 0.1755107, 
    0.346922, 0.2564588, 0.3380905, 0.4207843, 0.5500315, 0.2323039, 
    0.5298117, 0.2564288, 0.3454064, 0.3346179, 0.2374634, 0.1766451, 
    0.2457068, 0.1959069, 0.1207425, 0.4721346, 0.2681713, 0.5788395, 
    0.02652248, 0.2332639, 0.4650537, 0.07476665, 0.04967254,
  0.5137824, 0.3507872, 0.3707074, 0.3743837, 0.3704659, 0.3280808, 
    0.3902226, 0.4917314, 0.453281, 0.4575258, 0.5580782, 0.4462645, 
    0.4150782, 0.3646805, 0.3084046, 0.374893, 0.3914826, 0.4489671, 
    0.341489, 0.3692313, 0.4516852, 0.4167303, 0.4215328, 0.6617968, 
    0.1468384, 0.2034596, 0.1319584, 0.3077993, 0.527003,
  0.1813499, 0.1831295, 0.1849092, 0.1866888, 0.1884685, 0.1902481, 
    0.1920278, 0.1548532, 0.1560352, 0.1572172, 0.1583993, 0.1595813, 
    0.1607633, 0.1619453, 0.2071797, 0.2073352, 0.2074908, 0.2076463, 
    0.2078019, 0.2079574, 0.208113, 0.208149, 0.2050318, 0.2019146, 
    0.1987974, 0.1956801, 0.1925629, 0.1894457, 0.1799262,
  0.1586418, 0.1348162, 0.1043484, 0.1065873, 0.1126882, 0.1191175, 0.12288, 
    0.107506, 0.05603532, 0.04261462, 0.02975385, 0.01652538, 0.04880624, 
    0.005892667, 0.1971772, 0.2246817, 0.1644235, 0.1816061, 0.06806782, 
    0.07894631, 0.1495686, 0.3017095, 0.1561673, 0.07130957, 0.103465, 
    0.1252578, 0.0413298, 0.05045158, 0.1300971,
  0.1307728, 0.09598554, 0.1233671, 0.05023044, 0.0423483, 0.1431593, 
    0.02551841, 0.03867727, 0.06307673, 0.07466172, 0.06035016, 0.04314186, 
    0.04385073, 0.062776, 0.1685922, 0.1942042, 0.1304832, 0.1488687, 
    0.1423627, 0.1047725, 0.1102221, 0.1205417, 0.1660245, 0.3074568, 
    0.01556813, 0.177949, 0.2135187, 0.1902886, 0.1800233,
  0.1465744, 0.13429, 0.143785, 0.1253604, 0.1363721, 0.1268577, 0.09291448, 
    0.0796513, 0.1074332, 0.1219852, 0.09166142, 0.0769619, 0.1403826, 
    0.1138418, 0.09655331, 0.1827511, 0.1876424, 0.1815162, 0.154702, 
    0.1469708, 0.1232272, 0.09694038, 0.07018814, 0.07336731, 0.1067227, 
    0.1774699, 0.226166, 0.1706431, 0.1573104,
  0.1592044, 0.1115877, 0.1231035, 0.09162292, 0.09465764, 0.08343576, 
    0.08742697, 0.06918432, 0.09877645, 0.1156507, 0.06668279, 0.07016994, 
    0.02212466, 0.06538364, 0.08324782, 0.07220766, 0.03716738, 0.0477849, 
    0.0551502, 0.04716752, 0.06611803, 0.09984969, 0.06412186, 0.08313861, 
    0.0518841, 0.1222623, 0.2120318, 0.154039, 0.1703373,
  0.05548621, 0.01121226, 0.006178729, 0.04309183, 0.0305182, 0.02502617, 
    0.0325358, 0.0522298, 0.04690819, 0.02189146, 0.0177312, 0.005513864, 
    0.009217392, 0.04486251, 0.1352336, 0.03503748, 0.06206986, 0.01055479, 
    0.01627195, 0.08233625, 0.06928523, 0.08976384, 0.03586652, 0.08553011, 
    0.035173, 0.02541747, 0.02452898, 0.03639366, 0.05497119,
  0.005182929, 0.00568413, 0.01274402, 0.005953159, 0.002537822, 0.002805896, 
    0.001476975, 0.00464414, 0.01669008, 0.02381708, -2.81767e-06, 1.215e-07, 
    0.003442337, 0.001603798, 0.003576051, 0.008481424, 0.001243078, 
    0.006846115, 0.03674944, 0.01747012, 0.01070318, 0.001147011, 
    0.007962234, 0.02391252, -0.000247201, 0.005119361, 0.005331198, 
    0.001709241, 0.00335041,
  0.008122618, 0.01400778, 0.001616393, 0.0008912742, -0.001236637, 
    0.0003820748, 0.0007456269, 0.001918885, 0.01057515, -9.769647e-06, 
    9.178432e-08, -1.395922e-07, 0.002237407, 0.0004078779, 0.0004661307, 
    0.001003618, 0.0008671531, 0.002329554, 0.001303005, 0.001111343, 
    0.0004715115, 0.001551284, 0.0130758, 0.00933652, 0.01192492, 0.1052531, 
    0.0007188805, 0.0004188545, 0.002242209,
  0.02173591, 0.007977506, 0.03173296, 0.1654782, 0.0008953186, 0.0006800298, 
    0.0004142199, 0.0002524857, 0.0008858068, 0.0003256148, 0.0001937773, 
    0.0003903272, 0.0002173713, 7.920723e-05, 0.0003072706, 0.0001218469, 
    5.140273e-05, 0.0004555322, 5.559329e-05, 0.000185802, 0.001032265, 
    0.01229255, 0.02357777, 0.04245, 0.03464999, 0.01428191, 0.000220079, 
    0.0005453854, 0.005868686,
  0.0009150859, 0.0678597, 0.01946687, 0.06088526, 0.00142509, 0.0007345955, 
    0.0006561785, 0.00197302, 0.07389142, 0.1027427, 5.876864e-05, 
    0.0003604226, 0.0002425173, 0.0002304121, 0.0004939193, 0.0004318314, 
    0.0006218118, 0.001509099, 0.001500761, 0.001677486, 0.004530319, 
    0.02091607, 0.0304974, 0.04457462, 0.04584565, 7.907913e-05, 0.002884903, 
    0.0001763686, 0.003072815,
  -4.063821e-06, 1.248378e-08, 1.190533e-07, 0.001805328, 0.009309293, 
    0.0004243699, -0.000739989, 0.0002081719, -0.0002957229, 0.00114293, 
    0.001183313, 0.0002461641, 0.0004232763, 0.0007158603, 8.4164e-05, 
    0.0001309333, 0.001291685, 0.0007395628, 0.001013599, 0.001427589, 
    0.00178959, 0.0003506522, 0.1175739, 0.03073238, 4.598422e-05, 
    0.0001848901, 0.0006668985, 0.000317267, -0.0001632401,
  2.365534e-09, 4.498034e-10, 1.545699e-10, 1.032759e-05, -1.521605e-10, 
    0.0001333062, 0.0009674032, 0.0001403395, 0.01155433, 0.0009891267, 
    0.000592983, 0.0008323219, 0.0004000512, 0.0003461925, 0.0005063989, 
    0.0007241498, 0.001319964, 0.0008589158, 0.005605675, 0.003241813, 
    0.000252133, 0.06240557, 0.0004262424, -0.001214487, 0.0008665558, 
    3.368974e-05, 0.0003631287, 2.981562e-05, 1.616011e-08,
  -2.034791e-05, 0.000542652, 2.908325e-05, 0.01688738, 0.009382823, 
    0.007364349, 0.002126289, 0.006216832, 0.0484251, 0.01414673, 
    0.004046243, 0.002747744, 0.003062237, 0.003691419, 0.002805159, 
    0.001354025, 0.002240982, 0.0005269019, 0.01105515, 0.01299187, 
    2.292945e-05, 0.05439075, 0.04987023, 0.001546314, 0.001239954, 
    0.002631459, 0.0002669546, 0.001162766, 0.007407289,
  -0.00066071, 0.0003118058, 0.01078418, 0.1707996, 6.93877e-05, 
    0.0009037506, 0.09766417, 0.0007951796, -4.236258e-05, 0.004459408, 
    0.1294026, 0.01268238, 0.005066723, 0.008757588, 0.01971849, 0.03377295, 
    0.05636768, 0.03814795, 0.01412272, 0.16446, 0.001567695, 0.07213109, 
    0.1429432, 0.02011175, 0.01405773, 0.03378465, 0.02612406, 0.006998634, 
    0.01533746,
  0.02205956, 0.3218327, 0.2275557, 0.1952733, 0.1524279, 0.07688622, 
    0.06207479, 0.149219, 0.04661161, 0.1341867, 0.07812986, 0.3653969, 
    0.04244302, 0.04701068, 0.061163, 0.0943611, 0.09085125, 0.08177064, 
    0.08409945, 0.4426464, 0.1035246, 0.08322184, 0.1475664, 0.3931865, 
    0.09569433, 0.09691222, 0.08162436, 0.08491144, 0.02940738,
  0.02530765, 0.4518122, 0.3306076, 0.5742278, 0.5385363, 0.416503, 
    0.4629163, 0.4411611, 0.407136, 0.3083734, 0.3659516, 0.5147193, 0.39884, 
    0.2391496, 0.211391, 0.1284694, 0.4039769, 0.1261082, 0.266546, 
    0.3605201, 0.4345985, 0.1372162, 0.02855494, 0.5142668, 0.0445916, 
    0.05823524, 0.05976703, 0.03267788, 0.04382033,
  0.005140182, 0.005983995, 0.3798505, 0.02217917, 0.06788251, 0.1478942, 
    0.3196924, 0.258207, 0.3695073, 0.4295094, 0.6348248, 0.2488232, 
    0.4966646, 0.2266245, 0.3101412, 0.3127867, 0.2874792, 0.1580168, 
    0.2034519, 0.164945, 0.08794084, 0.4124655, 0.2487312, 0.5792084, 
    0.02324706, 0.2060239, 0.5128065, 0.06428698, 0.04213929,
  0.510744, 0.3507338, 0.3153281, 0.2598468, 0.3049161, 0.2778263, 0.2928402, 
    0.362324, 0.3289547, 0.3467885, 0.3792824, 0.3232245, 0.2946204, 
    0.2653522, 0.1860225, 0.2565001, 0.2856493, 0.3339429, 0.2572493, 
    0.2614388, 0.3183643, 0.4465349, 0.4856873, 0.713137, 0.1479894, 
    0.1929189, 0.1621467, 0.3130035, 0.4527495,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -1.138217e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -9.800518e-06, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -7.861276e-05, 0, 0, 0, 0,
  0, 0, 0, 0, -3.968773e-05, 0, 0, -1.970874e-05, 0, 0, 0, -5.643685e-05, 0, 
    0, 0.0001423138, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.349031e-05, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.495598e-05, -5.296782e-05, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.03109e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, -8.669944e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, -0.0001042122, 0, 0, 0, 0,
  0, 0, 0, 0, 0.0002039013, -1.20493e-05, -6.67663e-05, 0.002017465, 0, 0, 0, 
    0.0001826574, 0, -6.58538e-05, 4.883245e-05, 0, 0, 0, 0, 0, 0, 0, 0, 
    -1.748106e-05, 0.001791876, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 1.023877e-05, 0, 0, -5.306335e-07, 3.800426e-07, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5.444454e-05, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0.0003180573, 0, -3.717382e-10, 0, -9.593207e-06, 
    -9.79173e-05, -0.000158926, 0, 0, -6.959645e-06, 0, 0, -8.570663e-06, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002263848, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, -7.11349e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -4.78243e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, -0.000124516, 0, 0, 0, 0,
  0, 0, 0, 0, 0.0003656518, -4.329636e-05, -0.0003260972, 0.003231867, 0, 0, 
    4.972727e-06, 0.000913957, -2.840341e-05, 0.0003223257, 0.0006352871, 0, 
    0, 0, 0, 0, 0, 0, 0, -4.492389e-05, 0.004266388, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -3.428287e-05, 0.0002703622, 0, 0.002583209, 
    9.347022e-06, 0, 1.743166e-05, 0.001649699, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.001295727, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, -1.460231e-05, 0, 0, 0.004300561, 0.0001924297, 
    0.0002541722, -1.530014e-05, 0.0008731049, 0.000146523, -0.0002943696, 0, 
    0, 0.0001398146, -9.616686e-06, -2.285905e-05, -0.0001309318, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.00232332, -1.800154e-06, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, -1.214445e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, -2.660912e-10, 0, 0, 0,
  0, 0, 0, -9.339372e-05, 0, 7.966156e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0004188342, 0, 0.0001773836, 0, 0, 0, 0, 0, 0, 0, 0.0002432774, 0, 0, 0,
  0, 0, -7.919301e-05, 0, 0, 0, 0, 0, 0, 0, -1.85207e-05, 0, 0, 0, 0, 
    -7.597961e-06, 0, 0, 0, 0, 0, 0, 0, 0, 9.657419e-05, -1.649546e-05, 0, 0, 0,
  0, 0, 0, 0, 0.0004747432, -0.0001429544, -0.0002666366, 0.009351225, 0, 0, 
    9.870407e-06, 0.003311473, -0.0001022228, 0.001677625, 0.001043952, 
    -1.16587e-05, 0, 0, 0, 0, 0, 0, 0, -8.394045e-05, 0.006889476, 
    -4.006245e-06, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -4.436074e-06, 0.0007437892, 0, 0.006005459, 
    3.738809e-05, 0, 1.250111e-06, 0.007848411, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.004867509, 0, 0.0003906774, 0, 0, 0,
  0, 0, 0, 0, 0, -2.776785e-05, 0, 0, 0.006934865, 0.0007196103, 0.001173193, 
    -5.057141e-05, 0.004952475, 0.00191588, -0.0005644193, -5.232961e-05, 0, 
    0.001378585, -7.493592e-05, 0.0001051466, 0.0009127792, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.004888728, -1.939473e-05, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, -6.040682e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001377684, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0.001736352, 0, 0, 3.835647e-05, 0, 0, 0, 0, -5.244031e-05, 
    -4.291651e-05, 0, 0, 0, 0, 0, 0, -1.14269e-05, 0, 0, 0, 0, 0, 
    -8.749917e-06, 0.0001970587, 0, 0,
  0, 0, 0, -0.0001731127, 0, 0.004018475, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.001900905, 0, 0.006928907, -8.678668e-07, 0, 0, 0, 0, 0, -1.32705e-07, 
    0.002370973, 0.001592232, 0, 0,
  0, 0, 0.0004437942, 0, -3.377904e-05, 0, 0, 0, 0, 0, -4.63018e-05, 0, 0, 0, 
    0, -6.433963e-05, -3.461228e-05, 0.001151135, 0, 0, 0, 0, 0, 0, 
    0.0004442191, -0.0001506523, 0, 0, 0,
  0, 0, 5.067841e-05, -5.243139e-05, 0.007710775, 0.0004622182, 0.00167541, 
    0.01524097, 0, 0, 5.03033e-06, 0.004603947, -0.0001619995, 0.005908675, 
    0.002903094, 0.001981474, 0, 0, 0, 0, 0, 0, 0, 0.0007162479, 0.008223492, 
    0.0004203765, 0, 0, 0,
  0, 0, 0, 0, 0, 3.318413e-08, 0.001240183, 0.001832125, 5.617326e-07, 
    0.01424398, 0.0009918333, -2.456337e-05, 0.0003514473, 0.01301832, 0, 0, 
    0, -2.766062e-05, 0, 0, 0, 0, 0, 0.008935836, 0, 0.0005464507, 0, 0, 0,
  0, 0, 0, 0, 0, -5.030401e-05, 0, 0, 0.01123292, 0.007368704, 0.002025295, 
    -9.373123e-05, 0.01152965, 0.004451317, -0.0008578038, -0.0001046592, 0, 
    0.002941489, -0.000191754, 0.002362273, 0.003507652, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.006323283, -0.0001237662, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, -1.208136e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -4.911345e-07, 0, 0, 0, 0, 0, 0, 0, -3.340078e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0.002716417, 0, 0, 0, 0, 0, 0, 0, 0.003496203, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0.0001110382, 0.005544296, 0.0002424636, 0, 0.0008035921, 0, 0, 0, 
    -3.882498e-05, 0.0003281081, -0.000151944, -1.090893e-05, -5.04232e-06, 
    0, 0, 0, 0, -0.0001717872, 0, 0, 0, 0, 5.853676e-05, 0.001761321, 
    0.006274315, 0.0003393338, 0,
  0, 0, 0, 0.0006502501, -3.484084e-06, 0.01281734, -2.501e-05, 0, 0, 0, 0, 
    -1.521344e-05, 0, 0, -8.567553e-07, 0.004876326, -4.140817e-05, 
    0.01446479, -4.688736e-05, 0, 0, 0, 0, 0, -4.212089e-05, 0.005171211, 
    0.007650789, 0, 0,
  0, -8.60859e-06, 0.002107821, 0.0001472783, 0.0009469809, 0, 0, 0, 0, 0, 
    -0.0001129201, 5.869255e-05, 0, 0, -1.044666e-05, 0.002025056, 
    0.0004826898, 0.003986185, 0, 0, 0, 0, 0, 0, 0.0009011744, 0.001002511, 
    0, 0, 0,
  0, -7.312975e-05, 4.114506e-05, 0.0002904622, 0.01451078, 0.001046071, 
    0.006233099, 0.02639629, -1.569695e-05, -5.136649e-05, 1.086238e-07, 
    0.00647644, -0.000212614, 0.01510649, 0.01158834, 0.002823159, 0, 
    -4.720325e-07, 0, 0, 0, 0, 0, 0.002402747, 0.01016769, 0.002017933, 
    -1.710646e-05, 0, 0,
  0, -2.249574e-06, 0, 0, 0, -4.634742e-05, 0.004124275, 0.00200846, 
    -3.916972e-05, 0.02679086, 0.004228192, -0.0002563643, 0.00335636, 
    0.01736109, -1.03397e-05, -1.402806e-06, 0, 2.560623e-05, 0, 0, 0, 0, 0, 
    0.01202799, 1.676016e-05, 0.0007584669, -1.613822e-05, 0, 0,
  0, 0, 0, 0, -2.040066e-05, 0.002356025, 0, 0, 0.02038958, 0.01101717, 
    0.00383366, -0.0001465167, 0.02193787, 0.01607474, 0.0001449715, 
    0.002506416, 0.0003821972, 0.004513296, -0.0003318606, 0.004845988, 
    0.008418002, 0, 0, -1.975292e-06, 0, -5.542534e-06, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.007837872, 0.0005623864, 0, 0, 0, 0, 
    -6.450142e-06, 1.666261e-05, 0.0002455285, 0, 0, 0, 0, 0, 0.003119305, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0.000123413, 3.887249e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -4.279056e-05, 7.661896e-05, 0.0001794299, 0, 0, 0, 0, 0, 0, 0, 
    -4.12127e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -3.29278e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0.009628755, 0, 0, 0, 0, 0, 0, 0, 0.006985866, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, -2.661966e-05, 0, 0,
  0, 0, 0.003639916, 0.01388979, 0.003619708, 0.001508264, 0.001167461, 0, 0, 
    0, 0.0004809425, 0.01051467, 0.001441111, -3.744558e-05, 9.425898e-06, 0, 
    -1.919799e-05, 0, -7.976916e-05, 0.0003408936, 0, -8.167708e-05, 0, 0, 
    0.00387664, 0.004592516, 0.01122996, 0.002591036, 0,
  0, 0, 0, 0.00460115, -2.556238e-05, 0.01958862, 0.0002347973, 0, 0, 0, 0, 
    -9.42828e-05, -2.035213e-05, 0, 0.003414814, 0.00695906, 0.0001207757, 
    0.02308322, 0.001733989, 0.0002259451, 0, 0, 0, 0, 0.002025648, 
    0.007127889, 0.01555414, 0, 0,
  0, -1.596265e-05, 0.006648466, 0.0002998435, 0.006447611, 0, 1.655753e-05, 
    0, 0, 0, 0.0004953732, 0.0004833475, -1.682356e-05, 0, 0.0006688162, 
    0.006195877, 0.003473891, 0.009392868, 0, 0, 0, 0, 0, 0, 0.003191264, 
    0.002235554, 0, 0, 0,
  0, 0.0009971875, -1.865242e-05, 0.001937513, 0.03956347, 0.007600089, 
    0.01931052, 0.03938312, 0.0001392651, -0.0001310691, -1.133526e-05, 
    0.01069039, 0.0004591348, 0.04045695, 0.03370573, 0.00666806, 0, 
    -7.222644e-06, 0, 0, 0, 0, 0, 0.008421401, 0.01204528, 0.01053001, 
    0.0001447861, 0, 0,
  0, 0.0004230711, 8.192358e-06, 0, -6.852459e-06, -0.0001468718, 0.02089968, 
    0.004646315, 0.0002710565, 0.04507184, 0.007732647, 0.0005641487, 
    0.01232028, 0.03019584, -4.646495e-05, -3.788686e-06, -1.213226e-05, 
    0.000487804, 0, -2.103731e-07, 0, 0, 0, 0.02482928, 0.0008201169, 
    0.005856593, 0.000518674, 1.411398e-06, 0,
  0, 0, 0, 0, -9.669466e-05, 0.006808992, 0, -1.036344e-05, 0.03074425, 
    0.01595357, 0.01001779, -0.0001782449, 0.03679422, 0.02790517, 
    0.009151157, 0.01018313, 0.0004025378, 0.006260408, 0.0005556642, 
    0.01769449, 0.02158273, 0, 0, 3.480426e-05, -3.009552e-06, 0.0003396722, 
    -4.018879e-05, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01137306, 0.001580314, 0, 0, 0, 0, 
    0.001528782, 0.002422024, 0.0007951916, 0.000100914, 0, 0, 0, 0, 
    0.01835957, -5.191507e-05, 0, 0, 0,
  0, 0, 0, 0, 0.0001876827, 0.0005916921, 0, 0, 0, -3.997925e-06, 
    -3.191173e-06, -3.847375e-08, 0, 8.069645e-05, 0.001056622, 0.002436631, 
    0.00511507, 0.004492735, -2.041685e-05, 0, 0, 0, 0, 0, -7.497372e-05, 
    -5.094329e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.648408e-05, -2.723202e-05, 
    0.001790178, 0, 0, 0, 0, 0, 0, 0.0007122643, 0.0001880674, 0, 
    0.0009140857, 0.0004379798, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2.305285e-05, 6.8351e-06,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.205374e-07, 0.0007542556, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  -7.575732e-06, 0, 0, 0, 0.01428465, -3.987203e-06, 0, 0.001544107, 0, 0, 0, 
    -3.129204e-06, 0.01628353, 0, 3.541767e-06, 0, 0, 0, -2.284356e-05, 
    -1.351171e-08, 0, 0, 0, 0, 0, -1.431072e-05, -7.825028e-05, 
    -4.131617e-11, 0,
  0, 0, 0.007809438, 0.02558712, 0.00788957, 0.004798847, 0.005488659, 0, 0, 
    -9.244069e-06, 0.002102923, 0.02730497, 0.007459623, -8.6091e-05, 
    0.005443149, 0.003307374, 0.001696883, 0.001975182, 0.002712412, 
    0.007148316, 0.0004740269, 0.00416011, -6.081681e-06, 0, 0.01125587, 
    0.0130052, 0.0316648, 0.009092677, 0,
  0, 0, -2.062259e-05, 0.01594466, 0.005670078, 0.03357372, 0.007014187, 
    -1.093102e-06, 0, 0, 3.669801e-06, 0.0003615338, -2.233883e-05, 0, 
    0.01301936, 0.01334914, 0.004430815, 0.04126295, 0.007508366, 
    0.001098979, -1.853492e-05, 0, 0, 0, 0.01091078, 0.01081586, 0.02603894, 
    -5.572787e-06, 0,
  0, -0.0006405989, 0.01827555, 0.0009190254, 0.01311716, 3.53219e-05, 
    0.00303936, 0, 0, 0, 0.02519304, 0.002579361, 2.176216e-05, 0, 
    0.005268031, 0.02254655, 0.01142841, 0.02235119, -2.093865e-08, 0, 0, 0, 
    0, -5.837428e-06, 0.01196676, 0.003881308, -1.767113e-05, 0, -4.092418e-10,
  0, 0.004948414, 0.0002408013, 0.005802019, 0.05441263, 0.01269452, 
    0.05285545, 0.05934758, 0.001264697, 3.288368e-05, 0.0004101931, 
    0.01973041, 0.0039456, 0.08631663, 0.07367399, 0.01258358, -2.053141e-05, 
    -1.998871e-05, -9.241662e-11, 0, 0, 0, 0, 0.03575388, 0.02439761, 
    0.03020705, 0.0001688053, -6.021182e-10, 0,
  0, 0.0004972643, 0.0004107628, -1.183568e-05, -9.682248e-05, 0.0003433301, 
    0.03958571, 0.01111719, 0.002083343, 0.06486233, 0.01479785, 0.008420497, 
    0.05106942, 0.05112601, 0.00063144, -8.605421e-06, 0.0006701699, 
    0.001210451, -1.00261e-05, -1.013642e-05, 0, 0, 0, 0.04205707, 
    0.001661764, 0.02153489, 0.003440015, -1.51222e-07, 0,
  0, 0, 0, 5.47581e-05, 0.0002568137, 0.01291595, 0, -1.646669e-05, 
    0.04221257, 0.02390542, 0.01897541, 0.003681513, 0.0506697, 0.04486791, 
    0.02274453, 0.0232159, 0.002847862, 0.008202182, 0.003432107, 0.03168598, 
    0.03249879, 0, -2.285035e-05, 4.650576e-05, -2.560097e-05, 0.0007231022, 
    -3.447695e-05, 1.236855e-09, 0,
  0, 0, 0, 0, -6.23919e-09, 0, 0, 0, 0, -3.992517e-05, 0.01156369, 0.0019154, 
    -1.388047e-08, -4.409909e-09, 0, -5.500125e-09, 0.007583093, 0.01263304, 
    0.002680253, 0.0003378765, -1.89158e-05, 0.0001627353, 0, 0, 0.02682209, 
    -9.875535e-05, 0, 0, -1.620731e-05,
  0, 0, 0, 0, 0.001412819, 0.001502086, -1.179761e-06, 0, 0, 7.786284e-05, 
    0.003186944, 8.04605e-06, 1.890026e-05, 0.003552868, 0.008366167, 
    0.008286111, 0.02073096, 0.01947948, 0.01185466, 0.004583507, 0, 
    0.006384028, 0.0001536881, -6.404978e-07, 0.00362613, 0.002404005, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0007322597, 8.853557e-05, 
    0.007343402, 6.604754e-05, 5.229581e-05, 0, 0, 0, 0, 0.003793882, 
    0.001677025, 0.0009459222, 0.004435332, 0.002163085, 0.0001175149, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -8.316912e-09, 0, 0, 0, 0, 
    0, 0, -1.12881e-05, 0, 0.001221, 0.001066646, 0.001813818, 0.0009857033,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, -1.523246e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0.003110949, 
    -3.252802e-05, 0.002605237, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.0007582987, 0, 0.002464622, -4.804431e-05, 0.02010142, -0.0002234738, 
    -9.840417e-06, 0.00308537, -0.000171636, 0, 0, 0.001309805, 0.026154, 
    -1.120706e-05, 0.003451345, -3.7709e-06, 0, 0, -3.994986e-05, 
    5.824382e-05, 0.0003136594, -4.600645e-07, 0, 0, 3.44151e-05, 
    0.000524929, 0.004116623, 0.0003483426, -7.484047e-05,
  1.929646e-09, -3.432292e-05, 0.01187406, 0.03842812, 0.02412365, 
    0.01353283, 0.01186443, -4.658355e-05, -2.548367e-10, -2.957582e-05, 
    0.006871669, 0.041643, 0.01480965, 0.003193685, 0.01758384, 0.01520714, 
    0.007610492, 0.002985553, 0.0119228, 0.01314903, 0.008262226, 
    0.006380526, 9.968843e-05, 0, 0.02610612, 0.03166243, 0.05280895, 
    0.01695633, -0.0001254897,
  -7.190788e-09, 1.129241e-06, 0.0004746096, 0.04240362, 0.0352462, 
    0.04682259, 0.02977247, -1.61169e-05, 0.0001563945, -1.362155e-07, 
    0.0008875381, 0.003761168, 0.001060572, -6.78167e-05, 0.02497975, 
    0.03543168, 0.02381298, 0.06512035, 0.02226138, 0.008505129, 0.001149231, 
    0, 0, -1.540016e-08, 0.0291352, 0.02674324, 0.04631621, -2.866672e-05, 
    -7.646542e-08,
  -6.049778e-10, 0.00994935, 0.06380494, 0.01325492, 0.02091779, 
    2.168182e-05, 0.02946751, -2.858147e-07, 7.503249e-05, 4.353365e-06, 
    0.1153815, 0.01960876, 0.00221244, 0.0001956571, 0.09739076, 0.1067402, 
    0.04554953, 0.0472417, 0.00290526, -3.874861e-08, -2.446955e-05, 0, 
    -5.028548e-07, 0.009749105, 0.06438962, 0.01399591, 0.0002394633, 
    1.544907e-05, 0.0002356438,
  5.117307e-07, 0.02873719, 0.03183071, 0.0186075, 0.07909329, 0.02640055, 
    0.1162742, 0.08883455, 0.01050634, 0.01989686, 0.005675047, 0.09248292, 
    0.03918666, 0.2529309, 0.2515938, 0.1254628, 0.0002952678, 0.0002143316, 
    -2.851432e-05, 2.943336e-07, 0, 0, 1.146747e-06, 0.1224087, 0.1131552, 
    0.06873024, 0.005474485, 0.0005703332, -5.16859e-09,
  5.894316e-07, 0.002814929, 0.00649111, 0.00209493, 0.001375732, 
    0.003003375, 0.06374553, 0.02129284, 0.02639225, 0.1497669, 0.03403081, 
    0.02752209, 0.1884303, 0.1127076, 0.007325909, 0.007827622, 0.001060363, 
    0.007091342, -5.547866e-05, 0.011056, 2.187651e-09, 0, 2.139169e-06, 
    0.1226613, 0.0255826, 0.03804263, 0.01461887, -3.708003e-06, 0,
  3.764549e-06, 0, -3.50265e-08, 0.0006967907, 0.004827109, 0.01980015, 
    -1.43811e-08, 1.510951e-05, 0.04772224, 0.04374209, 0.06066145, 
    0.0242078, 0.1194631, 0.08588642, 0.05541405, 0.04064098, 0.006549051, 
    0.01280701, 0.02000228, 0.0361335, 0.04920938, 0.0007896521, 
    0.0001435548, 0.0009672035, 0.0003454813, 0.00226971, -9.4084e-05, 
    0.0003826657, 2.813661e-05,
  6.079752e-05, 0, 0, -3.471063e-06, -1.113144e-06, -8.658926e-10, 0, 0, 0, 
    0.001858751, 0.009166151, 0.01489685, -4.065507e-05, -1.098066e-06, 
    2.647129e-06, -4.412238e-07, 0.02486421, 0.0356605, 0.01903659, 
    0.01520706, 0.002921358, 0.002801194, 0, 0, 0.03788793, -0.0002338185, 
    2.195651e-07, 0, -0.0001133985,
  0, 0, 0, 0, 0.002091499, 0.005694067, -2.469939e-05, 0, 0, 0.01260871, 
    0.02195867, 0.002718635, 0.004863041, 0.00846559, 0.0168332, 0.01374592, 
    0.04188681, 0.03684002, 0.02922084, 0.01137022, -0.0001473799, 
    0.01803638, 0.002055927, 5.477235e-05, 0.01492638, 0.005848286, 0, 0, 0,
  0, 0, 3.608292e-06, -2.164129e-05, 0, 0, -1.360534e-05, 0, 0, 0, 0, 0, 
    0.0005692907, 0.002613547, 0.005511947, 0.01779145, 0.003265044, 
    0.002906642, 0, 0, 0, 0.0007595887, 0.01038167, 0.01751489, 0.01801584, 
    0.01590394, 0.01086443, 0.002131817, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -5.604747e-05, -1.836464e-06, 
    0.00204928, -7.729252e-06, -1.798546e-05, 0, 0, 0, 0, 0.0004027947, 
    0.0009566325, 0.0103421, 0.004606302, 0.006036902, 0.004150087,
  0, 1.865086e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.0007279041, 0, 0.0001348025,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.938165e-08, 0.0001200178, 0, 
    -5.368003e-10, -9.114291e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0.0004147071, -1.538146e-05, -7.484346e-06, 0, 0, 0, 0, 
    8.390621e-06, -2.278156e-05, 0.0001273011, 0.005742981, 0.001917648, 
    0.003815545, 0.0002188741, 0, 0, 0, 0, 0, -1.349623e-06, 5.001201e-05, 0, 
    0.002110448, 0, 0,
  0.006291689, 0, 0.00584847, 0.001050278, 0.04335534, 0.01082255, 
    0.005198679, 0.01589695, 0.001547089, 0.0002909096, -7.072552e-05, 
    0.003439655, 0.03144082, 0.001171818, 0.003990982, 0.000171084, 
    4.234144e-07, 2.117817e-05, -3.902511e-05, 0.00337345, 0.001077007, 
    0.002116009, 0.003353736, 9.903572e-05, 0.001481465, 0.004558542, 
    0.01773395, 0.01097224, 0.005563447,
  0.0005809736, 0.0005207623, 0.02068886, 0.07175279, 0.06148064, 0.04748983, 
    0.03464724, 0.007558462, 0.008055507, 0.0003752679, 0.02480711, 
    0.05182793, 0.03460812, 0.007592686, 0.02530382, 0.02604057, 0.01951573, 
    0.01052516, 0.02750766, 0.02292811, 0.02239674, 0.01221131, 9.827807e-05, 
    -1.597461e-06, 0.03591435, 0.05845828, 0.1097022, 0.03672919, 0.01278058,
  0.0004389279, 1.855901e-06, 0.02170772, 0.1613965, 0.1288791, 0.1062925, 
    0.08012125, 0.0249414, 0.03943024, 0.03142948, 0.007657018, 0.07604747, 
    0.0299731, 0.003901455, 0.04227755, 0.08666725, 0.08314227, 0.1122213, 
    0.1337868, 0.0235669, 0.006025682, 0.000906742, -7.340228e-05, 
    0.01896663, 0.07977819, 0.149559, 0.1418602, 0.04343144, 0.01895895,
  8.031197e-06, 0.04471185, 0.2847563, 0.05621329, 0.04609237, 0.02111573, 
    0.08600323, 1.840525e-05, 0.004044677, 9.508889e-06, 0.2424988, 0.111799, 
    0.0149394, 0.01232442, 0.1439705, 0.1983567, 0.2085444, 0.3198966, 
    0.07906881, 0.005442901, 0.00577725, 0.0005415444, 0.0008925473, 
    0.03890019, 0.1025612, 0.1565223, 0.06260638, 0.01488376, 0.005447309,
  0.00105324, 0.1754744, 0.3516198, 0.182702, 0.1559675, 0.1052442, 
    0.2499054, 0.1800678, 0.06172986, 0.05117839, 0.03895605, 0.1278352, 
    0.09338386, 0.2564584, 0.260237, 0.1435348, 0.06020899, 0.03682276, 
    0.007339616, 5.564301e-05, 0.0002853979, 5.478947e-07, 0.0177041, 
    0.326265, 0.3296216, 0.3164224, 0.2080316, 0.03623459, 1.896371e-06,
  0.00291297, 0.1446822, 0.1294311, 0.08045955, 0.06055841, 0.07910303, 
    0.1108857, 0.07731118, 0.3245514, 0.5037224, 0.123552, 0.06294923, 
    0.2015208, 0.126865, 0.02151606, 0.01195154, 0.02594738, 0.01862848, 
    0.001618658, 0.02221337, -2.391347e-07, 8.830382e-07, 0.002405019, 
    0.3172444, 0.2955022, 0.1201961, 0.2337136, 0.002730928, 1.240195e-06,
  0.002204113, 4.774879e-05, 2.157438e-06, 0.001291459, 0.04613509, 
    0.06356255, 2.422576e-06, 0.005726273, 0.09082808, 0.1264807, 0.0891426, 
    0.05033667, 0.1030179, 0.08176759, 0.06409369, 0.09095109, 0.06757203, 
    0.1316887, 0.05044896, 0.1148317, 0.2043909, 0.04787591, 0.01476677, 
    0.01096483, 0.04531718, 0.03642302, 0.002397071, 0.09390406, 0.002318268,
  0.0001920035, 0.0003030804, 0, -3.201755e-05, -4.106282e-05, 1.848117e-06, 
    -9.729381e-10, 0, -2.362016e-06, 0.02614715, 0.01085476, 0.07257491, 
    0.002245562, -9.561068e-05, 3.197261e-06, 6.439565e-06, 0.09213921, 
    0.1268791, 0.1443672, 0.08757934, 0.1547342, 0.04321309, 0.0103149, 
    0.000435318, 0.07137708, 0.01300047, 0.0001049676, 0.0003604078, 
    0.001117671,
  0, -4.103734e-06, -1.538596e-08, -5.677304e-07, 0.002931311, 0.02942379, 
    0.0003776625, 0, 0, 0.02613533, 0.05223262, 0.01493121, 0.0228986, 
    0.01516337, 0.02440909, 0.05458853, 0.05834874, 0.06850902, 0.0572753, 
    0.02584508, 0.001593266, 0.04416445, 0.01016446, 0.02740874, 0.03550202, 
    0.01219962, -7.821584e-07, 0, 0,
  -1.636282e-05, 0, -3.599876e-06, 0.0007144846, -0.0001005379, 
    -2.060507e-05, 0.001567998, 0, 0, 0, 0, 0.001361796, 0.002535472, 
    0.006379875, 0.02804916, 0.05046602, 0.01247927, 0.01200159, 
    -1.687595e-05, -3.27885e-12, 0, 0.003538283, 0.02234321, 0.04975428, 
    0.0514059, 0.02997581, 0.03139509, 0.01364215, -2.254779e-05,
  0.000566678, 0.0004555106, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0009558971, 0.0007839969, 0.007379359, 0.001554705, 0.001142825, 
    -4.973653e-06, -8.633552e-07, 0, -0.0001166692, 0.0007298603, 
    0.004626563, 0.02313004, 0.02109047, 0.01726195, 0.01235552,
  -0.0001586169, 3.005029e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -2.042814e-05, 0, 0, 0, -2.814732e-06, 0, 0, 0.00085045, 0, 0, 0, 0, 
    0.0009656346, 0.005141766, 0.000762449, 0.002450169,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0005299954, 0.0002119811, 
    0.001572431, -3.524811e-05, 1.130508e-05, -5.84317e-06, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  0.00308677, 0, 0, 0, 0.003419797, 0.003460679, 0.01358468, 1.604603e-05, 0, 
    0, -1.403226e-05, 0.005800589, -7.449843e-05, 0.01660694, 0.03617125, 
    0.02304738, 0.01071549, 0.00823546, -1.637699e-05, 0, 0, 0, 0, 
    0.0001358604, 0.002563515, 0.0001196532, 0.002880648, -9.758293e-06, 0,
  0.01314845, 0.002277695, 0.009592571, 0.009092279, 0.09800118, 0.08838134, 
    0.03386724, 0.05631921, 0.03760873, 0.003334183, 0.002394057, 0.0136274, 
    0.05065762, 0.04524241, 0.03190361, 0.03571036, 0.009362983, 0.004218276, 
    0.006702898, 0.006149147, 0.002922247, 0.006123481, 0.01780629, 
    0.000922351, 0.008146103, 0.0221163, 0.02974685, 0.04640077, 0.02936987,
  0.04678754, 0.0409194, 0.04892414, 0.1061218, 0.1052622, 0.104891, 
    0.1176314, 0.06365359, 0.04457455, 0.04869078, 0.1012064, 0.1255923, 
    0.08439878, 0.07832313, 0.03894647, 0.1336698, 0.1134007, 0.04647318, 
    0.1213258, 0.1350351, 0.1036643, 0.05387314, 0.007449654, 0.002607626, 
    0.06790289, 0.1486616, 0.2144936, 0.1199386, 0.06673758,
  0.001053426, 0.0005117753, 0.0462652, 0.1510275, 0.1288722, 0.1234722, 
    0.1011831, 0.02166934, 0.05141265, 0.03418883, 0.02928394, 0.1167913, 
    0.11596, 0.06946927, 0.1422356, 0.1787392, 0.1772926, 0.1433807, 
    0.258497, 0.2113859, 0.0414669, 0.04760095, 0.02534223, 0.00756836, 
    0.09190352, 0.1906705, 0.2034722, 0.06176082, 0.02135139,
  8.840241e-07, 0.02378466, 0.2594064, 0.04013189, 0.03544354, 0.01229794, 
    0.08049298, 0.002450205, 0.004786805, 3.60911e-05, 0.2120719, 0.08098724, 
    0.01369078, 0.004856614, 0.1461541, 0.1771258, 0.1602746, 0.2853609, 
    0.06239972, 0.02430736, 0.02819558, 0.0001260669, 0.004117537, 
    0.02937484, 0.07818422, 0.2372313, 0.07231552, 0.01338782, 0.0003188073,
  0.001524387, 0.142439, 0.3065177, 0.1448487, 0.1258779, 0.07924754, 
    0.1877212, 0.1442658, 0.03958496, 0.04635903, 0.02654106, 0.104446, 
    0.07132948, 0.2075152, 0.1986568, 0.08035055, 0.02252848, 0.009266222, 
    0.000442688, 1.32273e-05, 3.047376e-05, 9.475734e-08, 0.000464835, 
    0.2823631, 0.2693366, 0.2940972, 0.1843291, 0.0017906, 3.24511e-06,
  0.000152535, 0.1078441, 0.07376175, 0.03778245, 0.04353726, 0.06983802, 
    0.09661645, 0.0603192, 0.2636593, 0.4662485, 0.09466902, 0.04739236, 
    0.1441509, 0.115899, 0.01754544, 0.0109649, 0.0202673, 0.01753603, 
    0.000587234, 0.007234775, -7.124118e-08, 5.83404e-08, 0.00300701, 
    0.2445615, 0.1788375, 0.1107979, 0.1835136, 0.0002034659, 2.188168e-07,
  3.885845e-05, 5.101041e-05, -5.812512e-06, 0.01331008, 0.04207463, 
    0.03340995, 1.03421e-05, 0.001682309, 0.07104853, 0.09481534, 0.06599983, 
    0.03793756, 0.07650524, 0.07621852, 0.06669401, 0.07132311, 0.05650407, 
    0.1178605, 0.0417318, 0.07830565, 0.1489102, 0.02757756, 0.005038345, 
    0.003062516, 0.02926616, 0.02879449, 0.01174001, 0.1537781, 0.09000544,
  0.1378283, 0.02608551, -1.878234e-07, 5.001053e-07, 4.64933e-05, 
    0.002371192, -4.253851e-05, -7.886767e-12, 4.267543e-06, 0.02936535, 
    0.00695966, 0.05573924, 0.003514769, 0.002275685, 9.922655e-06, 
    0.0002903861, 0.1073958, 0.1375289, 0.1748655, 0.1029744, 0.1373744, 
    0.03723192, 0.007153849, 0.0008262252, 0.06519108, 0.06617839, 
    0.002076732, 0.0005909939, 0.1751438,
  -6.805375e-06, -0.0003378965, 0.001039135, -1.543415e-06, 0.003867667, 
    0.06664021, 0.01931754, 0, 0, 0.03113386, 0.06527648, 0.03868868, 
    0.03513641, 0.02750568, 0.0468534, 0.1593519, 0.1185997, 0.130781, 
    0.1301881, 0.1016307, 0.01447121, 0.1411903, 0.122719, 0.05489809, 
    0.1678412, 0.1719205, 0.04016247, 0.001037647, -1.329973e-05,
  0.001568137, 0.001237587, 0.001707394, 0.001721548, -0.0002071169, 
    0.0009089844, 0.001957571, 0, 0, 0, 0.0002146473, 0.003176916, 
    0.006042523, 0.01967395, 0.07323678, 0.08688215, 0.03407932, 0.06990654, 
    0.004967555, -0.0002817353, -1.699011e-05, 0.009515208, 0.0568255, 
    0.09989668, 0.1033735, 0.07512104, 0.09274341, 0.04409844, 0.002320336,
  0.001664322, 0.002728507, -1.554991e-05, -4.750901e-06, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, -3.917886e-05, 0.01859766, 0.007056606, 0.01232614, 0.005133721, 
    0.0177528, 0.003795653, 0.0002681158, -6.894917e-12, -0.0002842942, 
    0.004274349, 0.009157758, 0.03895585, 0.03821649, 0.04044969, 0.02374939,
  0.00322584, 0.001276386, -7.151029e-05, -3.597178e-08, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, -6.889366e-05, 0.002020898, 0.003393431, 0.0003032202, 
    -7.163486e-05, -2.602146e-05, -2.44016e-05, 0.003810409, -2.129386e-05, 
    0, 0, 0, 0.004068542, 0.01071947, 0.01190654, 0.01232096,
  0, 1.966135e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0.0003170591, 0.003417239, -2.591798e-06, 0, 0, 0, 0, 
    0.002061072, 0.001885731, 0.005731134, 0.005782903, 0.007680518, 
    0.006013444, 0.00116191, -1.545685e-05, 0, 0, 0, 0, 0.001686604, 0, 
    6.249773e-06, 0, 0,
  0.006785171, -7.962875e-05, -1.045399e-07, 0.001258916, 0.0118933, 
    0.01982295, 0.03734099, 0.01087823, 0.00862439, -2.772815e-05, 
    0.0001956518, 0.006543011, 0.01111476, 0.02648157, 0.06300981, 
    0.06656771, 0.0323625, 0.03210473, 0.02138707, 0.01016934, 0.002374386, 
    -4.11447e-05, 0.0003657858, 0.003167443, 0.0117449, 0.007545199, 
    0.007474275, 0.008512278, -0.0001344515,
  0.09684977, 0.07503981, 0.1008043, 0.1219303, 0.1715701, 0.1894938, 
    0.1434286, 0.1906345, 0.1476687, 0.05360879, 0.03698862, 0.07557503, 
    0.0916937, 0.1424198, 0.1231059, 0.138113, 0.1002515, 0.08258435, 
    0.08877163, 0.05803834, 0.06148574, 0.08420145, 0.1118142, 0.01785504, 
    0.03970822, 0.07313279, 0.07726904, 0.08796086, 0.09447248,
  0.0519908, 0.06695294, 0.05598597, 0.08802036, 0.1112259, 0.08840601, 
    0.1065979, 0.08196543, 0.07525845, 0.07379785, 0.130141, 0.1352227, 
    0.09548943, 0.09317529, 0.09004326, 0.1501855, 0.1761115, 0.09812734, 
    0.123782, 0.1698242, 0.1369069, 0.1602639, 0.05834875, 0.03042253, 
    0.1054401, 0.1512381, 0.2476097, 0.1688464, 0.08365735,
  0.001792739, 0.0004316303, 0.0593135, 0.1263922, 0.1392632, 0.1123926, 
    0.1132982, 0.02360478, 0.0393582, 0.04071448, 0.02947429, 0.1120668, 
    0.1161865, 0.0530653, 0.1126677, 0.1672489, 0.1457528, 0.1373487, 
    0.2120963, 0.2153296, 0.0337685, 0.03605313, 0.00203354, 0.0003478272, 
    0.06279122, 0.158163, 0.1642001, 0.04194244, 0.01386589,
  4.484019e-06, 0.01196622, 0.2394493, 0.04138711, 0.03349926, 0.01168465, 
    0.06858809, 0.0005041777, 0.003864739, 2.074e-05, 0.1818342, 0.06721242, 
    0.0100322, 0.001614559, 0.1474732, 0.1684712, 0.1299006, 0.2544676, 
    0.05723614, 0.02407378, 0.0176589, 1.248665e-05, 0.007850736, 0.01823401, 
    0.07075478, 0.1988146, 0.03361401, 0.004484606, 0.001411032,
  4.446973e-05, 0.108221, 0.2556277, 0.1274492, 0.1202808, 0.06336462, 
    0.1684867, 0.1407524, 0.04087418, 0.04304289, 0.02233224, 0.08160413, 
    0.07127258, 0.1745828, 0.1750091, 0.05991291, 0.009013551, 0.009583741, 
    0.0002191535, 3.926941e-06, 2.063568e-06, -8.420693e-09, 1.849862e-05, 
    0.2633913, 0.260304, 0.2720902, 0.1358393, -0.0001317239, 2.223474e-06,
  0.0001306294, 0.0766855, 0.03697428, 0.01861275, 0.03390152, 0.07019896, 
    0.09638516, 0.05783798, 0.2001336, 0.4208677, 0.07830641, 0.03212195, 
    0.1259499, 0.1228802, 0.0171156, 0.01012823, 0.01245998, 0.007274666, 
    0.0002205326, 0.0004118466, -4.431696e-08, 3.409557e-07, 0.004115901, 
    0.1657004, 0.1328943, 0.09916297, 0.1441307, -5.962721e-05, 2.535974e-07,
  3.746126e-06, 1.217928e-05, 4.670346e-05, 0.01324421, 0.05021924, 
    0.0233104, 2.602711e-06, 0.002106885, 0.07380777, 0.07932257, 0.05893837, 
    0.03510865, 0.06980626, 0.07144137, 0.07797415, 0.0631575, 0.05698662, 
    0.1088567, 0.0292301, 0.07905117, 0.1148997, 0.01860063, 0.003397917, 
    0.003074756, 0.01757296, 0.03011568, 0.0323212, 0.1490133, 0.05419998,
  0.1199946, 0.01169316, -5.828094e-08, 9.542716e-06, -3.369727e-06, 
    0.001107467, 0.0002691747, -4.071178e-11, 0.0005511391, 0.0341208, 
    0.01334198, 0.04057819, 0.001623187, 0.01221703, 4.78465e-05, 
    0.002727771, 0.1059825, 0.1347035, 0.1921098, 0.07624594, 0.1190285, 
    0.03077292, 0.005653062, 0.001707011, 0.07083587, 0.05904613, 
    7.401437e-05, 0.001373942, 0.2160635,
  0.01865505, 0.02872933, 0.02676405, 0.0006063718, 0.01914687, 0.1396486, 
    0.08228676, 0, 0, 0.03391675, 0.07512867, 0.04469935, 0.0343617, 
    0.04790761, 0.1036392, 0.203586, 0.1289832, 0.1810247, 0.1890912, 
    0.1143032, 0.06602781, 0.1861208, 0.1286116, 0.035481, 0.1432577, 
    0.1657991, 0.1134884, 0.01371286, 0.006381546,
  0.01894774, 0.00412599, 0.009870453, 0.007386645, 0.002213041, 0.002910644, 
    0.003523752, 0, 0, -6.805472e-10, 0.001408849, 0.004267962, 0.01289369, 
    0.05005986, 0.1390806, 0.1700941, 0.1041936, 0.1245588, 0.03989022, 
    0.01016284, 0.0008039258, 0.04241951, 0.1216081, 0.1857496, 0.1928347, 
    0.1808568, 0.1397852, 0.1228298, 0.0418666,
  0.03076134, 0.01177997, 0.0005021852, 0.004052324, -3.500977e-08, 0, 0, 0, 
    0, 0, 0, 0, -6.955783e-05, 0.003340977, 0.05859516, 0.04575116, 
    0.02218674, 0.02950316, 0.05659653, 0.01697044, 0.0001745644, 
    0.0003084724, 0.007045367, 0.007314149, 0.04177862, 0.07208411, 
    0.1038594, 0.1105238, 0.1019317,
  0.02814805, 0.01683853, 0.002642786, 0.0001851242, -7.040427e-06, 0, 0, 0, 
    0, 0, 0, 0, 0, 6.635107e-05, 0.008056157, 0.009867051, 0.004515106, 
    0.004502154, 0.000722624, 0.0003769617, 0.00526908, 0.0001618836, 0, 0, 
    -1.177989e-05, 0.009519137, 0.01477314, 0.03231736, 0.03865337,
  0.0007868338, 0.004179391, 1.390679e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0008798481, 0.002590872, -1.729852e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -4.439229e-06, 0.002011047,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.693567e-08, 0, 0, 0, 0, 
    0, 0, -0.0001089338, 0.007001211, -0.00230458, 0.002141327, 0, 0,
  0, 0, 0, 0, -2.110064e-10, 0.002898676, 0.02176606, -0.000191249, 0, 0, 0, 
    0, 0.008967004, 0.007426624, 0.0224215, 0.0269009, 0.03165263, 
    0.02606579, 0.02052541, 0.01082268, 0.007997793, 0.0002784311, 
    3.812945e-05, 0.0001741478, 0.01020466, 0.01823541, 0.007683631, 
    0.0006182212, 0.0004997943,
  0.04356242, 0.04179191, 0.02571791, 0.03715428, 0.05603043, 0.08089977, 
    0.06984179, 0.05556647, 0.04954056, 0.01391987, 0.005413795, 0.0194183, 
    0.05278571, 0.08094398, 0.1386985, 0.1521884, 0.1617828, 0.09721151, 
    0.07999907, 0.04874494, 0.03545614, 0.03184875, 0.02165274, 0.05846595, 
    0.09248732, 0.08134972, 0.07188039, 0.06485213, 0.03818214,
  0.1386133, 0.1367667, 0.1391414, 0.1826957, 0.1711441, 0.183623, 0.1457182, 
    0.2156536, 0.1925971, 0.1408739, 0.1012937, 0.124797, 0.1818062, 
    0.1885696, 0.1553236, 0.1587769, 0.117203, 0.1365176, 0.1645006, 
    0.1292498, 0.1206098, 0.1551749, 0.1919699, 0.06822486, 0.09652419, 
    0.1261489, 0.1082832, 0.1524601, 0.1421296,
  0.05120045, 0.06065071, 0.03936303, 0.07368075, 0.1019164, 0.07278816, 
    0.09179294, 0.07166905, 0.06492072, 0.06293497, 0.1331359, 0.1120731, 
    0.07986817, 0.07767466, 0.08409339, 0.1459522, 0.1751136, 0.1050223, 
    0.1145213, 0.1840814, 0.1619882, 0.1468721, 0.06727121, 0.07032315, 
    0.1009807, 0.1319924, 0.2433755, 0.1775457, 0.1015572,
  0.002473962, 2.729523e-06, 0.06765769, 0.1226596, 0.1355014, 0.09760077, 
    0.1043801, 0.03528859, 0.05164565, 0.01689676, 0.02796419, 0.104767, 
    0.1121525, 0.02399776, 0.09710324, 0.1338999, 0.1164603, 0.136956, 
    0.2219741, 0.2012927, 0.02865416, 0.03015815, -7.980524e-05, 
    2.210616e-05, 0.04614232, 0.1453476, 0.1238478, 0.02500094, 0.006716402,
  0.0001325647, 0.009291692, 0.2135576, 0.03505887, 0.03085754, 0.009466458, 
    0.05085036, 0.006400171, 0.0005320348, 1.488224e-05, 0.1209949, 
    0.05003207, 0.01015818, 0.002531174, 0.126556, 0.1456505, 0.09551462, 
    0.2326991, 0.02566994, 0.02279391, 0.006493357, 1.148522e-06, 0.01840743, 
    0.01113778, 0.05342996, 0.1923956, 0.01489701, 0.002639431, 0.01311247,
  4.960838e-05, 0.07982098, 0.2258841, 0.1046746, 0.1031704, 0.05977915, 
    0.1356863, 0.1337626, 0.0335957, 0.0400796, 0.01731402, 0.06145964, 
    0.06870344, 0.1581872, 0.143031, 0.05672607, 0.007930881, 0.008947863, 
    0.0002209789, 1.058901e-06, 2.594209e-06, -4.209173e-09, 1.443478e-05, 
    0.2180122, 0.2412749, 0.2418444, 0.08713242, -0.0003678536, 1.819059e-06,
  0.0005838571, 0.05723098, 0.02006928, 0.01404019, 0.02475929, 0.06404129, 
    0.1010076, 0.04402106, 0.118358, 0.3564202, 0.06149279, 0.02066527, 
    0.09653495, 0.1264312, 0.02060995, 0.005454839, 0.005881024, 
    1.783401e-05, 9.170617e-05, 1.313821e-05, -3.632989e-08, 1.030634e-07, 
    0.01703946, 0.1236185, 0.1126036, 0.09801056, 0.09762575, -1.277115e-06, 
    2.242536e-07,
  8.649071e-05, 9.172742e-06, 3.233924e-05, 0.004962304, 0.04166144, 
    0.0159161, 3.480568e-05, 0.002174858, 0.08077681, 0.06497578, 0.05402569, 
    0.02556963, 0.07467686, 0.06733676, 0.06662963, 0.04845827, 0.05944059, 
    0.09220298, 0.01839385, 0.0638078, 0.08368079, 0.01021732, 0.002762238, 
    0.002102562, 0.01159837, 0.04154472, 0.05243128, 0.1162581, 0.01294823,
  0.1077396, 0.005296261, -3.200662e-07, 1.10866e-05, 0.0001047912, 
    0.008516303, 0.001390607, -2.113482e-07, 0.01523925, 0.0460499, 
    0.02906592, 0.03438657, 0.0009224112, 0.01407077, 0.002310733, 
    0.005168029, 0.08851166, 0.1322496, 0.1524428, 0.02795227, 0.1123155, 
    0.0310867, 0.002975854, 0.002746273, 0.0693248, 0.03623846, 2.852756e-05, 
    0.005613575, 0.2376917,
  0.02958087, 0.04134696, 0.03772301, 0.02475194, 0.04560415, 0.170558, 
    0.09217959, -1.466469e-10, -2.782531e-11, 0.04338047, 0.0759067, 
    0.05527855, 0.04582144, 0.05175379, 0.1039455, 0.1509259, 0.110494, 
    0.1586031, 0.1788209, 0.08651915, 0.06700551, 0.1750575, 0.09773739, 
    0.02413906, 0.105572, 0.1533172, 0.09177088, 0.009874524, 0.02753937,
  0.07539953, 0.02511831, 0.03566223, 0.02202025, 0.02174777, 0.03483233, 
    0.005463635, -1.783622e-05, 0, 0.0007316847, 0.007783577, 0.02089014, 
    0.02627167, 0.09114614, 0.1703762, 0.2216875, 0.1759371, 0.1575412, 
    0.04828845, 0.03631518, 0.009218029, 0.06928448, 0.2113244, 0.1978684, 
    0.1775831, 0.1871808, 0.1785654, 0.1190156, 0.1044457,
  0.093292, 0.04815502, 0.02913769, 0.01455034, 0.00985979, -4.245041e-05, 
    -4.016035e-06, 0, 0, 0, 0, 0, 0.006566567, 0.03047634, 0.1744423, 
    0.1875997, 0.1174515, 0.04861726, 0.06705853, 0.03408046, 0.001540459, 
    0.008361077, 0.01295066, 0.02086086, 0.07712778, 0.1322231, 0.1590794, 
    0.1908219, 0.2011361,
  0.1101556, 0.05528391, 0.04504797, 0.003243613, 0.0004511299, 0.000766783, 
    0, 0, 0, 0, 0, 0, 0, 0.007142762, 0.0677615, 0.1280863, 0.02391406, 
    0.03401009, 0.005992375, 0.007503355, 0.01038912, 0.001446965, 0, 0, 
    -0.0002352927, 0.01464086, 0.03015329, 0.06111814, 0.1113845,
  0.009234942, 0.01533509, 0.0006642483, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -4.148134e-05, 0.007658831, 0.01005044, 0.01601397, -4.093232e-05, 
    -9.265856e-07, 0.0004976755, 0, 0, 0, 0, 0, 0, -2.668416e-09, 
    0.0003745155, 0.007637498,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.140857e-05, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002972207, 0.01351414, 0.01640985, 
    0.0127055, 0.003508277, 5.176782e-06, 0, 0, 0, 0.00162038, 0.03344413, 
    0.05819099, 0.05872425, 0.07459807, 0.002143971, 0,
  -0.002433851, 0.01108717, 0.0005782974, 0.00779421, -0.0002473267, 
    0.005091358, 0.05397974, 0.00313867, -0.0006774808, 0, 0, -7.877647e-05, 
    0.01063448, 0.05206628, 0.06838465, 0.07969056, 0.06131969, 0.04341543, 
    0.04257599, 0.04839324, 0.03921144, 0.06297554, 0.05549026, 0.038047, 
    0.04188358, 0.04941968, 0.1265048, 0.05000911, 0.02061091,
  0.08048561, 0.1059367, 0.08355469, 0.1140386, 0.1741199, 0.1384108, 
    0.1287802, 0.09562565, 0.09523404, 0.06606437, 0.06231964, 0.07730161, 
    0.1253145, 0.1364708, 0.1944094, 0.2007562, 0.2028621, 0.1330181, 
    0.1482169, 0.1316616, 0.1187174, 0.08691173, 0.108339, 0.1319495, 
    0.1767521, 0.1208487, 0.1245351, 0.08850559, 0.1097334,
  0.1455412, 0.1653405, 0.1657382, 0.2203234, 0.1558699, 0.1793961, 
    0.1399132, 0.1892529, 0.1877079, 0.1428051, 0.1428267, 0.1180092, 
    0.1730719, 0.1984726, 0.1626747, 0.1423248, 0.1119018, 0.1275254, 
    0.1459337, 0.1232657, 0.1624783, 0.1819231, 0.2274892, 0.1182803, 
    0.108541, 0.142439, 0.1214497, 0.1642035, 0.1473467,
  0.04293348, 0.05308487, 0.03761867, 0.0685019, 0.09755877, 0.0641757, 
    0.08815506, 0.06686146, 0.04773503, 0.06391895, 0.1228512, 0.1017587, 
    0.07050642, 0.06851934, 0.07257709, 0.1397937, 0.1613261, 0.08538196, 
    0.09667731, 0.1733898, 0.1528755, 0.1471989, 0.05705698, 0.06488083, 
    0.09008405, 0.1249411, 0.2294662, 0.1763196, 0.1024678,
  0.001216328, 5.250236e-06, 0.07788973, 0.1134737, 0.1535286, 0.08002942, 
    0.08598143, 0.03709836, 0.04892804, 0.009157214, 0.02909178, 0.1130254, 
    0.1068141, 0.01478133, 0.08470635, 0.09156831, 0.1003112, 0.1465015, 
    0.2163609, 0.2045739, 0.05213706, 0.03068217, -0.0005488341, 
    1.942429e-05, 0.03488524, 0.1615118, 0.108497, 0.01578693, 0.002276428,
  2.966515e-07, 0.009588582, 0.1822007, 0.02684335, 0.02897269, 0.007932095, 
    0.03921113, 0.01683442, 2.261919e-06, 1.653544e-05, 0.07806587, 
    0.03010518, 0.008355766, 0.004004543, 0.09519963, 0.1477604, 0.06941102, 
    0.2008088, 0.01619025, 0.01866058, 0.001039625, 9.408904e-08, 
    0.007697423, 0.002911792, 0.03790653, 0.1958807, 0.008873651, 
    0.001455348, 0.00540132,
  5.084571e-05, 0.05596325, 0.1723492, 0.07578472, 0.08704653, 0.04802505, 
    0.1037663, 0.1261325, 0.02138113, 0.02708265, 0.01111149, 0.0410446, 
    0.05673085, 0.1373718, 0.1063495, 0.05112204, 0.01250434, 0.0122077, 
    0.0001641582, 3.475059e-07, 4.931372e-07, -2.269688e-09, 2.262726e-05, 
    0.1818396, 0.2169622, 0.2061217, 0.05010739, -0.0002296586, 5.278787e-06,
  -6.983316e-06, 0.04541216, 0.01464716, 0.009913341, 0.01795385, 0.04743947, 
    0.09549289, 0.04092964, 0.06483532, 0.2943267, 0.04427346, 0.01240142, 
    0.07698774, 0.1150118, 0.01500826, 0.002993337, 0.001521702, 
    -8.837721e-05, 4.566735e-05, -1.159522e-05, -3.702375e-10, 6.270449e-08, 
    0.01901391, 0.09268452, 0.07865904, 0.09765272, 0.07651526, 9.088657e-05, 
    1.617381e-07,
  0.006868973, 5.385736e-06, 8.368545e-06, 0.004218205, 0.03227359, 
    0.01154816, 3.117161e-05, 0.003245498, 0.07571784, 0.04673618, 
    0.03689795, 0.02104122, 0.06840209, 0.06430322, 0.06542422, 0.0304187, 
    0.05479794, 0.07551225, 0.02163141, 0.07229767, 0.0572491, 0.007012837, 
    0.002429967, 0.00189492, 0.01207862, 0.03403905, 0.05684549, 0.1085934, 
    0.006945876,
  0.09296134, 0.004732963, -1.218344e-09, 1.281899e-05, 0.0001915252, 
    0.001224708, 0.001741765, -6.983365e-09, 0.03045299, 0.06295753, 
    0.03224612, 0.0253463, 0.0005319624, 0.005672577, 0.009075924, 
    0.008232649, 0.077119, 0.1380839, 0.1172666, 0.01458597, 0.1104325, 
    0.02978043, 0.001540525, 0.001838268, 0.07121988, 0.03097708, 
    2.442886e-06, 0.006050591, 0.20947,
  0.04226559, 0.04362222, 0.03568328, 0.02109286, 0.05479866, 0.1642828, 
    0.08433293, -3.953181e-08, -9.224469e-06, 0.04768786, 0.0808343, 
    0.0805794, 0.05349334, 0.06649052, 0.1064766, 0.1226516, 0.1008537, 
    0.1443172, 0.158106, 0.07566074, 0.07732809, 0.1669183, 0.06856735, 
    0.01062949, 0.0591874, 0.1405439, 0.07280792, 0.01745041, 0.03316011,
  0.1371808, 0.0478895, 0.08212847, 0.05014297, 0.0755187, 0.08735747, 
    0.008292365, 0.034898, -5.917919e-06, 0.004733895, 0.04599993, 0.0560119, 
    0.04894654, 0.1197504, 0.2032049, 0.2097217, 0.1862291, 0.1435077, 
    0.04299432, 0.06100875, 0.0672543, 0.1017238, 0.2173846, 0.1982087, 
    0.1919096, 0.1675452, 0.1720896, 0.1001982, 0.08881144,
  0.1372047, 0.08920497, 0.1229922, 0.08326136, 0.1383938, 0.09989521, 
    0.003917072, -5.515868e-06, 0, 0, 0, -6.305543e-07, 0.02191013, 
    0.05357974, 0.2215843, 0.2207531, 0.1136548, 0.06941619, 0.09119556, 
    0.05401845, 0.02528564, 0.03425171, 0.04919634, 0.05317108, 0.1046092, 
    0.14919, 0.1670997, 0.1776453, 0.2038304,
  0.1802086, 0.1306079, 0.1164558, 0.08243193, 0.05027988, 0.01045462, 
    0.001380763, 0.0004511868, 0, 0, 0, 0, -0.0007620504, 0.01579024, 
    0.2124023, 0.1917179, 0.103628, 0.1046932, 0.02548653, 0.02885406, 
    0.02542825, 0.003247767, 0.002046538, 0, 0.00350489, 0.03188189, 
    0.05929505, 0.104008, 0.1636538,
  0.042239, 0.04965597, 0.01299502, 0.003167081, 9.12054e-06, 0, 0, 0, 0, 0, 
    0, 0, 0, 9.42115e-05, 0.05220053, 0.09678984, 0.09677391, 0.05573395, 
    0.0551049, 0.01534292, 9.242314e-05, 0, 0, 0, 0, 0, -6.68753e-05, 
    0.02477967, 0.02647405,
  0, 0, -1.203404e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.569491e-05, 
    0.002931193, 0.006975109, 0.004740444, 0.000747023, -3.339847e-06, 
    -3.784309e-07, 0, 0, -3.251527e-05, -3.707846e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.03849905, 0.05527312, 0.08105693, 
    0.08310569, 0.04428117, 0.005675044, 3.005679e-05, 0, 0, 0.01321843, 
    0.1368535, 0.1409185, 0.1288341, 0.1393439, 0.0133461, 0,
  0.008205065, 0.09880811, 0.09685943, 0.08907651, -0.002186968, 0.02685457, 
    0.07786793, 0.02586332, -0.0008156543, -0.0003026793, -8.252827e-06, 
    -0.0004798755, 0.02682474, 0.08942463, 0.1061888, 0.1175627, 0.1212655, 
    0.07685619, 0.06762227, 0.07107591, 0.07263732, 0.1616705, 0.1674285, 
    0.09934463, 0.09202911, 0.1788779, 0.2828655, 0.116607, 0.03993824,
  0.121245, 0.1701834, 0.1440126, 0.1657677, 0.1998919, 0.1772658, 0.1669449, 
    0.1438375, 0.1569209, 0.1342581, 0.1108186, 0.1936973, 0.1774088, 
    0.1715677, 0.2073622, 0.2135156, 0.2141991, 0.1692637, 0.1771841, 
    0.1636364, 0.151431, 0.1442873, 0.1753506, 0.1604252, 0.1833382, 
    0.1730986, 0.1692859, 0.1216679, 0.1650833,
  0.1657327, 0.1839697, 0.1696656, 0.2388266, 0.1688213, 0.1618193, 
    0.1534798, 0.1707345, 0.1666199, 0.1308492, 0.1505788, 0.1191235, 
    0.1739716, 0.1967954, 0.1673638, 0.1235204, 0.1141245, 0.1184914, 
    0.1223402, 0.116588, 0.1449008, 0.1775568, 0.2107576, 0.1370467, 
    0.1036772, 0.1392488, 0.1216936, 0.136866, 0.1682584,
  0.04176592, 0.04772545, 0.04123687, 0.06162384, 0.08611257, 0.05706638, 
    0.08124818, 0.04991363, 0.04193379, 0.04245596, 0.1240127, 0.09632508, 
    0.06975646, 0.05934475, 0.07692061, 0.1560552, 0.1557367, 0.06719609, 
    0.08153871, 0.1294768, 0.1377468, 0.1330598, 0.05843891, 0.0422182, 
    0.07896081, 0.1327464, 0.2109919, 0.1615936, 0.09837993,
  0.0004517875, -8.443536e-06, 0.08959664, 0.1130188, 0.160432, 0.06745739, 
    0.06474714, 0.03625084, 0.04080456, 0.009419246, 0.03213879, 0.1102469, 
    0.08796407, 0.009650359, 0.06975777, 0.06029746, 0.08487982, 0.1604849, 
    0.223516, 0.2187959, 0.04689906, 0.01910338, 7.847149e-05, 0.002543656, 
    0.02401851, 0.1475519, 0.0681868, 0.009761217, 0.001745346,
  1.425297e-07, 0.0103028, 0.1419799, 0.02048929, 0.02590596, 0.005964492, 
    0.02889675, 0.00359776, 2.217762e-06, 3.58231e-06, 0.04472331, 
    0.02038676, 0.004854382, 0.006857339, 0.07309283, 0.1325836, 0.05275181, 
    0.1764681, 0.01117371, 0.008039639, 5.604327e-05, 1.03419e-08, 
    0.00262444, 0.0009268452, 0.03813497, 0.1847901, 0.007404367, 
    0.0002545852, 0.0003524204,
  6.157035e-05, 0.04285803, 0.1245352, 0.05668346, 0.07675896, 0.0325761, 
    0.0926552, 0.1248715, 0.01253873, 0.02219696, 0.01003147, 0.03828908, 
    0.04229157, 0.123835, 0.08083524, 0.03166485, 0.01143224, 0.00855635, 
    0.0001813149, 2.242271e-07, 2.021948e-07, -5.536633e-10, 1.675496e-05, 
    0.136015, 0.2025695, 0.1844709, 0.02135877, -4.125451e-06, 7.804428e-06,
  0.02156685, 0.03264703, 0.01469128, 0.007650401, 0.01084616, 0.03326533, 
    0.08836791, 0.0383713, 0.03993275, 0.24209, 0.03599087, 0.007743364, 
    0.05952489, 0.1080424, 0.01058587, 0.00180036, 0.0001595354, 0.000793922, 
    1.229463e-05, 0.001967261, 2.265547e-08, -2.368608e-09, 0.0229324, 
    0.0774448, 0.03980714, 0.09812719, 0.06816441, 0.0001220786, -2.329076e-06,
  0.01674961, 2.194227e-06, 6.808105e-06, 0.006452382, 0.03199493, 
    0.009629809, 7.457269e-05, 0.002516523, 0.07524268, 0.03652341, 
    0.02832762, 0.02141449, 0.06308119, 0.07019836, 0.06883517, 0.02371707, 
    0.05483046, 0.07616515, 0.03029847, 0.07132963, 0.04863841, 0.005504836, 
    0.001960447, 0.001966713, 0.008725557, 0.0323761, 0.02341436, 0.08426929, 
    0.01695208,
  0.0886834, 0.006393238, -1.624642e-09, 1.337269e-05, 0.0001487071, 
    -2.068236e-05, 0.0002902934, 7.404307e-08, 0.01333597, 0.0638333, 
    0.03464945, 0.02160867, 0.001590262, 0.003329971, 0.007484001, 
    0.005147147, 0.08308452, 0.1381404, 0.09017851, 0.007880645, 0.09678926, 
    0.02393775, 0.001395967, 0.001709871, 0.06848817, 0.01625923, 
    2.737542e-06, 0.01492575, 0.1716019,
  0.04603515, 0.0305876, 0.0331187, 0.01630275, 0.05016227, 0.1529801, 
    0.0808458, 9.731187e-07, 0.0008537545, 0.06974883, 0.07540977, 
    0.06108309, 0.07455505, 0.08592627, 0.08848644, 0.1077982, 0.09130472, 
    0.1491933, 0.13879, 0.07519375, 0.07367619, 0.1479465, 0.04047408, 
    0.009306131, 0.04424121, 0.1312332, 0.03537689, 0.01235744, 0.05571625,
  0.1322238, 0.04465596, 0.1043025, 0.1036005, 0.149995, 0.1278291, 
    0.01333354, 0.106494, 0.0417254, 0.0341629, 0.08780283, 0.07558393, 
    0.06381851, 0.1521384, 0.2126236, 0.1995235, 0.1769029, 0.1269851, 
    0.03918024, 0.06699002, 0.1007434, 0.09868045, 0.2072954, 0.1988213, 
    0.1892915, 0.1700902, 0.1679424, 0.1015035, 0.08419947,
  0.1602922, 0.1389999, 0.1420346, 0.1676476, 0.2360595, 0.2010984, 0.169426, 
    -0.0002957897, 0, 0.0002268733, -3.56209e-05, 7.163524e-05, 0.04751967, 
    0.07379207, 0.2535626, 0.259799, 0.09788586, 0.0724014, 0.1079618, 
    0.07144113, 0.04413697, 0.07559447, 0.1448602, 0.09388651, 0.1440029, 
    0.1615099, 0.1775885, 0.1763842, 0.193937,
  0.2364151, 0.1868568, 0.1663352, 0.1787399, 0.1467685, 0.1198082, 
    0.05810042, 0.01477888, -0.0001741043, 0, 0, 0, 0.01345569, 0.03173332, 
    0.2330389, 0.2231611, 0.1220771, 0.1427206, 0.07567849, 0.06071942, 
    0.0423579, 0.05484781, 0.01330446, 0.000150326, 0.01774026, 0.04703628, 
    0.09320798, 0.1280241, 0.1781735,
  0.1007698, 0.119365, 0.04803251, 0.0519459, 0.01805932, 0.01403236, 
    0.00673476, 0, 0, 0, 0, 0, -0.0005909011, 0.03536289, 0.1528018, 
    0.1764123, 0.1588418, 0.1190413, 0.1283461, 0.0914906, 0.02369505, 
    0.01634643, 5.803687e-05, 0, 0, 0, -7.730431e-05, 0.1013664, 0.08772331,
  0.01713734, 0.01621191, 0.001306395, 0.0004408071, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.0001027653, 0.008454815, 0.04556835, 0.06112821, 0.06192932, 
    0.04447439, 0.03814764, 0.008228581, -0.000242073, -0.0001375001, 
    0.001285866, -0.0001411717, -3.591325e-05, -3.261209e-07, -0.0001989159, 
    0.01528395,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -4.382915e-10, 0.0002882859, 0.05044032, 
    0.05985595, 0.07145152, 0.1381723, 0.1164013, 0.0418683, 0.004959236, 
    0.002124818, 0.0005127822, 0.05416074, 0.1550981, 0.199015, 0.2328758, 
    0.2052671, 0.06683595, 0.001525718,
  0.06828243, 0.2350626, 0.2207019, 0.2562925, 0.005631754, 0.06793985, 
    0.1260213, 0.04669243, -0.001868084, -0.003244528, 0.0005664529, 
    0.02189422, 0.05966883, 0.1881021, 0.1885007, 0.1750714, 0.1990893, 
    0.1558775, 0.114323, 0.1068193, 0.151719, 0.2643084, 0.2571037, 
    0.2072282, 0.2077358, 0.2570371, 0.2883945, 0.114716, 0.04329471,
  0.1316571, 0.2167999, 0.1869749, 0.2109029, 0.2300688, 0.1943517, 0.182103, 
    0.1615821, 0.2044169, 0.1977009, 0.1828377, 0.233033, 0.2440145, 0.2033, 
    0.2223235, 0.2134081, 0.2006767, 0.1743288, 0.1920376, 0.2251662, 
    0.2104912, 0.2221047, 0.243822, 0.203319, 0.2055616, 0.1819857, 
    0.2360027, 0.1374243, 0.1899121,
  0.1521651, 0.183827, 0.164712, 0.2258577, 0.1762334, 0.178425, 0.1638338, 
    0.1675955, 0.1595029, 0.1174362, 0.1645646, 0.1348498, 0.1735733, 
    0.1893931, 0.1542481, 0.1135964, 0.1085083, 0.1099623, 0.1196179, 
    0.1048153, 0.1430287, 0.1605858, 0.2060349, 0.1350543, 0.09488502, 
    0.1208175, 0.1059534, 0.120236, 0.1712391,
  0.04910717, 0.03270897, 0.02783133, 0.05817706, 0.08473869, 0.05213564, 
    0.09214126, 0.04179306, 0.03862312, 0.03352682, 0.1132696, 0.0814686, 
    0.06805772, 0.05031363, 0.0722909, 0.1315945, 0.1421994, 0.05322176, 
    0.06892309, 0.1299515, 0.09425903, 0.1552969, 0.06080515, 0.02998899, 
    0.07053695, 0.1282813, 0.1859877, 0.1491113, 0.08417971,
  5.525041e-05, -9.641788e-06, 0.09119276, 0.1174719, 0.1685473, 0.06247237, 
    0.05783074, 0.02234694, 0.03052648, 0.007222022, 0.03347394, 0.08431747, 
    0.06223998, 0.008732493, 0.05467965, 0.04760521, 0.06888794, 0.1792696, 
    0.2422037, 0.1258358, 0.04097334, 0.01028737, 0.0001955805, 0.0005660924, 
    0.01656682, 0.1271929, 0.06238678, 0.01243317, 0.002965463,
  9.770132e-08, 0.009074086, 0.1168691, 0.02097377, 0.02449991, 0.003786943, 
    0.03518898, -0.0002225524, 2.922742e-06, -2.080323e-06, 0.02827727, 
    0.01584109, 0.00507975, 0.006881182, 0.05349317, 0.1051694, 0.04433827, 
    0.1667458, 0.00684711, 0.003900002, 3.256636e-05, -5.717622e-10, 
    0.0001051476, 0.0001656352, 0.04571598, 0.1731223, 0.003349789, 
    7.90236e-05, 2.955896e-06,
  7.665616e-05, 0.04320047, 0.08896267, 0.04392052, 0.07055689, 0.02848129, 
    0.08361026, 0.1265351, 0.007013078, 0.01841583, 0.01388485, 0.03352702, 
    0.03288278, 0.1286163, 0.07435437, 0.02853348, 0.01077395, 0.008511174, 
    0.0003236214, 8.422203e-08, 3.553829e-08, 6.209171e-09, 9.698416e-06, 
    0.1215048, 0.1988827, 0.1730957, 0.01154518, 2.15078e-06, 1.04342e-05,
  0.09468033, 0.02282393, 0.01908461, 0.00663778, 0.008520198, 0.02177921, 
    0.06895324, 0.03986301, 0.03231435, 0.2296479, 0.03940277, 0.007299305, 
    0.04668438, 0.08575293, 0.01313856, 0.001705231, 0.0003088183, 
    -7.457685e-05, 0.0001340192, 0.001172608, -2.523281e-08, -7.591005e-09, 
    0.0284135, 0.07063727, 0.02888367, 0.103521, 0.07645546, 0.0002060178, 
    0.0006230699,
  0.0293519, 9.896031e-07, 0.0003439488, 0.002358587, 0.02981217, 
    0.009261619, 9.585837e-05, 0.001869809, 0.06903684, 0.03897604, 
    0.0252881, 0.02810878, 0.06152763, 0.07343062, 0.06675676, 0.02451281, 
    0.06801102, 0.06479012, 0.03896924, 0.08141879, 0.04506824, 0.005575025, 
    0.002010687, 0.003148984, 0.02047736, 0.01988471, 0.0008156231, 
    0.03986902, 0.02316554,
  0.08549673, 0.006587094, 1.218363e-08, 1.433163e-05, 0.0001756596, 
    0.003264219, 0.0004559884, 2.816342e-08, 0.008654967, 0.0618589, 
    0.04584249, 0.01370081, 0.0005047945, 0.002220678, 0.004355972, 
    0.001681212, 0.08794108, 0.1198213, 0.101619, 0.005543302, 0.07961703, 
    0.01667218, 0.001336382, 0.001635753, 0.06531471, 0.006211208, 
    1.450717e-06, 0.009928265, 0.1386029,
  0.02929031, 0.02831534, 0.02889854, 0.01726819, 0.04145949, 0.1582255, 
    0.07661775, 0.0004622825, 0.007521637, 0.0818151, 0.07810515, 0.04759234, 
    0.09512996, 0.08336338, 0.07810365, 0.09953935, 0.08981617, 0.1511577, 
    0.1401244, 0.06697284, 0.07047519, 0.1120475, 0.03522856, 0.005971782, 
    0.0329446, 0.1467619, 0.01162084, 0.008576637, 0.05580383,
  0.1032567, 0.03878219, 0.0943038, 0.159609, 0.1493935, 0.1141311, 
    0.02649172, 0.149649, 0.06042772, 0.1109625, 0.09850811, 0.07527842, 
    0.06604103, 0.1509129, 0.2204625, 0.2056642, 0.1575217, 0.1213991, 
    0.04715074, 0.08269731, 0.1036067, 0.08602663, 0.2085523, 0.199706, 
    0.1929799, 0.1470346, 0.1601336, 0.09013776, 0.1027455,
  0.1854108, 0.1456142, 0.1516975, 0.1710567, 0.2429458, 0.2181592, 
    0.2724871, -0.001002007, 0.003215545, 0.004136572, 0.002437871, 
    0.01229847, 0.1522988, 0.153001, 0.2767572, 0.2660973, 0.07981824, 
    0.07794825, 0.1038341, 0.07361685, 0.07388016, 0.1117755, 0.2086931, 
    0.1627437, 0.1536057, 0.1792194, 0.198974, 0.2025057, 0.1941403,
  0.2731553, 0.2277061, 0.2044269, 0.2139926, 0.1929259, 0.1821123, 0.138892, 
    0.1531036, 0.09371216, 0.03684176, -6.356068e-06, -6.289605e-05, 
    0.015878, 0.06032669, 0.2825865, 0.2461218, 0.1530446, 0.172542, 
    0.1264906, 0.1499828, 0.1010229, 0.09823655, 0.08306352, 0.05225497, 
    0.04586517, 0.09763087, 0.1734792, 0.2026443, 0.2358714,
  0.243081, 0.2513489, 0.1787991, 0.1544456, 0.08147754, 0.06201902, 
    0.06311707, 0.02465491, -5.843054e-05, 0, 0, -2.461826e-05, 0.01115665, 
    0.1136203, 0.1780335, 0.1955252, 0.2180329, 0.190975, 0.2068557, 
    0.1853069, 0.093254, 0.03821265, 0.01537907, -2.384365e-05, 0.0005379893, 
    -0.0001438675, -0.0003326633, 0.1757989, 0.2316415,
  0.1327761, 0.09842232, 0.05530159, 0.02387972, 0.0159293, 0.004008373, 
    0.002513378, 0.007679749, 0.01227958, 0.01007662, 0.01304636, 0.01208525, 
    0.0135252, 0.03685769, 0.09330061, 0.09327034, 0.09600337, 0.09125943, 
    0.08972802, 0.07986607, 0.0774127, 0.06427535, 0.01263599, 0.0004723419, 
    0.002612423, 0.0001848003, -0.0006507433, 0.001726583, 0.06807328,
  0.003990239, 0.002360163, 0.0007300873, -0.0008999886, -0.002530065, 
    -0.004160141, -0.005790216, -0.0002519356, -0.0001135386, 2.485845e-05, 
    0.0001632555, 0.0003016525, 0.0004400495, 0.0005784465, 0.003390337, 
    0.00341277, 0.003435203, 0.003457636, 0.003480069, 0.003502502, 
    0.003524935, -0.006913685, -0.005444439, -0.003975193, -0.002505947, 
    -0.001036701, 0.0004325454, 0.001901791, 0.0052943,
  -0.001139022, -2.046406e-05, 0, 0, 0, -0.0006758879, 0, 0, 0, 0, 0, 
    -2.399728e-05, 0.00239515, 0.07882516, 0.07126889, 0.1258411, 0.1696257, 
    0.1697955, 0.1103822, 0.03275169, 0.0202423, 0.03977493, 0.1373487, 
    0.1336874, 0.1832106, 0.2271752, 0.2471205, 0.1155661, 0.02554919,
  0.06533501, 0.2300999, 0.2294332, 0.3264087, 0.06275953, 0.1368529, 
    0.1958865, 0.07174329, 0.006235706, 0.03784668, 0.01276804, 0.03841843, 
    0.1334302, 0.2125449, 0.2265066, 0.2126219, 0.2306272, 0.2022461, 
    0.1346471, 0.1361215, 0.159078, 0.2686701, 0.2864582, 0.2499526, 
    0.2260912, 0.2553743, 0.2775495, 0.1145122, 0.04231213,
  0.1228263, 0.2240393, 0.2110861, 0.2354367, 0.2377368, 0.2009756, 
    0.1891661, 0.1668932, 0.2112143, 0.2240671, 0.240435, 0.28044, 0.2441746, 
    0.204616, 0.2296818, 0.2154759, 0.1968499, 0.1858603, 0.2254899, 
    0.2584325, 0.244862, 0.2711472, 0.268854, 0.2112025, 0.2212138, 
    0.2075691, 0.2246194, 0.1389591, 0.1977788,
  0.1561813, 0.1776106, 0.1688515, 0.2137991, 0.162361, 0.175649, 0.145585, 
    0.1667065, 0.1774843, 0.1412738, 0.1630313, 0.145336, 0.1666669, 
    0.1811112, 0.1549307, 0.1030462, 0.0846833, 0.1103528, 0.1157315, 
    0.09908962, 0.1363715, 0.1453051, 0.1793056, 0.1412174, 0.08861261, 
    0.1199087, 0.1192309, 0.1300592, 0.1712703,
  0.05389105, 0.02617789, 0.02571757, 0.06767813, 0.07827244, 0.05398549, 
    0.07290966, 0.03386662, 0.03346508, 0.0282819, 0.1146775, 0.07834887, 
    0.06166764, 0.04655004, 0.08054284, 0.1303198, 0.1414936, 0.03658292, 
    0.05618617, 0.1268474, 0.08992091, 0.135938, 0.05232078, 0.02171556, 
    0.064482, 0.1228732, 0.1762165, 0.1482091, 0.104139,
  -0.0001565681, 1.043303e-05, 0.09073874, 0.08510998, 0.1483798, 0.05695553, 
    0.0537779, 0.009051426, 0.0128791, 0.001172692, 0.04005047, 0.06936099, 
    0.06225067, 0.004639624, 0.04366501, 0.02573768, 0.05158934, 0.1638963, 
    0.2165117, 0.07106167, 0.01531545, 0.008777521, 0.0001563745, 
    2.725544e-06, 0.01622357, 0.1091828, 0.06767795, 0.01488311, 0.00588703,
  2.452205e-07, 0.007864556, 0.09991639, 0.0305084, 0.02051191, 0.003186332, 
    0.03935164, 0.001969973, 5.977446e-08, 1.288289e-05, 0.02056053, 
    0.01100306, 0.007395769, 0.01485295, 0.04181839, 0.09736323, 0.05117368, 
    0.1570721, 0.009694338, 0.00364903, 3.163381e-05, -7.216718e-10, 
    4.88802e-06, 0.0003283923, 0.05164923, 0.1426735, 0.002887252, 
    0.0002247306, 1.784818e-07,
  0.001127589, 0.04407576, 0.06352714, 0.04202233, 0.07071028, 0.02469416, 
    0.08650072, 0.1174106, 0.005185355, 0.02000929, 0.01659241, 0.02981075, 
    0.02706224, 0.1118088, 0.07486481, 0.03116015, 0.01352376, 0.006767894, 
    0.001012332, 3.409951e-08, 1.080815e-09, -2.229146e-12, 0.0005887869, 
    0.1058361, 0.2004171, 0.1489614, 0.01061607, -8.226957e-07, 0.0001433424,
  0.234577, 0.01482605, 0.0267632, 0.007023375, 0.01594191, 0.01571582, 
    0.06300125, 0.03000865, 0.03421107, 0.2086456, 0.0381388, 0.007001762, 
    0.03695622, 0.07501595, 0.01295243, 0.002683687, 9.276556e-05, 
    0.0001352241, 0.00070551, 0.0009338682, 3.944132e-07, -1.06323e-06, 
    0.04572133, 0.09253547, 0.03946105, 0.09510218, 0.05412004, 0.001852805, 
    0.03308034,
  0.03000078, 6.75856e-07, 0.01118198, 0.00153291, 0.02944021, 0.008699995, 
    0.0001157643, 0.001372675, 0.06806897, 0.03931188, 0.02624943, 0.0337356, 
    0.05635601, 0.06888888, 0.05631125, 0.02580069, 0.08893225, 0.03946424, 
    0.0547136, 0.07947833, 0.04357571, 0.00588277, 0.004412136, 0.005471975, 
    0.03195312, 0.01948073, 0.002025353, 0.01452229, 0.05436238,
  0.08889816, 7.356183e-05, -6.18324e-09, 1.451734e-05, 0.0003817468, 
    0.001513746, 0.0004955249, 1.923742e-09, 0.00341909, 0.05780608, 
    0.05915273, 0.01099033, 0.0007574628, 0.0009705552, 0.00059567, 
    0.003635405, 0.07911745, 0.09308527, 0.07565927, 0.004830504, 0.06376725, 
    0.01102263, 0.003483019, 0.002008678, 0.06370642, 0.003298485, 
    5.134357e-08, 0.001946506, 0.1283545,
  0.02999852, 0.02937385, 0.02391755, 0.02709077, 0.04008627, 0.1612006, 
    0.07905309, 0.002688678, 0.03459906, 0.07603334, 0.08888181, 0.05642824, 
    0.09160676, 0.09160749, 0.05893591, 0.09202968, 0.08159727, 0.1553573, 
    0.1280918, 0.07646279, 0.05923378, 0.09220458, 0.03178482, 0.003895437, 
    0.03454312, 0.1025083, 0.01021076, 0.009056931, 0.03926798,
  0.09163989, 0.03850273, 0.102293, 0.1666765, 0.1508114, 0.09197237, 
    0.07510433, 0.1571063, 0.0758135, 0.1222963, 0.08630943, 0.06459745, 
    0.076215, 0.1614648, 0.2183952, 0.1878704, 0.1515093, 0.1214739, 
    0.07388873, 0.1177659, 0.1122099, 0.08255541, 0.2216211, 0.1948686, 
    0.1943209, 0.1499354, 0.1495997, 0.08498175, 0.1193809,
  0.1865364, 0.155128, 0.1834602, 0.1769474, 0.2151996, 0.2126578, 0.2708162, 
    0.05622097, 0.04969931, 0.05092171, 0.04091543, 0.0390893, 0.231214, 
    0.2357245, 0.2793493, 0.2586766, 0.07396695, 0.08326165, 0.1158408, 
    0.09983662, 0.09787578, 0.1322763, 0.2188845, 0.1809629, 0.1534991, 
    0.1847807, 0.2084271, 0.2164273, 0.2044871,
  0.3125999, 0.2605316, 0.2466239, 0.2310318, 0.2027143, 0.2851511, 
    0.2528586, 0.2949392, 0.2031572, 0.1294186, 0.0443817, -0.000277109, 
    0.03075937, 0.1278556, 0.3370344, 0.2738095, 0.1751011, 0.2087515, 
    0.1606599, 0.2035451, 0.1713919, 0.1749277, 0.1355882, 0.1569458, 
    0.1073717, 0.2076819, 0.1838608, 0.2442217, 0.2675408,
  0.2499291, 0.3560562, 0.2464603, 0.2284575, 0.1817243, 0.1616468, 
    0.2238616, 0.1307998, 0.06150441, 0.05170617, 0.01620429, 0.01837752, 
    0.1082524, 0.2249647, 0.2320109, 0.2907419, 0.2796639, 0.2425825, 
    0.2644494, 0.2442461, 0.1409616, 0.05924603, 0.05810136, -0.00132204, 
    0.003366489, 0.001347867, 0.001828424, 0.2083257, 0.2565329,
  0.1602256, 0.184851, 0.0924677, 0.03621165, 0.0203563, 0.02019269, 
    0.02178503, 0.02580382, 0.05825746, 0.0799417, 0.08395804, 0.1062235, 
    0.08764321, 0.1182418, 0.1503113, 0.1154287, 0.09378588, 0.09229525, 
    0.08868729, 0.09484854, 0.08678689, 0.1115674, 0.03566495, -0.0003096948, 
    0.00292359, 0.0003966663, 0.0001758043, 0.01911873, 0.0981142,
  0.06727315, 0.06590822, 0.06454328, 0.06317835, 0.06181341, 0.06044848, 
    0.05908354, 0.06407852, 0.06107694, 0.05807535, 0.05507377, 0.05207218, 
    0.0490706, 0.04606901, 0.02471418, 0.02827971, 0.03184524, 0.03541077, 
    0.0389763, 0.04254184, 0.04610737, 0.07115003, 0.07195102, 0.072752, 
    0.07355299, 0.07435398, 0.07515497, 0.07595596, 0.0683651,
  0.03966309, -0.001063082, -0.0001946042, 0, 0.001579147, 0.003736655, 
    3.465553e-05, 0, 0, 0, -0.0001385093, 0.002947371, 0.02040004, 0.1292218, 
    0.06450079, 0.1344197, 0.1610285, 0.2037986, 0.1781977, 0.1264294, 
    0.1071818, 0.1357589, 0.2171769, 0.1304213, 0.1729774, 0.2186925, 
    0.2515773, 0.1696583, 0.09826604,
  0.06976331, 0.2045381, 0.2210599, 0.311024, 0.1868372, 0.1819283, 
    0.2189261, 0.07585524, 0.05140887, 0.07596651, 0.05681515, 0.05918045, 
    0.1903351, 0.2242731, 0.2409639, 0.2130283, 0.2480349, 0.2278609, 
    0.1524726, 0.1506549, 0.16252, 0.2554579, 0.2797156, 0.233321, 0.2381657, 
    0.2303691, 0.2662195, 0.1095953, 0.04349333,
  0.125245, 0.230278, 0.2273531, 0.2345544, 0.2443417, 0.2102503, 0.2037022, 
    0.1782295, 0.2116498, 0.2304419, 0.282503, 0.2674423, 0.2627065, 
    0.2040839, 0.2653728, 0.2153201, 0.1989928, 0.2119531, 0.2563493, 
    0.2677668, 0.2614856, 0.2793826, 0.2947356, 0.212393, 0.2157829, 
    0.2492473, 0.2271461, 0.1488646, 0.1894654,
  0.1500628, 0.176952, 0.1685677, 0.2008904, 0.1601143, 0.1564403, 0.1307995, 
    0.1711179, 0.1755327, 0.1578343, 0.1575186, 0.1353261, 0.1431914, 
    0.18343, 0.1420251, 0.1128364, 0.09217534, 0.1006173, 0.1218033, 
    0.08656854, 0.160511, 0.1462937, 0.1737363, 0.1239056, 0.08557073, 
    0.1209547, 0.1156849, 0.1300283, 0.1743367,
  0.048716, 0.01997038, 0.02193406, 0.07869601, 0.07523928, 0.04969458, 
    0.07646257, 0.03109821, 0.02660392, 0.04281881, 0.1129229, 0.0754725, 
    0.05821323, 0.04518865, 0.07227685, 0.1364172, 0.1260194, 0.02367513, 
    0.0407816, 0.1180533, 0.07825646, 0.1338338, 0.04726776, 0.0172568, 
    0.06850547, 0.1173647, 0.1646983, 0.1239938, 0.09162466,
  -6.273694e-05, 4.463409e-05, 0.08757159, 0.06149476, 0.1340493, 0.06687059, 
    0.05549277, 0.005340375, 0.007870398, 0.000925109, 0.05075226, 
    0.05636992, 0.0562152, 0.002524406, 0.03809404, 0.01914764, 0.04475023, 
    0.1666217, 0.1580835, 0.05057513, 0.0154831, 0.006258303, 2.947341e-05, 
    -3.369764e-08, 0.01943627, 0.08702671, 0.09652825, 0.01731679, 0.004558417,
  2.180471e-05, 0.01772523, 0.09213598, 0.03093361, 0.01641764, 0.00446637, 
    0.05192397, 0.005506143, 3.784826e-07, 0.0002049883, 0.02886957, 
    0.01593667, 0.01129926, 0.01423898, 0.04053754, 0.1096728, 0.05504008, 
    0.1516706, 0.01055667, 0.00375445, 3.514884e-06, 2.108697e-10, 
    4.926136e-06, 0.0007921652, 0.06458603, 0.1462561, 0.002078016, 
    1.385926e-05, 1.369642e-07,
  0.003355326, 0.0554035, 0.05359531, 0.04824051, 0.06656925, 0.02597972, 
    0.09769613, 0.122229, 0.004342271, 0.02432879, 0.01637007, 0.03317, 
    0.0245729, 0.116145, 0.07328364, 0.0359159, 0.01610973, 0.007168268, 
    0.001758646, 4.236254e-07, 9.905115e-09, -1.587887e-06, 0.0007233606, 
    0.09537674, 0.2317585, 0.1283416, 0.008112269, 0.0002199646, 0.00661356,
  0.3923626, 0.01512463, 0.05098205, 0.009104413, 0.03957753, 0.01573688, 
    0.07690959, 0.03026666, 0.03523652, 0.1910702, 0.03682435, 0.005324435, 
    0.03925228, 0.07496011, 0.01366841, 0.006708964, 9.45195e-05, 
    0.0007910891, 0.0001080306, 9.38455e-05, 8.336202e-07, -0.0001520685, 
    0.08957538, 0.09963515, 0.04658103, 0.07896756, 0.0366772, 0.02114331, 
    0.1424824,
  0.003890483, 5.485513e-07, 0.01708103, 0.001532005, 0.02647214, 
    0.008108701, 0.0001919489, 0.001140094, 0.06802757, 0.04207004, 
    0.02717717, 0.04055999, 0.05097836, 0.06426387, 0.04956849, 0.03312185, 
    0.1161036, 0.02690835, 0.05663919, 0.08565335, 0.04918043, 0.009987785, 
    0.003941973, 0.007620947, 0.03763935, 0.01840083, 0.00947476, 
    0.009343605, 0.01743311,
  0.08172306, 5.281544e-06, -5.587325e-09, 1.391879e-05, 0.0004037415, 
    0.0003038131, 0.0001862093, 6.642246e-05, 0.000207733, 0.07182639, 
    0.07840829, 0.01385982, 0.0005012672, 0.000648334, 0.0006690691, 
    0.00230753, 0.07028171, 0.08627638, 0.04464925, 0.00193564, 0.0391318, 
    0.009025618, 0.00311641, 0.002660801, 0.06148264, 0.002729871, 
    1.412877e-06, 4.435835e-06, 0.09134185,
  0.03282387, 0.02300178, 0.0189914, 0.03299592, 0.03663881, 0.1445955, 
    0.07729201, 0.01468102, 0.07843771, 0.08493094, 0.1024049, 0.08081091, 
    0.1048692, 0.09224186, 0.06074998, 0.09433649, 0.08810834, 0.1365948, 
    0.1113582, 0.05736459, 0.05148409, 0.07323737, 0.02650869, 0.001714517, 
    0.03576758, 0.08175793, 0.006506926, 0.007920882, 0.02878856,
  0.07490087, 0.03858435, 0.1087222, 0.165962, 0.1536579, 0.08416355, 
    0.1021781, 0.1514305, 0.07869516, 0.1125778, 0.08025473, 0.06336025, 
    0.07895759, 0.1467093, 0.2240046, 0.1718216, 0.1515408, 0.1016622, 
    0.07223427, 0.1339014, 0.1172053, 0.07891274, 0.2120435, 0.1769485, 
    0.1792711, 0.143278, 0.1503996, 0.06805101, 0.1097195,
  0.1744858, 0.1664464, 0.1458282, 0.1799094, 0.2115781, 0.1711712, 
    0.2764485, 0.1237623, 0.1148179, 0.1088578, 0.05128691, 0.06733566, 
    0.2269171, 0.2341094, 0.2815033, 0.2400546, 0.07338994, 0.07578494, 
    0.1326225, 0.1789812, 0.1222866, 0.1521416, 0.21354, 0.1854444, 
    0.1571164, 0.1854471, 0.2035291, 0.2246734, 0.1857924,
  0.2865953, 0.296415, 0.2377443, 0.2304242, 0.2399498, 0.3458222, 0.2977982, 
    0.3394802, 0.2398119, 0.1896546, 0.1438953, 0.0007356447, 0.09308617, 
    0.1512859, 0.3451869, 0.2736347, 0.1900535, 0.2119654, 0.2179772, 
    0.2526034, 0.1992415, 0.2040413, 0.184416, 0.2796714, 0.1159103, 
    0.2369237, 0.1978875, 0.2798016, 0.2651927,
  0.2640347, 0.3423505, 0.3118294, 0.2622723, 0.2592783, 0.2570383, 
    0.3351065, 0.3023766, 0.2026388, 0.1840946, 0.1103959, 0.1307521, 
    0.2092992, 0.2647093, 0.28225, 0.3094599, 0.3021996, 0.2864705, 0.293371, 
    0.2479013, 0.166983, 0.0928572, 0.08249252, 0.007478716, 0.04805413, 
    0.0142472, 0.004452249, 0.1995478, 0.2851644,
  0.2806033, 0.3017316, 0.1859996, 0.05903375, 0.03396276, 0.0693953, 
    0.0897109, 0.1222892, 0.1656831, 0.1998507, 0.2011674, 0.1969775, 
    0.2204502, 0.2378469, 0.2520364, 0.1476048, 0.148376, 0.1380842, 
    0.09351512, 0.1101783, 0.09078199, 0.1227471, 0.09301347, 0.009920505, 
    0.0171646, 0.004014751, 0.005766223, 0.006560443, 0.1902665,
  0.08475678, 0.08434079, 0.08392479, 0.0835088, 0.08309281, 0.08267681, 
    0.08226082, 0.08785783, 0.08745202, 0.0870462, 0.08664039, 0.08623457, 
    0.08582876, 0.08542294, 0.08130479, 0.08321545, 0.0851261, 0.08703676, 
    0.08894742, 0.09085807, 0.09276873, 0.0947281, 0.09363925, 0.0925504, 
    0.09146155, 0.0903727, 0.08928385, 0.088195, 0.08508957,
  0.1126059, 0.01425214, 0.007613398, 0.01449402, 0.02701701, 0.007654302, 
    0.0005907958, 0.01032371, 0.009467029, 0.002764474, 0.01067922, 
    0.05023815, 0.05499223, 0.139388, 0.07645407, 0.1550265, 0.1517758, 
    0.1955398, 0.2492831, 0.159948, 0.2163634, 0.3245367, 0.2329569, 
    0.1147977, 0.1580444, 0.2182256, 0.2457571, 0.1661399, 0.101936,
  0.07154284, 0.1907383, 0.2194, 0.2999404, 0.3176745, 0.2158697, 0.2270441, 
    0.1362685, 0.08065566, 0.1187129, 0.09390386, 0.08769207, 0.205916, 
    0.2303534, 0.253253, 0.2142098, 0.2534429, 0.2420343, 0.1762167, 
    0.1560905, 0.1648297, 0.2560937, 0.2779722, 0.2389389, 0.2525486, 
    0.2079977, 0.2638681, 0.09472691, 0.04140479,
  0.1268818, 0.2132403, 0.237755, 0.245822, 0.238801, 0.2231537, 0.2100559, 
    0.1771336, 0.2147887, 0.2279091, 0.2780986, 0.2711398, 0.2765234, 
    0.2156129, 0.2734268, 0.2088518, 0.2137954, 0.2172424, 0.2564475, 
    0.2545453, 0.2768519, 0.2607279, 0.2809612, 0.2351103, 0.2429078, 
    0.2654583, 0.2352834, 0.1529145, 0.197376,
  0.1701204, 0.1728104, 0.168208, 0.2041262, 0.157703, 0.1521484, 0.1266132, 
    0.157875, 0.1844403, 0.1862325, 0.1604612, 0.139107, 0.1504753, 
    0.1871065, 0.1380119, 0.1205411, 0.08837456, 0.09820368, 0.127105, 
    0.09519899, 0.1278632, 0.1426401, 0.1597602, 0.117226, 0.09793386, 
    0.1297568, 0.1245841, 0.1337626, 0.1759485,
  0.04883474, 0.01891296, 0.02262843, 0.08503902, 0.08348738, 0.05313718, 
    0.06838222, 0.03527883, 0.04185696, 0.03451418, 0.1069627, 0.06490052, 
    0.05388355, 0.03924911, 0.07285225, 0.1436246, 0.1071696, 0.01531888, 
    0.04019136, 0.1149937, 0.07534365, 0.1169015, 0.04373441, 0.01444908, 
    0.0745681, 0.1193556, 0.1502722, 0.1104998, 0.0809184,
  0.0008662273, -9.432658e-06, 0.1013276, 0.05627242, 0.1274915, 0.06738549, 
    0.05773789, 0.00219081, 0.0006351347, 0.001602706, 0.05263945, 
    0.06078258, 0.06610739, 0.004641879, 0.03359004, 0.01050606, 0.04241161, 
    0.1627135, 0.1271062, 0.04310642, 0.01951731, 0.003799888, 8.889735e-06, 
    3.822397e-06, 0.03622178, 0.08131649, 0.1200445, 0.01369305, 0.002479243,
  0.01245099, 0.05046882, 0.09877551, 0.03090161, 0.01689854, 0.007639392, 
    0.07629317, 0.002888202, 3.699362e-07, 1.228526e-05, 0.0385031, 
    0.03764907, 0.01011055, 0.0182719, 0.04135889, 0.1263875, 0.04658334, 
    0.1481177, 0.01350136, 0.00431906, -6.186439e-06, 7.188015e-10, 
    1.121467e-05, 0.001321838, 0.0833874, 0.1761632, 0.001336297, 
    3.628508e-06, 1.611774e-07,
  0.006281313, 0.1057705, 0.07092963, 0.07171807, 0.07522092, 0.03001213, 
    0.1100116, 0.1265798, 0.008429323, 0.0340614, 0.02263771, 0.03920321, 
    0.03406138, 0.1326368, 0.08269262, 0.04945979, 0.02035967, 0.00860061, 
    0.003438027, 7.510373e-06, 5.29118e-08, -2.683011e-07, 0.003379288, 
    0.1067572, 0.2726641, 0.1296237, 0.005409838, 0.0007694046, 0.001281817,
  0.4211332, 0.02887733, 0.07794567, 0.01429555, 0.0385949, 0.01975025, 
    0.09070067, 0.03507312, 0.04979709, 0.1938329, 0.04381934, 0.008199789, 
    0.05424678, 0.0805208, 0.01871916, 0.008595537, 5.335414e-05, 
    0.003200348, -6.376435e-05, 0.0001656546, 0.001676523, 0.01960539, 
    0.1436818, 0.1340368, 0.06065661, 0.06852131, 0.03439352, 0.02636878, 
    0.1200529,
  -6.204436e-05, 4.87142e-07, 0.01988005, 0.002729773, 0.03207142, 
    0.01018033, 0.0001358782, 0.001197695, 0.07103605, 0.04831784, 
    0.03501862, 0.05103766, 0.05103331, 0.07234085, 0.05498635, 0.05573151, 
    0.1218792, 0.03137689, 0.06873769, 0.09598774, 0.05735296, 0.01081945, 
    0.004485561, 0.01298449, 0.04205106, 0.01595879, 0.02701476, 0.01475769, 
    0.01950079,
  0.06592971, 1.207302e-05, 3.471009e-08, 8.007071e-06, 0.002060008, 
    0.001517199, 0.0002803006, 5.390619e-05, 1.088008e-05, 0.07071891, 
    0.08149003, 0.02299446, 0.0003500449, 0.0001947699, 0.0008310603, 
    0.005045163, 0.06089822, 0.08398288, 0.03375526, 0.001262464, 0.02448094, 
    0.009191389, 0.002704844, 0.003853971, 0.05781787, 0.003216937, 
    5.993266e-05, 8.448048e-07, 0.0680912,
  0.01016453, 0.02577545, 0.01420345, 0.02531976, 0.03863296, 0.1380817, 
    0.08227102, 0.03961388, 0.1106496, 0.103012, 0.1171617, 0.09462631, 
    0.1123483, 0.08499213, 0.05698965, 0.113069, 0.09292016, 0.1258413, 
    0.09226098, 0.05236739, 0.0562791, 0.06677889, 0.02323346, 0.0120504, 
    0.03794885, 0.0695755, 0.0108508, 0.005140598, 0.02964744,
  0.06212771, 0.03567863, 0.1114488, 0.1658166, 0.1579151, 0.06996746, 
    0.117803, 0.1304224, 0.07206928, 0.1147416, 0.0758651, 0.07817944, 
    0.07525164, 0.150484, 0.2077137, 0.1596894, 0.1513622, 0.07530253, 
    0.06663903, 0.1374021, 0.1322393, 0.07748955, 0.2006937, 0.1724797, 
    0.1659171, 0.1425457, 0.1469731, 0.07548588, 0.1080885,
  0.1759656, 0.1448803, 0.1337719, 0.174931, 0.1833815, 0.1818777, 0.2672748, 
    0.1677895, 0.1540729, 0.1088715, 0.05202456, 0.06791328, 0.2546448, 
    0.224272, 0.270341, 0.2304005, 0.08434884, 0.0704325, 0.1090574, 
    0.2513152, 0.1302987, 0.1511886, 0.188151, 0.2154565, 0.1621045, 
    0.1836794, 0.2156918, 0.2037434, 0.1710017,
  0.2920603, 0.2875259, 0.2399906, 0.2157446, 0.2596561, 0.3567441, 
    0.2985374, 0.3263927, 0.2701097, 0.2496051, 0.2159996, 0.0402242, 
    0.1959301, 0.2199652, 0.3440992, 0.2567909, 0.1856506, 0.2071061, 
    0.2721473, 0.2400981, 0.1963328, 0.1978181, 0.191247, 0.3449389, 
    0.1467131, 0.2335937, 0.1930218, 0.2750836, 0.271073,
  0.2752811, 0.3143134, 0.335232, 0.2682197, 0.2791465, 0.2823935, 0.409398, 
    0.3538556, 0.2875661, 0.241017, 0.1939683, 0.1724554, 0.2394528, 
    0.2873051, 0.2966578, 0.3002481, 0.2982534, 0.3300424, 0.3035663, 
    0.2494619, 0.1764039, 0.1231147, 0.138863, -0.001341661, 0.2430471, 
    0.059916, 0.07766833, 0.186162, 0.3057404,
  0.281789, 0.3330047, 0.1748661, 0.0701409, 0.04560691, 0.1012451, 
    0.1129699, 0.1038447, 0.1213563, 0.2477763, 0.2803694, 0.2495882, 
    0.2212656, 0.2581224, 0.2698271, 0.1729408, 0.1684839, 0.1946949, 
    0.1673681, 0.1513212, 0.1172485, 0.1788544, 0.1419962, 0.07347963, 
    0.06870464, 0.01394004, 0.04240727, 0.08848512, 0.2045432,
  0.1425587, 0.1371274, 0.1316961, 0.1262648, 0.1208335, 0.1154022, 
    0.1099709, 0.1297769, 0.1322683, 0.1347597, 0.1372511, 0.1397425, 
    0.1422339, 0.1447253, 0.1242124, 0.1290291, 0.1338458, 0.1386625, 
    0.1434792, 0.148296, 0.1531127, 0.1933501, 0.1914733, 0.1895965, 
    0.1877196, 0.1858428, 0.183966, 0.1820892, 0.1469038,
  0.1224593, 0.1008512, 0.01206676, 0.0184086, 0.03660408, 0.002450722, 
    -5.422613e-06, 0.007152546, 0.02740856, 0.03336051, 0.07835878, 
    0.1092943, 0.101617, 0.1521276, 0.04690773, 0.1727488, 0.1509384, 
    0.2052342, 0.2210055, 0.2104301, 0.2157951, 0.3500561, 0.2361342, 
    0.1194958, 0.1506286, 0.2142211, 0.2396155, 0.1680785, 0.0998005,
  0.09474145, 0.2198275, 0.2405236, 0.3402818, 0.3933396, 0.2602266, 
    0.2176992, 0.2166196, 0.1196074, 0.1936881, 0.1798121, 0.1546191, 
    0.208295, 0.2236457, 0.2199152, 0.2267787, 0.2431242, 0.2643053, 
    0.2222793, 0.2066864, 0.2028905, 0.3262148, 0.3727521, 0.3307368, 
    0.2673748, 0.1918554, 0.2389329, 0.08411425, 0.05079998,
  0.1337279, 0.2203542, 0.2999939, 0.2365741, 0.2418773, 0.2242524, 
    0.2053374, 0.2075107, 0.2193006, 0.206386, 0.2983476, 0.3120526, 
    0.2764348, 0.2175068, 0.204603, 0.2231418, 0.2253187, 0.222877, 
    0.2752109, 0.2906229, 0.2872671, 0.3110608, 0.3257226, 0.2253698, 
    0.2714631, 0.2701033, 0.233401, 0.1617968, 0.2194321,
  0.1846996, 0.1688236, 0.1518929, 0.1945841, 0.1519512, 0.1517031, 
    0.1342811, 0.1620789, 0.1785893, 0.1875649, 0.1731086, 0.156871, 
    0.1524531, 0.1950277, 0.1418741, 0.1192573, 0.08860109, 0.09291644, 
    0.1272747, 0.1002848, 0.1729687, 0.1322626, 0.1422365, 0.1161011, 
    0.1193866, 0.1278527, 0.1368757, 0.1308884, 0.1763864,
  0.03859322, 0.02319843, 0.0305386, 0.09345075, 0.09699239, 0.05138769, 
    0.07125582, 0.05535579, 0.04916299, 0.03677354, 0.08383605, 0.05882284, 
    0.05269234, 0.03790973, 0.08501504, 0.1327015, 0.1057873, 0.01303925, 
    0.04197627, 0.1152507, 0.0769675, 0.1006643, 0.04111314, 0.01010278, 
    0.08704814, 0.1282756, 0.1512753, 0.1114209, 0.07630505,
  0.002956114, 4.839599e-07, 0.1243147, 0.05307984, 0.1165702, 0.07145715, 
    0.06233214, 0.006454988, 1.510739e-05, 0.00685575, 0.04681574, 
    0.05105546, 0.08423715, 0.004848821, 0.04280196, 0.005703134, 0.03715971, 
    0.1681649, 0.1520597, 0.0417117, 0.02005443, 0.00189791, 7.566747e-06, 
    8.381524e-06, 0.04399006, 0.07752797, 0.1064705, 0.006966125, 0.001778921,
  0.005642916, 0.06921447, 0.1209707, 0.03692846, 0.01722459, 0.01158012, 
    0.09047917, 0.0003279038, 4.78444e-07, 0.002102867, 0.04973332, 
    0.06867824, 0.006054637, 0.03016426, 0.0456812, 0.1610234, 0.04925638, 
    0.1525409, 0.02351524, 0.006984742, -1.417746e-05, 7.559699e-10, 
    1.023018e-05, 0.000754445, 0.1016892, 0.2021373, 0.005200557, 
    5.12989e-06, 2.467928e-07,
  0.01853302, 0.1423986, 0.1119529, 0.09793544, 0.08123294, 0.03472444, 
    0.1318326, 0.1436577, 0.0145749, 0.04610804, 0.0333336, 0.0532306, 
    0.03505774, 0.145475, 0.1021179, 0.04717466, 0.02019895, 0.009143962, 
    0.007611872, 0.0002559993, 2.905734e-08, -2.069631e-05, 0.00742741, 
    0.1441126, 0.3184122, 0.127005, 0.007100657, 6.2064e-05, 0.003877195,
  0.4378321, 0.0526341, 0.09336591, 0.02048217, 0.04212787, 0.02941594, 
    0.1025899, 0.04263884, 0.1000214, 0.2315316, 0.05085547, 0.01005768, 
    0.07172694, 0.08939134, 0.02373411, 0.01299214, 0.0001114826, 
    -0.0001003398, -3.253605e-05, 0.005489613, 0.01331991, 0.04025423, 
    0.2072649, 0.1662781, 0.08814201, 0.07434782, 0.03492736, 0.02564042, 
    0.07106175,
  6.291953e-07, 3.071225e-06, 0.004916965, 0.006700892, 0.03437134, 
    0.01404482, 0.0001737902, 0.001492622, 0.08058279, 0.05405604, 
    0.04602606, 0.06081433, 0.0564125, 0.07144479, 0.07160784, 0.05883535, 
    0.1083143, 0.04849174, 0.07737452, 0.1031465, 0.07312962, 0.009428709, 
    0.005523511, 0.01837174, 0.06166174, 0.01473595, 0.02124297, 0.007596109, 
    0.008492161,
  0.02798569, 6.759513e-06, 7.324267e-08, 1.021968e-05, 0.01215482, 
    0.006967243, 0.0003885791, 9.745229e-07, 2.920504e-05, 0.08166358, 
    0.0748738, 0.03661354, 0.0002886844, 0.0004656666, 0.001415316, 
    0.005865328, 0.05601074, 0.09774669, 0.03230619, 0.0008924195, 
    0.02764024, 0.0120257, 0.002862669, 0.006229341, 0.05765062, 0.006994743, 
    0.0008502609, -1.824609e-06, 0.05109694,
  0.0008203969, 0.0213182, 0.01223904, 0.02409577, 0.04555869, 0.1400441, 
    0.07270028, 0.05547733, 0.1476465, 0.1532912, 0.1193346, 0.09170125, 
    0.1074882, 0.0873896, 0.06057859, 0.1149234, 0.09909043, 0.1164348, 
    0.08868363, 0.05108612, 0.07745047, 0.06544904, 0.02394882, 0.0143684, 
    0.05231307, 0.07536251, 0.01593611, 0.007539247, 0.04280106,
  0.05725009, 0.04141591, 0.134926, 0.1675157, 0.1466205, 0.07858832, 
    0.1355692, 0.1070099, 0.05485539, 0.118495, 0.05368171, 0.08712727, 
    0.08361152, 0.1612419, 0.2059086, 0.1386993, 0.1375891, 0.06319772, 
    0.09272645, 0.1514635, 0.1544683, 0.08518726, 0.1884384, 0.1656106, 
    0.1671968, 0.1524284, 0.1457482, 0.06798458, 0.1222835,
  0.1779032, 0.1537062, 0.1159596, 0.1370596, 0.1568004, 0.1706888, 
    0.2516649, 0.16816, 0.1776178, 0.105385, 0.05390345, 0.06029079, 
    0.2473448, 0.2093604, 0.2672226, 0.2160312, 0.08218381, 0.06667287, 
    0.1102311, 0.2911288, 0.1330925, 0.1405361, 0.1812947, 0.1922033, 
    0.1536974, 0.1693552, 0.2298244, 0.2212203, 0.1893935,
  0.3188591, 0.2950285, 0.2465742, 0.2145703, 0.2536921, 0.3344125, 
    0.2883532, 0.403367, 0.2760895, 0.2979332, 0.2418465, 0.09240174, 
    0.2670472, 0.2529185, 0.3369473, 0.2651588, 0.1641679, 0.2048902, 
    0.2723401, 0.2310941, 0.1901069, 0.1909665, 0.2001357, 0.3934716, 
    0.1650099, 0.2226174, 0.1896408, 0.2559896, 0.2833514,
  0.2803185, 0.3310972, 0.3229807, 0.3033306, 0.3409346, 0.3094964, 
    0.4151571, 0.4323036, 0.2845327, 0.1943538, 0.2475557, 0.199081, 
    0.3538458, 0.3180867, 0.3147137, 0.2863183, 0.2940269, 0.3465273, 
    0.3572291, 0.2863353, 0.2316304, 0.2017998, 0.1624775, 0.08042807, 
    0.2943622, 0.1657966, 0.1904754, 0.170746, 0.2989002,
  0.2945877, 0.3326252, 0.157823, 0.07934036, 0.05869424, 0.1157866, 
    0.1107841, 0.1023338, 0.1358296, 0.2164278, 0.2332894, 0.2507815, 
    0.1914818, 0.2433082, 0.2456095, 0.172266, 0.1661079, 0.2207674, 
    0.2723745, 0.2279045, 0.1924064, 0.2559513, 0.2394075, 0.07907064, 
    0.09672354, 0.04226491, 0.0264572, 0.109664, 0.2359347,
  0.2133387, 0.2105108, 0.207683, 0.2048551, 0.2020272, 0.1991993, 0.1963714, 
    0.2085183, 0.2091304, 0.2097424, 0.2103545, 0.2109666, 0.2115787, 
    0.2121907, 0.2076249, 0.2130489, 0.218473, 0.223897, 0.229321, 0.2347451, 
    0.2401691, 0.2336432, 0.230435, 0.2272267, 0.2240185, 0.2208103, 
    0.2176021, 0.2143939, 0.2156011,
  0.1348311, 0.1685959, 0.1224102, 0.04365751, 0.04323765, 0.008027693, 
    0.00358344, 0.0192174, 0.05997057, 0.1228514, 0.153238, 0.1799322, 
    0.2259888, 0.1449054, 0.05568902, 0.1402302, 0.159436, 0.2020425, 
    0.1942937, 0.1991351, 0.2031334, 0.3589931, 0.2529955, 0.1027902, 
    0.1326143, 0.2360052, 0.2433555, 0.1607205, 0.1104364,
  0.1071903, 0.2396239, 0.2582904, 0.4233003, 0.4169235, 0.2884804, 
    0.2135947, 0.2578904, 0.2278458, 0.2181733, 0.1702, 0.165601, 0.2244858, 
    0.2011912, 0.1993726, 0.2001668, 0.26962, 0.2468587, 0.2087732, 
    0.1763144, 0.2453974, 0.2813577, 0.3404925, 0.3597964, 0.2325307, 
    0.1912191, 0.1938732, 0.09867613, 0.02555415,
  0.1634079, 0.2360813, 0.3489994, 0.3351899, 0.2906868, 0.2861712, 
    0.2736046, 0.2209679, 0.2317372, 0.2479533, 0.276315, 0.2838134, 
    0.2603631, 0.2093163, 0.2093578, 0.2093039, 0.2091311, 0.2264294, 
    0.2792363, 0.2749096, 0.3002985, 0.2689113, 0.2964867, 0.2320416, 
    0.2678463, 0.292457, 0.2470218, 0.2215486, 0.2768998,
  0.2112884, 0.1981253, 0.1538085, 0.1908664, 0.1446351, 0.1403435, 
    0.1426505, 0.1796662, 0.2019336, 0.1908767, 0.1558759, 0.1549945, 
    0.1700784, 0.1785763, 0.1391596, 0.1099871, 0.09370661, 0.1063733, 
    0.1358214, 0.1114018, 0.1834134, 0.1525611, 0.1431892, 0.1144612, 
    0.1615896, 0.1255951, 0.140503, 0.1417485, 0.1902049,
  0.04477798, 0.02701457, 0.02949385, 0.08920028, 0.1192446, 0.04812978, 
    0.06831655, 0.0630201, 0.05629072, 0.03931816, 0.0754914, 0.06297188, 
    0.06320595, 0.04235438, 0.1009754, 0.1475354, 0.1211836, 0.01563026, 
    0.06090402, 0.1213128, 0.08774205, 0.1079044, 0.05037886, 0.008742182, 
    0.08799947, 0.1267221, 0.1426317, 0.1102394, 0.07062855,
  0.004075658, -2.906794e-07, 0.1264748, 0.06159246, 0.1115723, 0.07331952, 
    0.06948709, 0.003729362, 1.482772e-05, 0.0005778054, 0.02536526, 
    0.044324, 0.09729177, 0.00529705, 0.05745655, 0.007613251, 0.02740356, 
    0.1682124, 0.1437594, 0.04372475, 0.02796886, 0.002330561, 1.06014e-05, 
    2.177406e-05, 0.05778833, 0.08195668, 0.1009065, 0.00335985, 0.006627866,
  9.947196e-05, 0.04296298, 0.1568534, 0.03109969, 0.02250556, 0.01042631, 
    0.09149279, 1.186354e-06, 6.72228e-07, 0.002768778, 0.06356122, 
    0.07978622, 0.01080122, 0.04378127, 0.04608046, 0.120428, 0.04597892, 
    0.1512391, 0.02275237, 0.01208112, 0.0004807018, 6.107317e-09, 
    1.114099e-05, 0.0003871317, 0.1027061, 0.2152104, 0.007842021, 
    8.033499e-06, 2.508725e-07,
  0.01848259, 0.1115586, 0.1699653, 0.1067047, 0.08165928, 0.03826153, 
    0.1214086, 0.1384071, 0.01004416, 0.0303643, 0.0499615, 0.03348581, 
    0.03565626, 0.09958652, 0.07579861, 0.04015327, 0.02059802, 0.01314578, 
    0.005254738, 0.0009772306, 1.767411e-07, 1.182354e-07, 0.004203379, 
    0.1479962, 0.3280747, 0.1338989, 0.008100706, 7.400409e-06, 0.001337582,
  0.418967, 0.09410097, 0.1057061, 0.03672466, 0.04993371, 0.0336678, 
    0.1044789, 0.03773754, 0.1420321, 0.2508874, 0.04943542, 0.01076884, 
    0.04604383, 0.06819292, 0.01761303, 0.005502322, 0.00109598, 
    -5.565384e-05, 4.586032e-05, -9.399432e-05, 0.0165729, 0.03077128, 
    0.2349626, 0.2082801, 0.1041832, 0.07958963, 0.04062589, 0.02530148, 
    0.06043095,
  -1.028714e-05, 2.738403e-06, 0.01337506, 0.0243102, 0.03366876, 0.0124972, 
    0.0003570023, 0.002229402, 0.08909488, 0.0486416, 0.04586881, 0.05719448, 
    0.04755486, 0.07115165, 0.06194288, 0.05162055, 0.08957785, 0.05535807, 
    0.09890748, 0.1018512, 0.06671283, 0.01091973, 0.01175709, 0.02014299, 
    0.06866506, 0.01766413, 0.01825812, 0.004995991, 0.0004227472,
  0.0008334047, 1.793951e-06, 9.701439e-07, 2.679922e-05, 0.02651178, 
    0.007917689, 0.0004668216, 9.43079e-07, 1.723749e-05, 0.07793402, 
    0.0926433, 0.03836627, 6.498126e-05, 0.001558891, 0.002882671, 
    0.007309697, 0.05844878, 0.1088348, 0.03446466, 0.0008183604, 0.02881676, 
    0.01768234, 0.005636503, 0.01076884, 0.05707769, 0.01500998, 
    0.0008978946, 1.415611e-05, 0.03514871,
  0.0002758316, 0.01098892, 0.01310986, 0.03891364, 0.06152747, 0.1449656, 
    0.07129582, 0.08561929, 0.1797399, 0.1983426, 0.1260493, 0.09149811, 
    0.09539688, 0.09093551, 0.05922535, 0.1280988, 0.109122, 0.1108448, 
    0.092965, 0.04468438, 0.1118041, 0.06875733, 0.02650387, 0.01139498, 
    0.05322669, 0.08198514, 0.01849361, 0.009202858, 0.03935325,
  0.0531822, 0.04536282, 0.1658371, 0.1759989, 0.1529964, 0.0968194, 
    0.1447306, 0.08074448, 0.04735369, 0.1147079, 0.04905719, 0.09057718, 
    0.07995953, 0.1765904, 0.190467, 0.1420831, 0.135591, 0.06870504, 
    0.09458768, 0.1673479, 0.1771989, 0.08957943, 0.1841441, 0.1657731, 
    0.1830853, 0.1589865, 0.1332622, 0.07091115, 0.1368065,
  0.1823905, 0.1363487, 0.1013225, 0.1799296, 0.1646183, 0.1461866, 
    0.1924406, 0.1762788, 0.1802209, 0.08699152, 0.06176047, 0.05601876, 
    0.2464704, 0.1839686, 0.258857, 0.2370376, 0.08092103, 0.06257087, 
    0.129549, 0.3219072, 0.1341612, 0.1452992, 0.2096083, 0.2509708, 
    0.1699386, 0.1736895, 0.2434413, 0.2211815, 0.2042943,
  0.296379, 0.2958961, 0.2407453, 0.2047321, 0.2627639, 0.3411379, 0.3032918, 
    0.4185621, 0.3015596, 0.3235247, 0.3130132, 0.09509153, 0.320648, 
    0.2553071, 0.336232, 0.2649518, 0.185211, 0.2104256, 0.2760354, 
    0.2821446, 0.2048246, 0.2227836, 0.1662816, 0.3741437, 0.205438, 
    0.2305997, 0.1975012, 0.2712633, 0.30445,
  0.3121304, 0.3147791, 0.349377, 0.2893282, 0.3375816, 0.3388442, 0.4267591, 
    0.4359991, 0.2999941, 0.2487181, 0.2514626, 0.2608978, 0.3631947, 
    0.3281666, 0.3527422, 0.2743041, 0.2859853, 0.354234, 0.3894939, 
    0.3285774, 0.2882544, 0.2415071, 0.2056371, 0.1307121, 0.271429, 
    0.2611225, 0.315897, 0.2055969, 0.3014203,
  0.3212165, 0.3356033, 0.1439908, 0.07623159, 0.07600901, 0.1386486, 
    0.1172149, 0.1415816, 0.1324802, 0.2416528, 0.187413, 0.2353968, 
    0.1826437, 0.2381374, 0.2471875, 0.1759197, 0.1727629, 0.237445, 
    0.2884507, 0.245322, 0.2287736, 0.304717, 0.2792512, 0.08402103, 
    0.1010601, 0.04836548, 0.04932566, 0.1730944, 0.2861776,
  0.2245434, 0.2263062, 0.2280689, 0.2298317, 0.2315944, 0.2333572, 
    0.2351199, 0.2520762, 0.2548577, 0.2576393, 0.2604208, 0.2632023, 
    0.2659838, 0.2687654, 0.2815106, 0.2864562, 0.2914018, 0.2963474, 
    0.301293, 0.3062386, 0.3111842, 0.282798, 0.2733082, 0.2638183, 
    0.2543284, 0.2448385, 0.2353486, 0.2258587, 0.2231332,
  0.1282396, 0.1872784, 0.1950679, 0.1326868, 0.0889495, 0.05585773, 
    0.01719507, 0.03268135, 0.1320803, 0.2117315, 0.1996794, 0.2383634, 
    0.2741697, 0.1488848, 0.1129334, 0.1068407, 0.1573456, 0.2029873, 
    0.186432, 0.1911826, 0.1959793, 0.3702277, 0.2482489, 0.1060924, 
    0.1214486, 0.2062632, 0.2391036, 0.1612981, 0.1269298,
  0.1279431, 0.2734445, 0.2998877, 0.4520567, 0.4434319, 0.2901924, 
    0.2044593, 0.2854053, 0.2429363, 0.2232576, 0.167819, 0.1633235, 
    0.2406256, 0.221942, 0.265522, 0.2458835, 0.3304362, 0.3134539, 
    0.2603908, 0.2999281, 0.2229574, 0.3284139, 0.4012936, 0.4037164, 
    0.2108329, 0.1779055, 0.1736785, 0.2199146, 0.05998966,
  0.2813805, 0.3182682, 0.4004187, 0.3367898, 0.3274438, 0.2593967, 
    0.2551661, 0.2495003, 0.2618424, 0.2501472, 0.3397336, 0.3223642, 
    0.3070431, 0.2187815, 0.1983339, 0.2211563, 0.2116918, 0.2188969, 
    0.2733395, 0.2688975, 0.300104, 0.2603438, 0.2835295, 0.1876911, 
    0.3002444, 0.3252612, 0.29099, 0.2498063, 0.3241685,
  0.2095966, 0.1926752, 0.1415133, 0.2030961, 0.1363338, 0.1443827, 
    0.1478214, 0.1849468, 0.2223768, 0.2084645, 0.1579061, 0.1410833, 
    0.1712036, 0.1682903, 0.1266927, 0.1094093, 0.09053168, 0.122427, 
    0.1314781, 0.1152677, 0.1854987, 0.1430335, 0.1259428, 0.1211873, 
    0.1469808, 0.1153631, 0.1428316, 0.1163949, 0.1649826,
  0.05713147, 0.03021304, 0.02998499, 0.0720538, 0.1242748, 0.05093426, 
    0.07279754, 0.06378971, 0.07906043, 0.03860611, 0.0591356, 0.06427716, 
    0.05165564, 0.05796049, 0.1160674, 0.1552795, 0.1151376, 0.01681998, 
    0.06767634, 0.1337387, 0.1075504, 0.1199351, 0.06425346, 0.008717353, 
    0.07662009, 0.1282963, 0.137391, 0.1249353, 0.06540246,
  0.006918339, -4.797348e-08, 0.1310437, 0.06741943, 0.1021458, 0.07312521, 
    0.06549792, 0.00242687, 3.739237e-06, 6.675008e-05, 0.008027675, 
    0.02454943, 0.09330592, 0.006467952, 0.07663627, 0.008670243, 0.02357135, 
    0.1710244, 0.1240929, 0.03807693, 0.04630854, 0.004348724, 1.359754e-05, 
    2.235308e-05, 0.03820163, 0.08392978, 0.08895186, 0.004892848, 0.008825754,
  7.408604e-06, 0.02008198, 0.1563164, 0.02687426, 0.02731525, 0.009816788, 
    0.08450417, 4.80914e-06, 1.353528e-06, 0.001906238, 0.05687405, 
    0.04737418, 0.01857267, 0.05293558, 0.04986399, 0.07788335, 0.0446107, 
    0.09914953, 0.02572584, 0.02107441, 0.006127011, 1.601356e-08, 
    7.269652e-06, 0.0002073845, 0.1003169, 0.2397635, 0.01054993, 
    4.552959e-06, 1.535209e-07,
  0.006046288, 0.04620581, 0.1978368, 0.0841087, 0.08627594, 0.03450796, 
    0.1085421, 0.1224264, 0.009912034, 0.02260796, 0.04323162, 0.02586851, 
    0.03448965, 0.08780538, 0.06083757, 0.0410276, 0.02150373, 0.0189582, 
    0.009344826, 0.0004521372, -2.833705e-07, -1.267902e-06, 0.002061097, 
    0.09928057, 0.2256595, 0.1172766, 0.009500532, 2.310686e-06, 0.0004575749,
  0.3823668, 0.08574432, 0.1031137, 0.05123971, 0.05321707, 0.02946959, 
    0.09749974, 0.02997659, 0.1252774, 0.1960455, 0.04705567, 0.01062046, 
    0.0299405, 0.06217985, 0.01402027, 0.003628331, 0.009955543, 
    -2.449904e-05, 0.0001466447, 7.619389e-06, 0.01249769, 0.02161124, 
    0.2032787, 0.192523, 0.1072095, 0.06210996, 0.04341993, 0.01817869, 
    0.04027889,
  4.526552e-06, 1.680231e-06, 0.003407505, 0.09515464, 0.03900961, 
    0.008056276, 0.002030232, 0.004792673, 0.08261003, 0.04200256, 
    0.04848947, 0.05101521, 0.04518092, 0.07170296, 0.05763778, 0.03566213, 
    0.07935771, 0.06878299, 0.1029598, 0.1055379, 0.06363314, 0.01459291, 
    0.03311608, 0.02500945, 0.06945643, 0.01642652, 0.006351535, 
    0.0006841589, 0.0007520278,
  7.499359e-05, 7.463546e-07, 8.703276e-07, 0.0001240332, 0.02661835, 
    0.0001810373, 0.001189039, -1.856553e-06, 2.581278e-06, 0.04879707, 
    0.1167953, 0.04036593, 5.495668e-05, 0.002753181, 0.005724495, 
    0.01008321, 0.05165959, 0.1378216, 0.03260023, 0.0006525647, 0.01475162, 
    0.01696226, 0.01472537, 0.0240257, 0.06489715, 0.0170692, 0.0006867744, 
    0.001862781, 0.01284549,
  9.409363e-05, 0.005060607, 0.0102538, 0.03929314, 0.08116195, 0.1462454, 
    0.06497414, 0.08580122, 0.2006339, 0.2102272, 0.1231854, 0.08632664, 
    0.09069739, 0.09619657, 0.06109133, 0.1501247, 0.1175885, 0.1195392, 
    0.1068475, 0.05285297, 0.1451449, 0.07963277, 0.02306388, 0.005113926, 
    0.0615389, 0.08816856, 0.02591571, 0.01403487, 0.03459187,
  0.0508752, 0.05321816, 0.156769, 0.2105737, 0.1692025, 0.09603305, 
    0.1638746, 0.06251016, 0.04667728, 0.1055879, 0.05518059, 0.08262819, 
    0.08527616, 0.1785926, 0.1927808, 0.1505234, 0.1465411, 0.08132491, 
    0.09996168, 0.2016945, 0.193739, 0.0930851, 0.1785689, 0.1663653, 
    0.1905547, 0.1771191, 0.1423448, 0.09155658, 0.1474712,
  0.1788554, 0.1362617, 0.1001635, 0.1639712, 0.1584038, 0.1642659, 
    0.2072344, 0.1791389, 0.1665275, 0.07362603, 0.06633864, 0.05059224, 
    0.2609121, 0.2192866, 0.2527429, 0.2334669, 0.08130776, 0.05582757, 
    0.1280971, 0.3327733, 0.1605935, 0.1298211, 0.2221864, 0.2901326, 
    0.1526112, 0.1859529, 0.2714055, 0.2091207, 0.2050648,
  0.2914166, 0.286086, 0.2432008, 0.2526807, 0.3336744, 0.4023907, 0.316947, 
    0.4201756, 0.2697179, 0.328276, 0.340928, 0.09249809, 0.3303452, 
    0.2810676, 0.339543, 0.2910875, 0.1939274, 0.2198134, 0.2602583, 
    0.2920166, 0.229671, 0.2080079, 0.2369877, 0.4131069, 0.2193954, 
    0.2282165, 0.2231707, 0.2952866, 0.307279,
  0.333055, 0.3547881, 0.3736758, 0.3693262, 0.3532301, 0.4696627, 0.5619112, 
    0.4753084, 0.3147826, 0.239639, 0.3053684, 0.2534806, 0.3999265, 
    0.3401216, 0.3597668, 0.288389, 0.2888923, 0.3572621, 0.4092575, 
    0.3880441, 0.3155158, 0.2050081, 0.2457876, 0.1599234, 0.2502836, 
    0.3217756, 0.4041639, 0.3525793, 0.3228376,
  0.4043815, 0.3413097, 0.1814714, 0.09072074, 0.07462935, 0.1612915, 
    0.1701266, 0.2155869, 0.1594545, 0.2737891, 0.2024621, 0.2630633, 
    0.2415155, 0.2512451, 0.25803, 0.1961711, 0.1710654, 0.238859, 0.3018489, 
    0.2777458, 0.2269952, 0.3142766, 0.2876682, 0.1027848, 0.07762937, 
    0.07715271, 0.09470129, 0.1964527, 0.3867711,
  0.2106881, 0.2120548, 0.2134215, 0.2147882, 0.2161549, 0.2175216, 
    0.2188883, 0.2248279, 0.2327773, 0.2407265, 0.2486759, 0.2566251, 
    0.2645744, 0.2725238, 0.2800113, 0.2814701, 0.2829289, 0.2843877, 
    0.2858466, 0.2873054, 0.2887642, 0.2703517, 0.2595769, 0.2488021, 
    0.2380272, 0.2272524, 0.2164776, 0.2057028, 0.2095948,
  0.1223254, 0.180681, 0.2149562, 0.1759423, 0.1175277, 0.1130017, 
    0.05060038, 0.1187935, 0.1939757, 0.223161, 0.2202625, 0.2470463, 
    0.2615833, 0.1479137, 0.05981699, 0.04034652, 0.1357329, 0.2032031, 
    0.174655, 0.2357364, 0.2053151, 0.3625994, 0.2476939, 0.1059303, 
    0.1486961, 0.2899455, 0.2655443, 0.1733563, 0.127941,
  0.1498908, 0.3553434, 0.3222931, 0.4528313, 0.4446029, 0.3007318, 
    0.1987745, 0.2756217, 0.2562005, 0.247896, 0.1636284, 0.1761859, 
    0.259116, 0.228305, 0.2548269, 0.2680975, 0.3928919, 0.3020729, 
    0.2207872, 0.3050613, 0.3565164, 0.3850766, 0.3994961, 0.4230168, 
    0.2153231, 0.1641548, 0.1973943, 0.1955495, 0.1145922,
  0.38979, 0.4915627, 0.4865275, 0.4041512, 0.3676815, 0.3420614, 0.3224455, 
    0.2536795, 0.3131947, 0.3104669, 0.3288614, 0.2873532, 0.3259121, 
    0.2349999, 0.2195984, 0.2157657, 0.2144336, 0.2224668, 0.2745863, 
    0.2875004, 0.3333421, 0.2576394, 0.2978662, 0.2116856, 0.2699849, 
    0.265911, 0.2503772, 0.2628285, 0.3790919,
  0.2542723, 0.1942834, 0.1437166, 0.2088224, 0.1320832, 0.142538, 0.1638485, 
    0.1841247, 0.2167185, 0.2334573, 0.1836659, 0.1718587, 0.1779684, 
    0.1741638, 0.1327062, 0.1053183, 0.09049726, 0.1359938, 0.1505835, 
    0.1326551, 0.1936402, 0.1597214, 0.1451679, 0.1475223, 0.1398712, 
    0.1171266, 0.1484689, 0.1403792, 0.1889432,
  0.06273812, 0.03708386, 0.03523028, 0.07418704, 0.1415223, 0.06400598, 
    0.08966348, 0.06558599, 0.08262773, 0.04151122, 0.04511783, 0.06398465, 
    0.04409182, 0.04265516, 0.1318576, 0.1664331, 0.1214432, 0.0307174, 
    0.07430855, 0.1460957, 0.1090273, 0.1435126, 0.08928055, 0.01189122, 
    0.06343805, 0.1264823, 0.1433928, 0.1324681, 0.0712563,
  0.02062617, 9.5738e-10, 0.1268194, 0.05755826, 0.05858101, 0.07763581, 
    0.05681703, 0.01114975, 3.308099e-06, 3.160933e-06, 0.0007743063, 
    0.01817174, 0.05305071, 0.00612672, 0.08435237, 0.02193854, 0.0244002, 
    0.1703761, 0.1016913, 0.03593218, 0.05304697, 0.009349448, 1.038845e-05, 
    1.245431e-05, 0.02612341, 0.0678833, 0.07143337, 0.00624011, 0.01274534,
  1.16524e-06, 0.0094953, 0.1191252, 0.02449686, 0.03619161, 0.01398975, 
    0.08543679, 4.827466e-06, 2.962394e-07, 6.19668e-05, 0.05089154, 
    0.04141817, 0.03459682, 0.05180398, 0.05489876, 0.06529091, 0.04125743, 
    0.06197964, 0.03710794, 0.03899971, 0.02083801, -3.264112e-07, 
    4.919872e-06, 4.667463e-05, 0.1015133, 0.2272811, 0.01638019, 
    0.0008671114, 1.661294e-07,
  0.0008056894, 0.0203923, 0.169433, 0.08110634, 0.08114487, 0.03303606, 
    0.1079034, 0.1189396, 0.01089754, 0.01667136, 0.03850866, 0.01981914, 
    0.03212802, 0.08407038, 0.0558644, 0.04195859, 0.02791373, 0.03098193, 
    0.02322264, 0.001227126, 1.617262e-06, 1.306207e-07, 0.001135001, 
    0.09487981, 0.1871779, 0.0939054, 0.01156481, 2.195792e-06, 7.571422e-06,
  0.3275318, 0.05684722, 0.09803123, 0.06869332, 0.05755147, 0.03586861, 
    0.09270856, 0.02633501, 0.1291177, 0.1713458, 0.04243658, 0.009039353, 
    0.02846905, 0.0534234, 0.01506706, 0.004105689, 0.005587059, 
    -0.0004058517, 0.000803167, 0.0002190134, 0.008936057, 0.01881512, 
    0.1657536, 0.1995386, 0.1097244, 0.04733797, 0.04412803, 0.01934451, 
    0.03093567,
  9.506462e-07, 5.872769e-07, 0.001879958, 0.1654508, 0.04836267, 
    0.008629548, 0.002625356, 0.005111658, 0.08581887, 0.04425715, 
    0.05878477, 0.05052878, 0.04627771, 0.07312143, 0.07062281, 0.02505344, 
    0.06498932, 0.08398157, 0.1095544, 0.1025627, 0.06101236, 0.01855345, 
    0.04602349, 0.03074088, 0.07423539, 0.01906788, 0.00188373, 3.158427e-05, 
    0.0006738799,
  8.953779e-05, 6.690896e-07, 4.166819e-07, 0.000146881, 0.02851119, 
    0.00319133, 0.001145745, -1.857346e-06, 9.783664e-05, 0.05023679, 
    0.119293, 0.04298032, 0.00117506, 0.003997155, 0.01203883, 0.01236177, 
    0.04682093, 0.1634989, 0.03398917, 0.001836804, 0.01645089, 0.03671601, 
    0.024673, 0.04620746, 0.06543032, 0.02950128, 0.008563883, 0.007510012, 
    0.000614245,
  8.195278e-06, 0.003754268, 0.01463613, 0.04207315, 0.09650981, 0.152206, 
    0.0801857, 0.07573079, 0.2039227, 0.2018116, 0.1202911, 0.07960582, 
    0.08196911, 0.09286876, 0.07435078, 0.1687279, 0.1332885, 0.1265999, 
    0.1315871, 0.07393351, 0.1735907, 0.07292796, 0.01580123, 0.006302074, 
    0.06164631, 0.08046185, 0.02749768, 0.0258293, 0.03611212,
  0.06629161, 0.07555501, 0.1667937, 0.2824208, 0.1919836, 0.05383854, 
    0.1682019, 0.0499981, 0.04484176, 0.10464, 0.06709076, 0.09939142, 
    0.1175144, 0.1889086, 0.1869157, 0.1589688, 0.1555345, 0.1144765, 
    0.103408, 0.2335903, 0.2019919, 0.0858176, 0.1681419, 0.1732426, 
    0.211797, 0.2087807, 0.1660968, 0.1241324, 0.1598744,
  0.1839659, 0.1282796, 0.08541704, 0.1778197, 0.1757602, 0.1922905, 
    0.215527, 0.1714761, 0.1642101, 0.06962258, 0.06720903, 0.04642696, 
    0.2823302, 0.2166469, 0.256019, 0.2314541, 0.09969729, 0.06603803, 
    0.1357097, 0.3488183, 0.1774279, 0.1248742, 0.2242697, 0.2852941, 
    0.1452972, 0.1774852, 0.2831694, 0.2237766, 0.2218021,
  0.2711633, 0.3142421, 0.2344636, 0.2269529, 0.3792288, 0.4697331, 
    0.4002311, 0.4185114, 0.2878883, 0.3351571, 0.3834419, 0.1102508, 
    0.3521846, 0.2627237, 0.322173, 0.3012994, 0.2023091, 0.2314741, 
    0.2495791, 0.3284277, 0.2269368, 0.1951531, 0.272729, 0.4016697, 
    0.195874, 0.2302427, 0.2502499, 0.2976174, 0.304421,
  0.339557, 0.3164373, 0.4585217, 0.4168463, 0.3758239, 0.4669311, 0.5794992, 
    0.5144405, 0.282015, 0.240429, 0.3096192, 0.2752824, 0.4232775, 
    0.3521792, 0.3678695, 0.2662159, 0.2758796, 0.3853752, 0.3803184, 
    0.4049235, 0.3495738, 0.219584, 0.2863573, 0.1776777, 0.2366772, 
    0.3609447, 0.4302319, 0.4240524, 0.3368098,
  0.3254744, 0.3249723, 0.1778055, 0.1082189, 0.1143169, 0.1740976, 
    0.1579678, 0.2278438, 0.1574243, 0.236988, 0.2544665, 0.3171678, 
    0.3201482, 0.2810957, 0.2824462, 0.2151289, 0.1960468, 0.256184, 
    0.3648123, 0.3191742, 0.2537623, 0.2972151, 0.2918577, 0.1244939, 
    0.06600873, 0.08974443, 0.1118697, 0.2147436, 0.4016651,
  0.1849882, 0.1856724, 0.1863566, 0.1870407, 0.1877249, 0.188409, 0.1890932, 
    0.2118551, 0.221373, 0.230891, 0.2404089, 0.2499268, 0.2594447, 
    0.2689627, 0.2666764, 0.2668773, 0.2670783, 0.2672793, 0.2674803, 
    0.2676812, 0.2678822, 0.2420392, 0.2316362, 0.2212331, 0.2108301, 
    0.200427, 0.190024, 0.1796209, 0.1844409,
  0.1176915, 0.1657309, 0.2352078, 0.1929036, 0.168942, 0.1331067, 0.1110287, 
    0.1894689, 0.2104648, 0.1965354, 0.2113777, 0.2357565, 0.245425, 
    0.09404441, 0.04210798, 0.105726, 0.09971575, 0.1901118, 0.1792948, 
    0.2177207, 0.2129613, 0.3957721, 0.2891699, 0.1216379, 0.1660108, 
    0.2770659, 0.2334404, 0.1705147, 0.1160617,
  0.1415627, 0.2380612, 0.3100672, 0.4333051, 0.4328553, 0.2989261, 
    0.1758934, 0.2668678, 0.2419039, 0.2565748, 0.1754287, 0.1668743, 
    0.2426037, 0.1878195, 0.2632368, 0.2614962, 0.3130581, 0.3128948, 
    0.3224578, 0.2657825, 0.2364445, 0.3295549, 0.4492245, 0.4296551, 
    0.1740928, 0.1428997, 0.1802594, 0.1894424, 0.1280581,
  0.2378608, 0.3725888, 0.3943331, 0.4328159, 0.3169603, 0.3195345, 
    0.2913388, 0.3164366, 0.2835828, 0.2833959, 0.3295871, 0.302838, 
    0.3292026, 0.2813852, 0.2161377, 0.2245733, 0.2215537, 0.2776283, 
    0.2984998, 0.2822604, 0.3043565, 0.2837571, 0.2890811, 0.2263767, 
    0.2886311, 0.2449501, 0.2249007, 0.2462843, 0.2832173,
  0.2566663, 0.2183609, 0.1705996, 0.2077952, 0.1424645, 0.1552967, 
    0.1715189, 0.2069667, 0.2546018, 0.2687005, 0.20711, 0.1943079, 
    0.2062731, 0.174674, 0.1361857, 0.1164969, 0.1173445, 0.1461469, 
    0.1638546, 0.1393082, 0.2161001, 0.1852054, 0.1699731, 0.1595219, 
    0.1212699, 0.1005091, 0.1456913, 0.1363168, 0.1960393,
  0.07542076, 0.046546, 0.04575924, 0.08229671, 0.1109149, 0.07751531, 
    0.09229179, 0.07023491, 0.08900241, 0.04979347, 0.05281589, 0.06418507, 
    0.04285906, 0.03448853, 0.1443718, 0.1562485, 0.1363448, 0.0260823, 
    0.07502161, 0.1273802, 0.1094429, 0.1690461, 0.09216935, 0.01478592, 
    0.06153534, 0.1270526, 0.1424489, 0.1303499, 0.08177148,
  0.0278824, 2.236717e-08, 0.1096264, 0.06814013, 0.02722469, 0.0801243, 
    0.05488944, 0.01110473, 2.541576e-06, 6.156227e-07, 0.0001712321, 
    0.01354416, 0.03061357, 0.0121114, 0.08636548, 0.0548908, 0.03729724, 
    0.1782969, 0.08186138, 0.03183581, 0.06285168, 0.01129783, 0.0001269219, 
    6.461883e-06, 0.02299698, 0.07170396, 0.07356816, 0.02092825, 0.01627932,
  7.802406e-07, 0.003212928, 0.1024067, 0.02090117, 0.04127311, 0.01731626, 
    0.08482084, 0.002412186, -5.549133e-08, 1.410942e-06, 0.03757602, 
    0.02700607, 0.05592633, 0.04674989, 0.05781546, 0.06317342, 0.03642715, 
    0.04560654, 0.03505997, 0.05365742, 0.03915971, 0.000496732, 
    1.496383e-06, 2.572119e-05, 0.09933326, 0.2110703, 0.02333601, 
    0.009491332, 2.521483e-06,
  1.356196e-05, 0.01075, 0.1668189, 0.07791346, 0.07491165, 0.03549328, 
    0.1011305, 0.1106256, 0.01345241, 0.01434292, 0.03956053, 0.01662926, 
    0.03481129, 0.07763429, 0.04950917, 0.04008655, 0.03391364, 0.03362398, 
    0.02910603, 0.0033646, 1.529729e-08, 8.790727e-08, 3.712676e-05, 
    0.1013209, 0.1649817, 0.08008872, 0.01778676, 6.067476e-06, 3.395058e-06,
  0.2910362, 0.03759564, 0.09388086, 0.08862605, 0.05601262, 0.0357716, 
    0.08808489, 0.02791945, 0.1387334, 0.169085, 0.03820473, 0.008730464, 
    0.02853916, 0.0459233, 0.01674638, 0.005750247, 0.002434873, 
    0.0006189077, 0.001463351, 0.0002438345, 0.001401155, 0.01253975, 
    0.1340676, 0.1856244, 0.1213639, 0.03795126, 0.04531685, 0.02918954, 
    0.03084435,
  3.185733e-07, 1.51868e-07, -8.433872e-05, 0.1593198, 0.0597102, 0.01667973, 
    0.005877868, 0.008116751, 0.09448574, 0.04298981, 0.07219664, 0.05685055, 
    0.05545983, 0.08661683, 0.09206942, 0.03077446, 0.06153004, 0.09689464, 
    0.1198315, 0.1047221, 0.05736125, 0.02391822, 0.05022291, 0.03532759, 
    0.07024332, 0.02169563, 0.0009623105, 0.000112659, 4.313615e-05,
  7.808914e-06, 7.175313e-07, 1.09652e-07, 0.002750237, 0.01689654, 
    0.01030443, 0.002657976, -7.034399e-06, 0.00936715, 0.07705427, 0.115026, 
    0.05646589, 0.01755347, 0.008894453, 0.0162436, 0.01923962, 0.04126568, 
    0.1475057, 0.03457957, 0.005771207, 0.02173644, 0.06778795, 0.02704284, 
    0.04740328, 0.05870929, 0.0695717, 0.05780347, 0.006636519, 6.505757e-06,
  1.255604e-06, 0.01426931, 0.02966882, 0.05493395, 0.1034923, 0.1590662, 
    0.04720616, 0.05293657, 0.1795349, 0.1909611, 0.1196178, 0.0716588, 
    0.08440901, 0.1014718, 0.0767144, 0.182725, 0.1531271, 0.1289749, 
    0.1499798, 0.07885276, 0.1685866, 0.06348291, 0.01970156, 0.01041822, 
    0.06546265, 0.0794747, 0.03955191, 0.03254007, 0.05574545,
  0.05621494, 0.09960991, 0.1994055, 0.3092544, 0.1886313, 0.05904908, 
    0.1824824, 0.04311473, 0.04226021, 0.08528041, 0.06299347, 0.1266471, 
    0.1627113, 0.1946077, 0.2034303, 0.1908348, 0.1852198, 0.1220423, 
    0.1191305, 0.2397785, 0.2208091, 0.07781491, 0.173897, 0.1801988, 
    0.2361059, 0.2177862, 0.1832718, 0.1400497, 0.1779592,
  0.1773952, 0.1340231, 0.08605464, 0.1763674, 0.167483, 0.1921189, 0.179666, 
    0.1589258, 0.1652885, 0.07527865, 0.06618325, 0.03973012, 0.3245666, 
    0.2351403, 0.3021185, 0.2240085, 0.1580281, 0.07860775, 0.1502105, 
    0.3445769, 0.1384434, 0.1247292, 0.195706, 0.2445634, 0.1500746, 
    0.2150103, 0.2903005, 0.2431524, 0.2100616,
  0.2460382, 0.2731104, 0.246159, 0.264661, 0.3780629, 0.4477364, 0.3812849, 
    0.4819314, 0.2879519, 0.369636, 0.4181185, 0.133662, 0.4020995, 
    0.2746076, 0.3051574, 0.2763285, 0.2197158, 0.2373599, 0.2463288, 
    0.3069659, 0.2555893, 0.2105949, 0.2063279, 0.3608328, 0.2109015, 
    0.2323716, 0.2461858, 0.301481, 0.2962962,
  0.3635351, 0.3162385, 0.3618099, 0.3668675, 0.4073585, 0.476043, 0.5172926, 
    0.5359262, 0.2666412, 0.2628241, 0.2931131, 0.2711233, 0.4380771, 
    0.3548208, 0.3401217, 0.2248709, 0.2869072, 0.404884, 0.3601041, 
    0.4037149, 0.3443903, 0.1934225, 0.3030692, 0.1701723, 0.1866914, 
    0.3980065, 0.4582863, 0.3962487, 0.3250492,
  0.3454848, 0.4521009, 0.2624436, 0.1141067, 0.0693688, 0.1504282, 
    0.1250257, 0.1236525, 0.1189331, 0.2106086, 0.261777, 0.2625242, 
    0.2992034, 0.2949787, 0.2659715, 0.2464713, 0.2193299, 0.2692763, 
    0.358648, 0.2989082, 0.2547392, 0.2995592, 0.2766418, 0.1356692, 
    0.05680995, 0.06829368, 0.1270092, 0.2612748, 0.4473844,
  0.1654041, 0.1652822, 0.1651603, 0.1650384, 0.1649165, 0.1647945, 
    0.1646726, 0.2009898, 0.2110285, 0.2210672, 0.231106, 0.2411447, 
    0.2511834, 0.2612221, 0.2497094, 0.2508593, 0.2520091, 0.253159, 
    0.2543088, 0.2554587, 0.2566085, 0.2588316, 0.2477649, 0.2366982, 
    0.2256315, 0.2145649, 0.2034982, 0.1924316, 0.1655017,
  0.1161799, 0.1485025, 0.2305062, 0.2190278, 0.1852999, 0.1535667, 
    0.1539229, 0.2521155, 0.2424963, 0.1942248, 0.2080633, 0.2190441, 
    0.2719715, 0.06321286, 0.06274096, 0.06611771, 0.1309869, 0.1716229, 
    0.1361026, 0.2095218, 0.2454127, 0.3883342, 0.3228347, 0.1721232, 
    0.1181614, 0.236936, 0.2018438, 0.1486519, 0.1107567,
  0.09646098, 0.1900852, 0.2532487, 0.3943173, 0.4312745, 0.293145, 
    0.1728127, 0.2430339, 0.2410445, 0.2735488, 0.1719131, 0.1689532, 
    0.2314207, 0.1728874, 0.2345428, 0.2408119, 0.2896998, 0.2752235, 
    0.3168975, 0.2317625, 0.1875969, 0.3295005, 0.3546277, 0.4423125, 
    0.1176802, 0.1323653, 0.1329577, 0.1585038, 0.09903111,
  0.1692359, 0.2545, 0.4006061, 0.3783992, 0.2981757, 0.2894231, 0.2559308, 
    0.2946917, 0.2937089, 0.2853391, 0.3170182, 0.2715421, 0.3157772, 
    0.2463927, 0.2206377, 0.2409203, 0.2278556, 0.2490136, 0.2721464, 
    0.2794737, 0.2665414, 0.2860976, 0.2803827, 0.2514991, 0.2989512, 
    0.2334956, 0.2620372, 0.2146821, 0.2587439,
  0.2817624, 0.2376325, 0.19861, 0.2175823, 0.1667785, 0.1644484, 0.1683948, 
    0.2245651, 0.2571139, 0.3045219, 0.2259994, 0.2252871, 0.2329871, 
    0.2058624, 0.1387832, 0.1130422, 0.1416168, 0.1617481, 0.1899927, 
    0.155113, 0.2262429, 0.2208211, 0.1739348, 0.1589177, 0.08645701, 
    0.09640922, 0.1444507, 0.1449362, 0.2063468,
  0.08923073, 0.06630723, 0.06554338, 0.0977026, 0.1009471, 0.07026854, 
    0.09545758, 0.07954656, 0.1045919, 0.06254724, 0.0510022, 0.05814698, 
    0.03621767, 0.0454733, 0.1847535, 0.1503895, 0.1224279, 0.03850719, 
    0.0825708, 0.1222688, 0.1234244, 0.1398747, 0.0897531, 0.02302495, 
    0.0541533, 0.124749, 0.1489152, 0.137106, 0.09430678,
  0.03788286, -2.358046e-06, 0.08843642, 0.05640716, 0.0266226, 0.08269181, 
    0.06488951, 0.02723776, 0.001135294, 8.309196e-05, 9.569858e-05, 
    0.005657134, 0.01945569, 0.01332474, 0.1003613, 0.06558011, 0.05206835, 
    0.1825988, 0.06154851, 0.03533305, 0.07653822, 0.01514691, 0.0008766171, 
    1.455185e-05, 0.02080726, 0.06165011, 0.1062411, 0.03003345, 0.02737282,
  8.502112e-07, 0.0003416291, 0.10382, 0.01871576, 0.04360555, 0.02695252, 
    0.08452103, 0.02304104, 5.785825e-05, -4.458919e-07, 0.03044887, 
    0.01696698, 0.0668671, 0.0494661, 0.06288859, 0.07272173, 0.03989255, 
    0.03541375, 0.02837894, 0.04287809, 0.07731275, 0.02230242, 9.372263e-07, 
    3.095804e-05, 0.1008255, 0.1885125, 0.02518018, 0.02527898, 0.002299016,
  1.03168e-05, 0.01169257, 0.161426, 0.06995293, 0.06202295, 0.03450767, 
    0.08689524, 0.1129863, 0.01762469, 0.01347336, 0.04215661, 0.0141615, 
    0.0356796, 0.0659752, 0.03861158, 0.03503099, 0.02863193, 0.02775552, 
    0.024318, 0.01017584, 0.0001618792, -3.038679e-08, 1.662893e-05, 
    0.09890277, 0.1434878, 0.05144669, 0.04862593, 0.0002710716, 6.323978e-06,
  0.2460627, 0.02408592, 0.08711288, 0.1140318, 0.04825528, 0.0292154, 
    0.08137687, 0.02995144, 0.1437634, 0.1676464, 0.03890311, 0.009248627, 
    0.02851146, 0.03574349, 0.01665166, 0.01018175, 0.003714213, 0.002453734, 
    0.004983821, 0.000375438, 0.002323189, 0.02335495, 0.1020048, 0.180152, 
    0.1073475, 0.03282718, 0.04235585, 0.0308091, 0.0457863,
  1.969015e-07, 5.048155e-08, -1.058381e-06, 0.1099625, 0.07634914, 
    0.01913908, 0.01062243, 0.01736438, 0.08994789, 0.04383788, 0.07157752, 
    0.05629165, 0.06270568, 0.08311392, 0.1038577, 0.03584195, 0.05677002, 
    0.1027272, 0.1249642, 0.1042722, 0.05162179, 0.02192884, 0.05138022, 
    0.03789404, 0.05888426, 0.02330865, 0.00156021, 2.925526e-05, 
    -3.112889e-06,
  4.174723e-06, 4.487259e-07, 4.829385e-08, 0.02114003, 0.002632513, 
    0.02492052, 0.003977394, 3.853862e-05, 0.01483373, 0.102498, 0.1010763, 
    0.08824071, 0.03426348, 0.02976934, 0.04792033, 0.0323936, 0.03713387, 
    0.1273221, 0.04759178, 0.02177475, 0.02811191, 0.1001994, 0.03091495, 
    0.03529167, 0.04315561, 0.04858675, 0.07094814, 0.007551356, 5.367483e-06,
  -4.799696e-05, 0.03811714, 0.0431035, 0.07497398, 0.1050355, 0.1615928, 
    0.01706199, 0.03871686, 0.140263, 0.1766246, 0.09135985, 0.07612578, 
    0.09772956, 0.1085385, 0.08163656, 0.1791396, 0.1686178, 0.1240654, 
    0.1672986, 0.07868155, 0.1502647, 0.07110659, 0.02700579, 0.03590828, 
    0.06474967, 0.07748368, 0.05742225, 0.03164351, 0.06353332,
  0.04253766, 0.1048205, 0.1897825, 0.3042728, 0.1795558, 0.0622477, 
    0.191016, 0.04153967, 0.03620037, 0.06090531, 0.05372918, 0.2080434, 
    0.2204642, 0.2091288, 0.2256145, 0.2121201, 0.2002703, 0.1235059, 
    0.1852004, 0.2259712, 0.2666246, 0.07056883, 0.1705511, 0.1772969, 
    0.2667355, 0.2157217, 0.20749, 0.1465895, 0.2200388,
  0.1761356, 0.1711752, 0.09896603, 0.2174796, 0.1626782, 0.1865885, 
    0.173413, 0.150012, 0.1440633, 0.07648841, 0.07399492, 0.03732345, 
    0.3862104, 0.2888455, 0.3045958, 0.2304942, 0.1377198, 0.1026993, 
    0.1753107, 0.3291851, 0.1673707, 0.1476432, 0.2141178, 0.3039357, 
    0.1814441, 0.2900542, 0.3140196, 0.2399688, 0.2008725,
  0.2586773, 0.2644569, 0.2944352, 0.3571399, 0.3724687, 0.3852179, 
    0.3402721, 0.4325771, 0.2630412, 0.3869848, 0.4412845, 0.1281332, 
    0.4272165, 0.2778473, 0.3130849, 0.2986116, 0.2294254, 0.2157776, 
    0.221435, 0.253868, 0.2782318, 0.2045823, 0.1876241, 0.3081209, 
    0.2663692, 0.2584148, 0.2716489, 0.2861755, 0.2995718,
  0.348669, 0.3178771, 0.3245586, 0.3670106, 0.3322957, 0.43578, 0.5218698, 
    0.5049444, 0.277324, 0.3259352, 0.2699312, 0.2726244, 0.4575843, 
    0.3855758, 0.3825113, 0.2289002, 0.3046224, 0.4227488, 0.38606, 
    0.3860514, 0.389596, 0.1635854, 0.3275052, 0.1969984, 0.1628176, 
    0.4274367, 0.4791356, 0.4473016, 0.3374133,
  0.4706406, 0.3868977, 0.2256314, 0.1671701, 0.1720048, 0.1676295, 
    0.1251013, 0.1320164, 0.1565597, 0.2165859, 0.255201, 0.2797278, 
    0.3089806, 0.2780302, 0.2631108, 0.2852593, 0.2923437, 0.3101508, 
    0.3850311, 0.3690752, 0.3215136, 0.311054, 0.2794024, 0.1163287, 
    0.05819121, 0.05320961, 0.1375965, 0.2757534, 0.4208642,
  0.1573271, 0.1572207, 0.1571143, 0.1570079, 0.1569015, 0.1567951, 
    0.1566887, 0.1684985, 0.1778727, 0.1872469, 0.1966211, 0.2059954, 
    0.2153696, 0.2247438, 0.2194737, 0.2216336, 0.2237935, 0.2259534, 
    0.2281133, 0.2302732, 0.2324331, 0.2528448, 0.2414171, 0.2299894, 
    0.2185617, 0.2071339, 0.1957062, 0.1842785, 0.1574122,
  0.1193676, 0.1459998, 0.218403, 0.2123191, 0.1835776, 0.1627416, 0.2050741, 
    0.2729991, 0.2127258, 0.1934071, 0.2169859, 0.2103538, 0.2663773, 
    0.04321722, 0.06439593, 0.06596489, 0.0817231, 0.1731959, 0.1351658, 
    0.2057104, 0.2403258, 0.3975143, 0.3370927, 0.208867, 0.1884329, 
    0.2758003, 0.2065936, 0.1297985, 0.121151,
  0.114185, 0.1794062, 0.2611245, 0.3228616, 0.4071828, 0.307361, 0.1660084, 
    0.1880642, 0.2597677, 0.3068238, 0.2026023, 0.1561025, 0.2048631, 
    0.2046501, 0.2263296, 0.2351259, 0.3641627, 0.3956425, 0.3020279, 
    0.258951, 0.1959036, 0.3600222, 0.3315538, 0.4915627, 0.08572894, 
    0.1516422, 0.1653039, 0.1591385, 0.09546087,
  0.2491263, 0.2515515, 0.4308996, 0.3361838, 0.3621067, 0.2712716, 
    0.3054819, 0.2979677, 0.368985, 0.3411779, 0.3541467, 0.279786, 
    0.2967715, 0.2589489, 0.2452205, 0.2535143, 0.2379611, 0.2402882, 
    0.2941263, 0.3209433, 0.2813486, 0.3065102, 0.3396672, 0.3082023, 
    0.3456823, 0.3016682, 0.2711969, 0.2549337, 0.34232,
  0.290335, 0.2696993, 0.2399511, 0.2484097, 0.1947331, 0.1764508, 0.1816835, 
    0.2399025, 0.2946727, 0.3508532, 0.2951416, 0.255357, 0.2460541, 
    0.2243975, 0.1313348, 0.1099386, 0.1414706, 0.1944156, 0.2291704, 
    0.1890725, 0.2906605, 0.2611216, 0.1975103, 0.1578123, 0.06639588, 
    0.09011131, 0.1664712, 0.1630478, 0.2219287,
  0.1321424, 0.1380714, 0.1213137, 0.1487372, 0.1167646, 0.09221458, 
    0.1071775, 0.1030704, 0.1445708, 0.1016136, 0.06539666, 0.0638387, 
    0.04234842, 0.0497053, 0.2199616, 0.1559469, 0.1161577, 0.06152478, 
    0.1170159, 0.1306016, 0.1714001, 0.1518439, 0.120816, 0.02902992, 
    0.03930837, 0.1602928, 0.1777097, 0.1686415, 0.1022137,
  0.06533869, 1.915142e-05, 0.08161264, 0.05703582, 0.03500725, 0.09096488, 
    0.08643089, 0.05545574, 0.02041049, 0.001673243, 6.654268e-05, 
    0.001982884, 0.01780236, 0.03147329, 0.1170525, 0.08222122, 0.07444017, 
    0.1931386, 0.05211105, 0.03344521, 0.08614875, 0.02351071, 0.009103611, 
    2.063476e-05, 0.01834077, 0.06069991, 0.1074252, 0.04646887, 0.05307685,
  0.0003026413, -0.0003569874, 0.09850553, 0.02120984, 0.04020818, 0.0318813, 
    0.09160121, 0.03470584, 0.001831661, 5.574093e-08, 0.02766892, 
    0.01214314, 0.06265403, 0.0452481, 0.0696031, 0.07418165, 0.04690712, 
    0.02993445, 0.02706719, 0.03205522, 0.07581974, 0.04222342, 2.943306e-05, 
    0.0001479839, 0.09696683, 0.1838601, 0.03606512, 0.05891316, 0.01355222,
  1.367457e-05, 0.01634148, 0.1625789, 0.06374986, 0.05772768, 0.03268344, 
    0.06784385, 0.1049988, 0.0230264, 0.01773689, 0.04432163, 0.01136919, 
    0.03485379, 0.05256603, 0.03070451, 0.03119548, 0.02556805, 0.02447184, 
    0.02535924, 0.02358507, 0.01013925, 0.0009671993, 4.294369e-06, 
    0.09091777, 0.1222478, 0.04138456, 0.07061814, 0.009954589, 0.000419757,
  0.2168145, 0.0208943, 0.1048395, 0.1234104, 0.04284417, 0.02228836, 
    0.07198843, 0.02989477, 0.1546582, 0.1560971, 0.03622756, 0.009907275, 
    0.02682332, 0.02521026, 0.01812431, 0.0115707, 0.008328088, 0.009189074, 
    0.0143204, 0.008496248, 0.01065292, 0.01693384, 0.07258938, 0.16279, 
    0.08921774, 0.03014456, 0.03715743, 0.02667488, 0.03867088,
  4.404052e-08, 1.271286e-08, -1.873656e-08, 0.07132313, 0.1148891, 
    0.02440611, 0.01400252, 0.02445003, 0.0923635, 0.03731726, 0.05895374, 
    0.04415141, 0.06754287, 0.06911416, 0.1028558, 0.03481769, 0.05054439, 
    0.09684925, 0.1214072, 0.09683324, 0.04652435, 0.01982388, 0.05128061, 
    0.04183656, 0.05044708, 0.02816454, 0.005737544, -6.699892e-05, 
    -2.624307e-06,
  1.309589e-06, 2.904873e-07, 3.441499e-08, 0.07286454, 0.001533732, 
    0.05788564, 0.01253874, 0.005462918, 0.04582831, 0.1445973, 0.1083857, 
    0.102399, 0.03772242, 0.05894955, 0.06116859, 0.03520541, 0.03882689, 
    0.1271446, 0.06752443, 0.02536728, 0.03336327, 0.1443474, 0.03271633, 
    0.0315159, 0.03703713, 0.03798308, 0.07013288, 0.01148672, -9.406345e-07,
  0.002522142, 0.03206228, 0.07598595, 0.06414796, 0.1133963, 0.1462206, 
    0.007504114, 0.02503108, 0.1101775, 0.1626841, 0.09177104, 0.1595901, 
    0.1737755, 0.1560374, 0.1246165, 0.1810739, 0.1912758, 0.1201721, 
    0.2082841, 0.1260069, 0.17122, 0.08550252, 0.04013395, 0.08339477, 
    0.08796762, 0.08831734, 0.06731062, 0.05436277, 0.04618044,
  0.04196879, 0.1076959, 0.1815668, 0.3187139, 0.1560812, 0.08521915, 
    0.1755145, 0.03910792, 0.02896738, 0.04906539, 0.06125483, 0.3070614, 
    0.2316874, 0.2191246, 0.250834, 0.2263454, 0.2449837, 0.2250952, 
    0.2625735, 0.2586716, 0.2850297, 0.07102597, 0.1664603, 0.1922692, 
    0.2906346, 0.2185541, 0.2236478, 0.1713236, 0.2491652,
  0.2115071, 0.2067374, 0.1818269, 0.2543453, 0.1718495, 0.2229651, 
    0.1907154, 0.156864, 0.1036392, 0.08622248, 0.0802076, 0.03565592, 
    0.3941923, 0.3544572, 0.3339354, 0.2319775, 0.1459443, 0.1504931, 
    0.2416018, 0.331109, 0.2032126, 0.2182293, 0.2363718, 0.2991721, 
    0.2308966, 0.3399796, 0.3137826, 0.2438432, 0.2203217,
  0.2333516, 0.2605795, 0.3361734, 0.3247716, 0.3736808, 0.3309649, 
    0.3756184, 0.4057846, 0.3221793, 0.4083347, 0.4626573, 0.1313827, 
    0.4541848, 0.2776074, 0.3546502, 0.3273483, 0.2411539, 0.2147183, 
    0.225877, 0.2685552, 0.329566, 0.2474519, 0.2479766, 0.328395, 0.4076933, 
    0.2450782, 0.2858509, 0.2772977, 0.307268,
  0.3521969, 0.3199123, 0.3408702, 0.4467954, 0.4051408, 0.5108097, 
    0.5277484, 0.4482726, 0.2747589, 0.3889539, 0.267171, 0.314238, 
    0.5006534, 0.4489209, 0.40861, 0.2383714, 0.3202529, 0.466942, 0.3921163, 
    0.4026459, 0.4043459, 0.228705, 0.3752896, 0.2337851, 0.1607369, 
    0.4624613, 0.4893786, 0.4221838, 0.400362,
  0.4907472, 0.2697937, 0.1861986, 0.1979723, 0.176682, 0.1741168, 0.1482064, 
    0.1712508, 0.1558993, 0.2034538, 0.2340912, 0.3302178, 0.3316436, 
    0.3044325, 0.2785073, 0.2993907, 0.3352891, 0.3366207, 0.3947924, 
    0.4081534, 0.3258398, 0.376371, 0.2850011, 0.1146908, 0.0604673, 
    0.04654094, 0.1290182, 0.3160371, 0.4809149,
  0.1429823, 0.1426574, 0.1423325, 0.1420076, 0.1416827, 0.1413578, 
    0.1410329, 0.1482412, 0.1573051, 0.166369, 0.175433, 0.1844968, 
    0.1935608, 0.2026247, 0.2102686, 0.2140703, 0.2178719, 0.2216735, 
    0.2254752, 0.2292768, 0.2330785, 0.2543429, 0.2418022, 0.2292616, 
    0.2167209, 0.2041803, 0.1916396, 0.179099, 0.1432422,
  0.1207952, 0.1669818, 0.2251404, 0.2248784, 0.1802054, 0.1610184, 
    0.2029004, 0.2786167, 0.1925125, 0.1922144, 0.235708, 0.2421087, 
    0.2791563, 0.0294248, 0.1537487, 0.1541052, 0.2312962, 0.1898448, 
    0.1615429, 0.2129609, 0.229324, 0.4234637, 0.3593145, 0.1433994, 
    0.1413808, 0.2697079, 0.208025, 0.1177563, 0.1170388,
  0.1139866, 0.1553322, 0.2161858, 0.2612507, 0.356427, 0.3302541, 0.1596152, 
    0.1828592, 0.2761213, 0.2864452, 0.2622298, 0.1410994, 0.174693, 
    0.2037367, 0.2782342, 0.3224596, 0.4524652, 0.4672477, 0.321448, 
    0.2788209, 0.2561053, 0.3453134, 0.3508899, 0.4913896, 0.1010123, 
    0.1801892, 0.2317515, 0.2537826, 0.1430579,
  0.3198319, 0.3036489, 0.4590085, 0.418969, 0.4149943, 0.4095933, 0.4103582, 
    0.404805, 0.3430353, 0.3740462, 0.3803293, 0.3396465, 0.3188337, 
    0.3032728, 0.3027437, 0.2943859, 0.3182216, 0.3280161, 0.351454, 
    0.4024141, 0.3463837, 0.369545, 0.4062622, 0.3281505, 0.3640953, 
    0.3233243, 0.3301976, 0.3372716, 0.4625806,
  0.3423125, 0.3353901, 0.285013, 0.3022798, 0.2241687, 0.2040611, 0.2148412, 
    0.2856348, 0.374248, 0.4312202, 0.3734872, 0.2952558, 0.2583337, 
    0.2543513, 0.1653354, 0.1445423, 0.1826428, 0.2432512, 0.2858856, 
    0.2557164, 0.3380433, 0.2825266, 0.2496322, 0.1443599, 0.05727298, 
    0.1232616, 0.2312196, 0.2158715, 0.2435431,
  0.1468533, 0.2357355, 0.2124472, 0.1809591, 0.1713402, 0.1828452, 
    0.1856556, 0.1443264, 0.2002853, 0.1803853, 0.1518684, 0.08753031, 
    0.05459039, 0.05796772, 0.2129178, 0.1868908, 0.1512994, 0.1090737, 
    0.1380481, 0.1496838, 0.2336963, 0.224033, 0.2360589, 0.03332783, 
    0.04849527, 0.1886711, 0.2212334, 0.220536, 0.1501038,
  0.09041547, 0.002708408, 0.05415619, 0.06343105, 0.07701252, 0.1384273, 
    0.1008541, 0.09795176, 0.106135, 0.02624108, 7.252672e-05, 0.0009044393, 
    0.01539223, 0.09364954, 0.1372018, 0.1105766, 0.1113244, 0.1968223, 
    0.04997851, 0.0566355, 0.1192052, 0.07015067, 0.06117256, 1.823534e-05, 
    0.01552626, 0.05948246, 0.1161841, 0.06141495, 0.1018979,
  0.008610812, -0.0001796625, 0.07805146, 0.02415991, 0.04230076, 0.03783192, 
    0.09317036, 0.05350982, 0.01844623, 3.966267e-08, 0.0225529, 0.0106082, 
    0.06802365, 0.04062833, 0.07097206, 0.08215404, 0.05422438, 0.02913044, 
    0.0299921, 0.03351635, 0.05834749, 0.151163, 0.007662695, 0.0005061014, 
    0.09027094, 0.1679778, 0.05265354, 0.1295003, 0.0697622,
  0.001102232, 0.02905644, 0.1419783, 0.0633883, 0.0539709, 0.03445233, 
    0.0580632, 0.0782406, 0.02961432, 0.02772698, 0.04527325, 0.0119674, 
    0.04017939, 0.04388839, 0.02992792, 0.0323837, 0.02598383, 0.02526206, 
    0.03053058, 0.04302925, 0.0644224, 0.01998984, 0.001820595, 0.08142018, 
    0.1037785, 0.03424145, 0.07253806, 0.05386726, 0.01677511,
  0.1652502, 0.02799608, 0.07555727, 0.1121829, 0.04201559, 0.0202038, 
    0.06237193, 0.03187547, 0.136949, 0.146299, 0.03933451, 0.01346439, 
    0.02795758, 0.02509969, 0.02265402, 0.01490026, 0.008825433, 0.01028482, 
    0.0161276, 0.02754783, 0.02217099, 0.03429759, 0.04783753, 0.1390906, 
    0.08233571, 0.03033575, 0.03311084, 0.02472345, 0.02860177,
  4.244888e-09, 4.192483e-09, -1.776974e-07, 0.0497052, 0.1568109, 
    0.02890151, 0.01203504, 0.08510361, 0.1326078, 0.03423707, 0.05759929, 
    0.0421356, 0.06403928, 0.05988958, 0.09321759, 0.04277513, 0.04651401, 
    0.09214968, 0.1259786, 0.09080461, 0.04453683, 0.01998784, 0.05592541, 
    0.04930677, 0.04786301, 0.03849806, 0.0454678, -0.0001026936, 
    -1.364799e-06,
  4.309362e-07, 1.691508e-07, 1.194263e-08, 0.04614601, 0.0002215282, 
    0.07057878, 0.01093522, 0.02841857, 0.04472131, 0.2160025, 0.1331777, 
    0.1239316, 0.1005777, 0.08717457, 0.07315232, 0.06066873, 0.07057759, 
    0.1133041, 0.1002637, 0.09726975, 0.03110505, 0.190767, 0.05966303, 
    0.03826622, 0.04183916, 0.04558045, 0.08831294, 0.02016249, -7.249421e-06,
  0.02423444, 0.05643697, 0.1217081, 0.08187349, 0.1313674, 0.1278042, 
    0.001629922, 0.01782624, 0.08495982, 0.1728789, 0.1952084, 0.2344962, 
    0.1170346, 0.1594048, 0.1457025, 0.1905747, 0.2664361, 0.1267275, 
    0.2238845, 0.1631955, 0.1790543, 0.1093442, 0.08630688, 0.1227085, 
    0.1384242, 0.1040884, 0.09603719, 0.08932944, 0.04522318,
  0.05600181, 0.1010181, 0.1943016, 0.3131883, 0.1454449, 0.06394807, 
    0.1611375, 0.02700198, 0.02032305, 0.02905527, 0.1066407, 0.4063478, 
    0.23414, 0.2173579, 0.2480701, 0.2552443, 0.2855383, 0.3690785, 
    0.2130608, 0.3002394, 0.2774073, 0.08120531, 0.1898005, 0.2068387, 
    0.3123066, 0.2174221, 0.2608393, 0.2514625, 0.2557798,
  0.2057318, 0.2179818, 0.19598, 0.2791556, 0.2178818, 0.2180269, 0.2072331, 
    0.168167, 0.08110684, 0.07255659, 0.1114067, 0.04856235, 0.3905949, 
    0.2684519, 0.310757, 0.2136144, 0.1989946, 0.1715514, 0.3058136, 
    0.3498227, 0.1887334, 0.2013582, 0.275299, 0.3586318, 0.2326189, 
    0.3056799, 0.2916436, 0.2438672, 0.2228263,
  0.2192902, 0.2858527, 0.3700346, 0.3303849, 0.3527168, 0.3650293, 
    0.3481905, 0.4074836, 0.3486817, 0.446981, 0.4960161, 0.1251808, 
    0.4650656, 0.2450338, 0.4333497, 0.3872011, 0.2668548, 0.2123167, 
    0.2148121, 0.2807288, 0.4006089, 0.2596233, 0.2864073, 0.3615404, 
    0.6079923, 0.2130567, 0.2575405, 0.2439523, 0.2729049,
  0.3522773, 0.3578198, 0.3149264, 0.4786218, 0.4418451, 0.5437282, 
    0.5148022, 0.4484495, 0.2697638, 0.4213849, 0.3497541, 0.387327, 
    0.5536425, 0.4944289, 0.4502633, 0.2494084, 0.3540202, 0.4975799, 
    0.4155897, 0.4486643, 0.4135534, 0.3465121, 0.417081, 0.2411169, 
    0.1708255, 0.4623554, 0.5264595, 0.3964949, 0.4225251,
  0.3787297, 0.3041724, 0.1940642, 0.1302237, 0.1271736, 0.150383, 0.2129163, 
    0.2219559, 0.1706832, 0.2401786, 0.2974965, 0.3688285, 0.3903649, 
    0.3877098, 0.3048622, 0.3542581, 0.3764898, 0.4032559, 0.4449985, 
    0.4141674, 0.3198742, 0.3810665, 0.3147055, 0.1310985, 0.06899639, 
    0.04304955, 0.1376613, 0.3749257, 0.5684041,
  0.139992, 0.1406398, 0.1412876, 0.1419355, 0.1425833, 0.1432311, 0.1438789, 
    0.1444827, 0.1517099, 0.1589371, 0.1661644, 0.1733916, 0.1806189, 
    0.1878461, 0.2146063, 0.219774, 0.2249417, 0.2301094, 0.2352771, 
    0.2404448, 0.2456125, 0.2340844, 0.2210416, 0.2079988, 0.194956, 
    0.1819133, 0.1688705, 0.1558278, 0.1394737,
  0.1649158, 0.192272, 0.2288964, 0.2153431, 0.1721347, 0.151458, 0.1912434, 
    0.2622871, 0.1920159, 0.2191593, 0.2360831, 0.2707638, 0.2524018, 
    0.02694003, 0.2331444, 0.1780337, 0.2583918, 0.2524904, 0.1946152, 
    0.1988257, 0.2364561, 0.4003487, 0.3848343, 0.1446657, 0.1456947, 
    0.2591555, 0.1887923, 0.09337644, 0.1254601,
  0.1363726, 0.15462, 0.2182727, 0.2444372, 0.3167189, 0.3945317, 0.172277, 
    0.171301, 0.2723961, 0.269152, 0.3157206, 0.1523622, 0.1600531, 
    0.2051993, 0.2974316, 0.4301952, 0.4377662, 0.4773316, 0.4478658, 
    0.3534888, 0.3488068, 0.4019633, 0.467548, 0.5283496, 0.08967677, 
    0.1800191, 0.400194, 0.3237563, 0.1242898,
  0.4690627, 0.4377928, 0.5017321, 0.469042, 0.4775771, 0.4719398, 0.4351933, 
    0.418718, 0.368941, 0.4166836, 0.3704936, 0.409626, 0.3926573, 0.3784618, 
    0.3481699, 0.3699424, 0.3820329, 0.3757004, 0.3896533, 0.4025398, 
    0.3986076, 0.4141973, 0.4279745, 0.3820176, 0.4227276, 0.3510878, 
    0.4095781, 0.4475115, 0.5598329,
  0.3900896, 0.4066496, 0.3224316, 0.3927634, 0.3059049, 0.2934178, 0.277352, 
    0.3878719, 0.4423548, 0.4229454, 0.3870089, 0.3376264, 0.3006479, 
    0.2954586, 0.1996015, 0.2065873, 0.2422782, 0.3693229, 0.3393175, 
    0.3526638, 0.3224617, 0.3065718, 0.3138479, 0.146529, 0.05028762, 
    0.1746613, 0.2824602, 0.2961749, 0.3519614,
  0.2187359, 0.2220586, 0.2363722, 0.2598107, 0.2368042, 0.2985709, 
    0.2659855, 0.2382996, 0.3434231, 0.1886549, 0.1897429, 0.1423815, 
    0.09843998, 0.1624352, 0.2234792, 0.2576479, 0.1913657, 0.197658, 
    0.1995759, 0.2522019, 0.2827517, 0.294076, 0.2485127, 0.0381408, 
    0.0488801, 0.1903271, 0.3269925, 0.2893727, 0.2065453,
  0.2648869, 0.06687166, 0.04525752, 0.1108363, 0.1090548, 0.1783642, 
    0.116137, 0.1563475, 0.24634, 0.06217358, 0.0015739, 0.0003321992, 
    0.01069759, 0.1161438, 0.1897889, 0.106341, 0.1361662, 0.232132, 
    0.1101781, 0.06073482, 0.1168276, 0.1109331, 0.2469765, 6.431308e-05, 
    0.01191259, 0.06576791, 0.1204055, 0.09336617, 0.1745509,
  0.1688673, 7.286965e-05, 0.05919958, 0.0273383, 0.06771439, 0.05720356, 
    0.08373421, 0.1160286, 0.1952897, -3.070501e-07, 0.01505249, 0.006621064, 
    0.0800213, 0.04675969, 0.08509649, 0.07198688, 0.08153024, 0.03149794, 
    0.04005092, 0.04722626, 0.06348067, 0.2031522, 0.1442143, 0.001748887, 
    0.06455145, 0.1316104, 0.05747224, 0.1734917, 0.3170359,
  0.02468504, 0.04818331, 0.1120313, 0.05047609, 0.05505497, 0.04113167, 
    0.05086477, 0.07267393, 0.03955, 0.03470645, 0.04664466, 0.01760195, 
    0.04663078, 0.04491426, 0.03352197, 0.03872976, 0.03236232, 0.03548812, 
    0.04659233, 0.07254913, 0.1451234, 0.1071085, 0.01409418, 0.06719586, 
    0.08202986, 0.02466777, 0.1001207, 0.08438114, 0.08721156,
  0.1424664, 0.01088255, 0.0496823, 0.09718439, 0.05210559, 0.02260912, 
    0.06236048, 0.04361378, 0.1191845, 0.1394435, 0.04785014, 0.01896691, 
    0.03058308, 0.02870228, 0.04203683, 0.05359216, 0.009455564, 0.006850712, 
    0.03851017, 0.03040841, 0.05472078, 0.06572286, 0.03862253, 0.1000031, 
    0.07203522, 0.03452903, 0.0348438, 0.02685201, 0.02422576,
  1.205789e-09, 1.924487e-09, -1.267028e-07, 0.02850413, 0.1651068, 
    0.09943451, 0.003618354, 0.1038807, 0.135015, 0.0544938, 0.06866279, 
    0.04935627, 0.06023079, 0.09786288, 0.09642712, 0.05349704, 0.04934692, 
    0.1011772, 0.1182082, 0.07907644, 0.04633101, 0.01970896, 0.09322482, 
    0.06597766, 0.05726621, 0.061584, 0.2171307, 0.0103938, -1.272085e-06,
  1.39582e-07, 6.71162e-08, -1.420173e-08, 0.01417573, 2.06617e-05, 
    0.1771699, 0.003043965, 0.0320071, 0.03850297, 0.2962866, 0.1375214, 
    0.1793104, 0.1139851, 0.09578994, 0.1008501, 0.06191601, 0.1133291, 
    0.108478, 0.2011063, 0.2160939, 0.02402444, 0.2159262, 0.05945187, 
    0.04672243, 0.04930413, 0.06645222, 0.05887285, 0.005620019, -4.881897e-06,
  0.01122642, 0.1122028, 0.04734182, 0.08932119, 0.1409645, 0.1327983, 
    -0.002386534, 0.01165603, 0.06630995, 0.201374, 0.3751819, 0.1088088, 
    0.0768391, 0.09028632, 0.1162026, 0.2300074, 0.2921685, 0.1410578, 
    0.1874598, 0.1575954, 0.176249, 0.1465648, 0.1202608, 0.1276684, 
    0.1339938, 0.09329096, 0.137499, 0.1331291, 0.03716374,
  0.0797647, 0.1209404, 0.2444876, 0.3051013, 0.1247682, 0.06835625, 
    0.1542008, 0.009645517, 0.01791109, 0.02910431, 0.1900445, 0.289703, 
    0.1318341, 0.1525304, 0.2554395, 0.2444921, 0.3586146, 0.3867335, 
    0.1314804, 0.3158144, 0.2679089, 0.09454802, 0.2479156, 0.2683753, 
    0.3222874, 0.2255318, 0.2273239, 0.2220953, 0.2830825,
  0.2436554, 0.2746206, 0.1859587, 0.3277257, 0.2936273, 0.2276758, 
    0.2056081, 0.1886047, 0.06930107, 0.0943397, 0.1395353, 0.06050269, 
    0.3087624, 0.1892789, 0.2865764, 0.2274172, 0.3373098, 0.1401032, 
    0.235122, 0.3549874, 0.1690801, 0.2014114, 0.2705473, 0.4466675, 
    0.2784892, 0.2701094, 0.2456399, 0.2106226, 0.2095733,
  0.1946471, 0.3136942, 0.3687984, 0.3433889, 0.4211696, 0.381772, 0.3994241, 
    0.4685847, 0.4335299, 0.489556, 0.550475, 0.1623041, 0.5075421, 0.264928, 
    0.5376064, 0.3609824, 0.3361721, 0.2045189, 0.2561861, 0.2662833, 
    0.5102613, 0.3356, 0.2978154, 0.3813759, 0.5918018, 0.1364168, 0.1611602, 
    0.1877103, 0.235553,
  0.3530406, 0.3624978, 0.4074376, 0.4469577, 0.4780557, 0.6126721, 
    0.5508301, 0.5032353, 0.283614, 0.4270404, 0.3576204, 0.4528227, 
    0.600979, 0.539167, 0.514247, 0.2571232, 0.3936053, 0.4968189, 0.4302808, 
    0.5238625, 0.45648, 0.402954, 0.4479211, 0.2354759, 0.1384172, 0.4404655, 
    0.5681881, 0.3599485, 0.4706273,
  0.3355889, 0.2818578, 0.2366039, 0.2059266, 0.1743853, 0.1864277, 
    0.2945158, 0.3345875, 0.2288948, 0.3302527, 0.4136986, 0.3889938, 
    0.4274889, 0.4468655, 0.3843482, 0.4491529, 0.431854, 0.4503056, 
    0.4479458, 0.4105537, 0.3174022, 0.3819344, 0.3259059, 0.1501416, 
    0.06869079, 0.04952693, 0.1429456, 0.3985247, 0.5296386,
  0.2284337, 0.2263003, 0.2241669, 0.2220335, 0.2199001, 0.2177667, 
    0.2156333, 0.2060852, 0.2120168, 0.2179483, 0.2238798, 0.2298113, 
    0.2357429, 0.2416744, 0.2894132, 0.2980576, 0.3067019, 0.3153463, 
    0.3239906, 0.332635, 0.3412793, 0.3074223, 0.2949798, 0.2825374, 
    0.2700949, 0.2576524, 0.2452099, 0.2327675, 0.2301404,
  0.1803104, 0.2126425, 0.2503165, 0.1801268, 0.1728698, 0.1296751, 
    0.1651893, 0.236938, 0.2262778, 0.2324917, 0.2730833, 0.2727628, 
    0.3324935, 0.02605778, 0.2171256, 0.2676017, 0.231482, 0.3198364, 
    0.1905443, 0.1795614, 0.284063, 0.3659296, 0.4122165, 0.1712441, 
    0.2479823, 0.2835419, 0.1727381, 0.1083433, 0.1384572,
  0.1144739, 0.2001892, 0.2427802, 0.1998723, 0.2311142, 0.4126596, 
    0.1647895, 0.1396168, 0.2028087, 0.2172122, 0.2707647, 0.1825155, 
    0.1090942, 0.2377149, 0.3607327, 0.4672244, 0.4914085, 0.4481103, 
    0.4381558, 0.3562441, 0.3719461, 0.4445061, 0.5603921, 0.5479174, 
    0.07585377, 0.1795793, 0.3988177, 0.3750801, 0.1330966,
  0.5430575, 0.4691924, 0.5612427, 0.4993275, 0.5558177, 0.5317271, 
    0.4675333, 0.3754108, 0.3424065, 0.3783792, 0.3538291, 0.3909848, 
    0.515176, 0.4255652, 0.3776446, 0.394125, 0.4150979, 0.3857286, 0.455064, 
    0.3925573, 0.3985089, 0.4424856, 0.4217752, 0.4008311, 0.4352618, 
    0.4134625, 0.4483221, 0.5249321, 0.6517093,
  0.4159817, 0.4137787, 0.4129474, 0.4438939, 0.3670681, 0.4123498, 
    0.3783519, 0.461581, 0.4945585, 0.4066707, 0.3769449, 0.3510806, 
    0.3164854, 0.314643, 0.1788248, 0.252527, 0.3685335, 0.4316811, 
    0.3268329, 0.34211, 0.2965565, 0.3375871, 0.3284385, 0.1455909, 
    0.04603312, 0.1594832, 0.3221915, 0.3493164, 0.4343811,
  0.2258816, 0.1971228, 0.1404549, 0.2291948, 0.2603135, 0.319145, 0.4073135, 
    0.335608, 0.3404636, 0.2120606, 0.2239349, 0.135065, 0.09560524, 
    0.3454858, 0.2319423, 0.2757432, 0.3708396, 0.3415339, 0.3281999, 
    0.2871795, 0.2699116, 0.2651832, 0.2081974, 0.04568804, 0.05966241, 
    0.2214274, 0.3041085, 0.2313616, 0.2033623,
  0.3185573, 0.1102515, 0.03646556, 0.1571826, 0.114507, 0.1424614, 
    0.1450926, 0.198311, 0.3390561, 0.0532254, 0.02024033, 6.045549e-05, 
    0.003474966, 0.1098881, 0.1842375, 0.1406979, 0.09167748, 0.2251939, 
    0.0786346, 0.1150826, 0.1553327, 0.2310918, 0.3380491, 0.0003058598, 
    0.01112991, 0.1277401, 0.1179386, 0.129894, 0.1461403,
  0.5996327, -5.809449e-05, 0.0429358, 0.05526551, 0.07697211, 0.07281534, 
    0.09823348, 0.1039847, 0.2920283, -5.26319e-05, 0.01193732, 0.002352561, 
    0.1219569, 0.06213133, 0.09196045, 0.07709891, 0.07016594, 0.04113737, 
    0.04878091, 0.04658402, 0.04999417, 0.1325461, 0.6107917, 0.004771565, 
    0.04594173, 0.1257018, 0.05509234, 0.06790533, 0.3113842,
  0.2232237, 0.09783056, 0.08315845, 0.04438955, 0.05593508, 0.05100562, 
    0.05680071, 0.1018365, 0.1169295, 0.1516792, 0.08686551, 0.1284411, 
    0.0615232, 0.06750197, 0.05222259, 0.04653803, 0.0391276, 0.04583609, 
    0.03899852, 0.03550559, 0.2089845, 0.3079985, 0.03842745, 0.04607248, 
    0.06235346, 0.01544114, 0.1037365, 0.09403887, 0.2452561,
  0.08825669, 0.002727506, 0.02907157, 0.08622517, 0.07972956, 0.05586237, 
    0.1440739, 0.1270611, 0.1139855, 0.1304837, 0.1044234, 0.1949917, 
    0.05282458, 0.09007447, 0.08439624, 0.09883605, 0.03184953, 0.01255059, 
    0.04667623, 0.04441192, 0.09509207, 0.09056131, 0.04434649, 0.06170124, 
    0.0439739, 0.04111379, 0.04125365, 0.05752626, 0.02887224,
  7.493967e-10, 8.096843e-10, -3.631114e-08, 0.0139029, 0.1828535, 0.1158631, 
    0.0009064478, 0.09163733, 0.1245477, 0.06170553, 0.06743144, 0.0503002, 
    0.05002231, 0.07513095, 0.1383705, 0.09994942, 0.06808928, 0.1076547, 
    0.1135732, 0.09037714, 0.05110485, 0.04358995, 0.2693663, 0.1267916, 
    0.05260935, 0.02762095, 0.0938276, 0.0003332732, -1.968917e-06,
  4.603802e-08, 2.388639e-08, 5.945848e-10, 0.004180306, 1.746713e-05, 
    0.06934343, 0.001617616, 0.01590511, 0.03422423, 0.3471038, 0.1622706, 
    0.1482474, 0.07082355, 0.06173973, 0.06457511, 0.03086983, 0.06675711, 
    0.1014794, 0.1687587, 0.203013, 0.0242474, 0.2537005, 0.06001568, 
    0.03602975, 0.03448987, 0.02588241, 0.0355695, 0.000741057, -4.409432e-07,
  0.002715837, 0.07160968, 0.009369398, 0.07600144, 0.1258637, 0.1572455, 
    -0.003930359, 0.008075952, 0.04681542, 0.2234076, 0.2250961, 0.04777342, 
    0.05782291, 0.05541514, 0.0816453, 0.213775, 0.2050702, 0.128711, 
    0.1998423, 0.1145228, 0.1588041, 0.2059781, 0.1421546, 0.1667646, 
    0.157368, 0.118113, 0.07853253, 0.2211792, 0.02235555,
  0.05619591, 0.1303589, 0.2600928, 0.3094412, 0.1085793, 0.1015387, 
    0.1679965, 0.001917516, 0.01204477, 0.03248976, 0.251144, 0.1290224, 
    0.07491664, 0.1139983, 0.2595304, 0.3143714, 0.4457535, 0.2524664, 
    0.07067285, 0.3215541, 0.2384223, 0.08510296, 0.3303992, 0.2788618, 
    0.3017355, 0.2137383, 0.2741265, 0.1970839, 0.3115269,
  0.300683, 0.3013675, 0.2676584, 0.4436139, 0.3338504, 0.2646094, 0.2188704, 
    0.2231033, 0.06272525, 0.1404407, 0.1756175, 0.05907599, 0.1987099, 
    0.1201791, 0.289234, 0.2777031, 0.355548, 0.3075646, 0.1636391, 
    0.3527843, 0.1592448, 0.2297254, 0.2792113, 0.4987094, 0.3067131, 
    0.2228753, 0.2161143, 0.1973553, 0.2016706,
  0.1804847, 0.3328221, 0.4535224, 0.4287468, 0.5600166, 0.4275266, 
    0.5143635, 0.5579001, 0.4966814, 0.532548, 0.6511488, 0.2151851, 
    0.4989204, 0.2368951, 0.5148986, 0.3369011, 0.3857825, 0.2080172, 
    0.3302078, 0.2603354, 0.5986494, 0.4163448, 0.3560033, 0.3779821, 
    0.435395, 0.07316172, 0.1075369, 0.157512, 0.2032045,
  0.3217218, 0.3500674, 0.3681572, 0.3719883, 0.5333812, 0.6674932, 
    0.6442552, 0.5360028, 0.2794888, 0.4624401, 0.3605327, 0.4995979, 
    0.6313503, 0.5678827, 0.5325522, 0.250019, 0.3948422, 0.4885337, 
    0.4354776, 0.6417178, 0.4916143, 0.4621131, 0.4444389, 0.2350549, 
    0.1686033, 0.4175056, 0.5834892, 0.3228665, 0.4337342,
  0.3559289, 0.2163685, 0.2800208, 0.1984946, 0.228703, 0.2849211, 0.4331814, 
    0.4513436, 0.4168485, 0.4090486, 0.4537019, 0.4066097, 0.4763144, 
    0.5109651, 0.4351898, 0.4787766, 0.4839132, 0.4880942, 0.568164, 
    0.501785, 0.4003983, 0.4189211, 0.358607, 0.1963184, 0.07764361, 
    0.04769662, 0.1481085, 0.3806622, 0.6084014,
  0.3125763, 0.3141736, 0.315771, 0.3173684, 0.3189658, 0.3205632, 0.3221605, 
    0.3024939, 0.3076315, 0.3127691, 0.3179068, 0.3230444, 0.3281821, 
    0.3333197, 0.4003515, 0.4077883, 0.4152251, 0.4226619, 0.4300987, 
    0.4375354, 0.4449722, 0.3809198, 0.366748, 0.3525762, 0.3384044, 
    0.3242326, 0.3100608, 0.295889, 0.3112984,
  0.2280552, 0.2292765, 0.2445742, 0.1871328, 0.1854486, 0.08537415, 
    0.1229788, 0.2302245, 0.3166682, 0.2744124, 0.300051, 0.2754445, 
    0.3270495, 0.02473152, 0.1359739, 0.1796233, 0.1579917, 0.3023468, 
    0.1907725, 0.1519949, 0.2718787, 0.3595006, 0.3632056, 0.1885285, 
    0.2945354, 0.3130756, 0.1635, 0.09693182, 0.1155696,
  0.2392401, 0.1917227, 0.2720483, 0.1943942, 0.1654418, 0.3554642, 
    0.1219296, 0.1047375, 0.1374947, 0.1493974, 0.2038306, 0.196746, 
    0.09165908, 0.2254135, 0.4199403, 0.4649218, 0.4818621, 0.4403903, 
    0.3870042, 0.327254, 0.3802014, 0.5185705, 0.5606615, 0.5957891, 
    0.08155001, 0.2464829, 0.3340981, 0.41687, 0.2772468,
  0.5099866, 0.4761165, 0.5756388, 0.5547442, 0.578559, 0.5779119, 0.5019621, 
    0.3326996, 0.3340626, 0.3334743, 0.3462975, 0.3925671, 0.5538633, 
    0.4871644, 0.3430731, 0.4035835, 0.4114996, 0.4347917, 0.4493842, 
    0.3599213, 0.3434887, 0.3988714, 0.425088, 0.4028251, 0.4379357, 
    0.4345261, 0.5283355, 0.617472, 0.6280558,
  0.4257083, 0.4086681, 0.4256824, 0.3921531, 0.3611373, 0.4271247, 
    0.4512414, 0.5348817, 0.4718961, 0.374068, 0.3465215, 0.3390785, 
    0.3129165, 0.3156327, 0.133526, 0.2522963, 0.3742329, 0.3954982, 
    0.3433028, 0.3037397, 0.2680967, 0.31386, 0.3025415, 0.1417007, 
    0.04378211, 0.1316989, 0.3367293, 0.3658222, 0.4579245,
  0.1766668, 0.1237311, 0.09498245, 0.2146043, 0.2414701, 0.1910359, 
    0.3713927, 0.2575713, 0.2177351, 0.1829605, 0.1852141, 0.09783701, 
    0.09450126, 0.2414324, 0.2599825, 0.2786266, 0.2558951, 0.2426196, 
    0.3493594, 0.2598187, 0.233142, 0.267983, 0.1816006, 0.06137617, 
    0.07412958, 0.2149494, 0.2392521, 0.1827742, 0.1549279,
  0.1712636, 0.09008916, 0.02517751, 0.1750682, 0.07464986, 0.09222843, 
    0.1593975, 0.1553751, 0.151499, 0.02087777, 0.02334451, -7.246324e-06, 
    0.0005731249, 0.1008819, 0.1482644, 0.0938025, 0.07026652, 0.213171, 
    0.06022344, 0.1653443, 0.1408994, 0.10786, 0.1892895, 0.01342437, 
    0.006929716, 0.1075946, 0.115837, 0.07915865, 0.08678787,
  0.3379984, 0.02796143, 0.03236983, 0.0896408, 0.02143212, 0.06808307, 
    0.04200592, 0.02902363, 0.2240772, 3.639025e-06, 0.01192691, 
    0.0007768433, 0.04708281, 0.04803073, 0.0765733, 0.05416064, 0.09067146, 
    0.04500169, 0.03488937, 0.006231171, 0.00836389, 0.03839104, 0.4382023, 
    0.09520882, 0.03238049, 0.1112089, 0.01198266, 0.01375559, 0.1214925,
  0.461679, 0.1881702, 0.05520494, 0.04549569, 0.03433821, 0.05623263, 
    0.04826142, 0.05835003, 0.05961516, 0.06372455, 0.02747006, 0.0193682, 
    0.04318707, 0.0288458, 0.03038463, 0.01549242, 0.01972416, 0.02089874, 
    0.007148963, 0.007379268, 0.05546956, 0.2550837, 0.4678085, 0.03009571, 
    0.04331134, 0.01339036, 0.02703448, 0.03393229, 0.2109345,
  0.07253713, 0.001056486, 0.02037134, 0.07273693, 0.1045238, 0.06218594, 
    0.06037184, 0.0565319, 0.07199293, 0.1138345, 0.02520631, 0.1221284, 
    0.01523313, 0.02841262, 0.02979118, 0.04410859, 0.08428555, 0.03685194, 
    0.01140078, 0.04340659, 0.08959319, 0.15323, 0.09839348, 0.0390107, 
    0.01996902, 0.01799523, 0.03986115, 0.1469762, 0.03760028,
  6.900134e-10, 4.704951e-10, -3.129797e-09, 0.01255849, 0.2070705, 
    0.02538232, 0.0001556786, 0.01964661, 0.07109036, 0.03584836, 0.05605901, 
    0.03871509, 0.02224152, 0.02947089, 0.05552513, 0.06579664, 0.04173733, 
    0.07372927, 0.09008002, 0.09818148, 0.06879558, 0.04521226, 0.4144341, 
    0.1582467, 0.026071, 0.007055003, 0.02760839, 9.720532e-06, -2.606831e-06,
  2.211029e-08, 9.20478e-09, 1.997198e-11, 0.0006244104, 0.00393066, 
    0.01794975, 0.001202567, 0.002407887, 0.0368559, 0.3111848, 0.08298477, 
    0.06325625, 0.01796707, 0.02556788, 0.01861485, 0.02394226, 0.03417577, 
    0.09115534, 0.09807835, 0.1792065, 0.01963659, 0.2412086, 0.008128444, 
    0.01464501, 0.01970227, 0.006801297, 0.009386749, 0.0002607907, 
    -1.856331e-08,
  0.00019242, 0.03548701, 0.001425359, 0.05233351, 0.109933, 0.125358, 
    -0.003053508, 0.00451841, 0.03132866, 0.2078854, 0.1232644, 0.02583796, 
    0.04042388, 0.0355706, 0.06272476, 0.1904647, 0.1858635, 0.1042561, 
    0.1729035, 0.1007833, 0.1390507, 0.2716291, 0.1480871, 0.1626324, 
    0.12398, 0.08203511, 0.03973821, 0.1315628, 0.009814088,
  0.05126185, 0.07497014, 0.1996172, 0.3059573, 0.05566726, 0.1106807, 
    0.1755375, 0.0002682345, 0.00946665, 0.05258636, 0.2517255, 0.06769638, 
    0.03762792, 0.08800022, 0.2612371, 0.3254175, 0.3961721, 0.1254981, 
    0.05735144, 0.3205319, 0.2171906, 0.08873023, 0.3411767, 0.2484298, 
    0.2399005, 0.2361884, 0.2517098, 0.1751232, 0.2769058,
  0.3028971, 0.3269869, 0.2942822, 0.5498402, 0.3784668, 0.2667837, 
    0.2609488, 0.244319, 0.06208131, 0.171051, 0.1944776, 0.07383571, 
    0.1253116, 0.07785892, 0.2862245, 0.3484688, 0.2982008, 0.2536468, 
    0.1205992, 0.3777374, 0.1742969, 0.2157669, 0.2626703, 0.4760827, 
    0.3105676, 0.1918374, 0.1813105, 0.1886213, 0.1957579,
  0.143878, 0.3515781, 0.5436881, 0.5089952, 0.5810483, 0.4972355, 0.624009, 
    0.7036306, 0.5859006, 0.6156796, 0.7178912, 0.2771201, 0.4673237, 
    0.216321, 0.4680389, 0.3545713, 0.4388925, 0.2075232, 0.3506151, 
    0.2629147, 0.668941, 0.3842469, 0.4070562, 0.3667913, 0.3416734, 
    0.04120275, 0.09000796, 0.1323621, 0.1837097,
  0.2602202, 0.297581, 0.3347107, 0.3011573, 0.5478455, 0.7212987, 0.7311115, 
    0.5722034, 0.2887388, 0.4760194, 0.3769706, 0.5384997, 0.6340977, 
    0.6299987, 0.5181241, 0.2551984, 0.3605155, 0.4277106, 0.4799439, 
    0.6995789, 0.4725061, 0.4642466, 0.4631885, 0.2663989, 0.1455841, 
    0.4246604, 0.5891558, 0.3127275, 0.3783084,
  0.3690292, 0.1896686, 0.3167672, 0.2229825, 0.2766505, 0.4278438, 
    0.4947702, 0.5225357, 0.4705015, 0.4574571, 0.4896799, 0.4917881, 
    0.5685384, 0.5779207, 0.4795519, 0.5332366, 0.5143561, 0.4889507, 
    0.5641081, 0.5067787, 0.4981211, 0.4403786, 0.3954664, 0.2132103, 
    0.1084468, 0.04929949, 0.1530598, 0.3846885, 0.667814,
  0.3295633, 0.3325611, 0.3355589, 0.3385566, 0.3415544, 0.3445522, 0.34755, 
    0.3310375, 0.3360687, 0.3410999, 0.3461312, 0.3511624, 0.3561936, 
    0.3612248, 0.416387, 0.4208802, 0.4253734, 0.4298666, 0.4343598, 
    0.4388531, 0.4433463, 0.3969068, 0.3843845, 0.3718623, 0.3593401, 
    0.3468179, 0.3342957, 0.3217734, 0.3271651,
  0.2022519, 0.2286711, 0.1941483, 0.1850928, 0.1649441, 0.05366306, 
    0.08628345, 0.2204107, 0.3439411, 0.3118029, 0.278275, 0.2136529, 
    0.2571053, 0.007266257, 0.1012068, 0.1662728, 0.1518193, 0.2498984, 
    0.1599903, 0.1176513, 0.2003318, 0.3006281, 0.329319, 0.2000854, 
    0.2117284, 0.2832466, 0.1293902, 0.06665768, 0.114607,
  0.2108014, 0.1560401, 0.2840167, 0.180299, 0.09925073, 0.2857799, 
    0.1034042, 0.08006629, 0.09709747, 0.09217387, 0.1306223, 0.1583062, 
    0.05371436, 0.2295756, 0.4316573, 0.4088801, 0.4433587, 0.3923121, 
    0.3463289, 0.3522798, 0.3938642, 0.5314236, 0.5623212, 0.6157995, 
    0.08725522, 0.3339644, 0.3437322, 0.4172786, 0.3724767,
  0.4497033, 0.4633175, 0.5490188, 0.548096, 0.516495, 0.5300608, 0.4832829, 
    0.2908978, 0.305041, 0.307963, 0.3144639, 0.3677429, 0.5371845, 
    0.4334871, 0.3085122, 0.37283, 0.3695941, 0.4460026, 0.4040459, 
    0.3018977, 0.3109046, 0.3422286, 0.4085309, 0.3868196, 0.4064898, 
    0.4504938, 0.5729032, 0.6107128, 0.5603491,
  0.3842132, 0.3650365, 0.3683336, 0.3415082, 0.3482185, 0.4114863, 
    0.4341052, 0.4552308, 0.429386, 0.3644606, 0.3025205, 0.3388075, 
    0.2802572, 0.317423, 0.1246443, 0.2548618, 0.3301635, 0.3320862, 
    0.2875138, 0.2535151, 0.2343173, 0.2729825, 0.2670614, 0.1309608, 
    0.04392637, 0.1258492, 0.3350789, 0.3462042, 0.4009737,
  0.1360931, 0.08181478, 0.06018951, 0.2013836, 0.2261921, 0.1745424, 
    0.270912, 0.2011641, 0.1552458, 0.1359181, 0.1657063, 0.07923001, 
    0.04897722, 0.1434991, 0.2643221, 0.2230226, 0.1689678, 0.163482, 
    0.2841175, 0.2403192, 0.2305126, 0.2475702, 0.1411206, 0.07417175, 
    0.1039883, 0.1771194, 0.2455534, 0.1956594, 0.1350833,
  0.08780055, 0.06930084, 0.02233174, 0.1247783, 0.05952472, 0.05663918, 
    0.08594793, 0.04992185, 0.05820755, 0.007290572, 0.01827239, 
    0.0002899484, -0.0008917333, 0.03657469, 0.138429, 0.04898308, 
    0.06633396, 0.1878432, 0.1197436, 0.09612014, 0.07396727, 0.02766454, 
    0.07153429, 0.02578776, 0.002077837, 0.06452874, 0.1019047, 0.02209027, 
    0.05022398,
  0.1155917, 0.07292597, 0.02249076, 0.02291481, -0.0004162929, 0.02100853, 
    0.01453155, 0.005024746, 0.1111568, 0.002400763, 0.00906137, 
    0.0006338623, 0.01148603, 0.03021571, 0.0562764, 0.03097504, 0.03543384, 
    0.02158544, 0.005177921, 8.785585e-05, 0.0003358103, 0.01003225, 0.15586, 
    0.3000222, 0.0316353, 0.1039327, 0.0008073648, 0.00347007, 0.03763975,
  0.1604539, 0.1064383, 0.03991181, 0.06566846, 0.01330535, 0.01774397, 
    0.02066365, 0.0258501, 0.02475683, 0.01039546, 0.01049977, 0.005529531, 
    0.01644534, 0.01245715, 0.00609798, 0.002909299, 0.001335035, 
    0.002046806, 0.0002373634, 0.0003645795, 0.01476658, 0.07840011, 
    0.3840621, 0.02439808, 0.0310702, 0.01210267, 0.0003035129, 0.003973005, 
    0.05425324,
  0.08371715, 0.0006640821, 0.0152765, 0.06892644, 0.03636793, 0.01333932, 
    0.02918219, 0.01388936, 0.06073247, 0.08762078, 0.01508202, 0.02089983, 
    0.006901333, 0.005484137, 0.004064974, 0.005791517, 0.01459234, 
    0.01353982, 0.001717827, 0.01076908, 0.06756366, 0.3895484, 0.3192225, 
    0.03297078, 0.01111369, 0.003044019, 0.01492616, 0.07590909, 0.05688949,
  6.523075e-10, 3.697856e-10, 2.554435e-09, 0.01691705, 0.1930974, 
    0.005948095, -0.00137779, 0.004720032, 0.03140783, 0.01357914, 
    0.02682681, 0.009351988, 0.008980603, 0.008188566, 0.02525225, 
    0.02933891, 0.02642029, 0.03705552, 0.06813483, 0.05180325, 0.01994593, 
    0.01033247, 0.3641875, 0.1222185, 0.0117486, 0.00132853, 0.009408977, 
    -1.280472e-05, -1.401626e-06,
  1.258838e-08, 5.175152e-09, -7.143064e-10, -0.0002204997, 0.004597791, 
    0.004748222, 0.002710486, 0.0009306835, 0.03441216, 0.2363771, 
    0.03649225, 0.02834671, 0.00720934, 0.003080246, 0.005994019, 
    0.002681458, 0.01888996, 0.06383917, 0.04850008, 0.153507, 0.01175878, 
    0.2548681, 0.001084363, -0.001763302, 0.01192358, 0.0006698674, 
    0.003018591, 0.0001277388, 2.823068e-08,
  -3.896403e-05, 0.03015351, 0.000910393, 0.02443059, 0.09775325, 0.08592354, 
    -0.003572922, 0.002574249, 0.01952791, 0.1999263, 0.07533798, 0.01549394, 
    0.02699765, 0.0249334, 0.04655794, 0.1447309, 0.1798407, 0.0478591, 
    0.1052735, 0.1082514, 0.124285, 0.2647107, 0.1344924, 0.08451328, 
    0.08809792, 0.06555609, 0.01557128, 0.04408988, 0.003795119,
  0.02803309, 0.03712441, 0.1487213, 0.3142738, 0.02989749, 0.07804669, 
    0.1776707, 0.000265882, 0.003115661, 0.07331926, 0.241315, 0.04071684, 
    0.02520005, 0.06935988, 0.2285397, 0.2640647, 0.3153253, 0.1062087, 
    0.06390844, 0.3112228, 0.1910761, 0.08697234, 0.3111913, 0.2415952, 
    0.19112, 0.2098531, 0.2113407, 0.1435465, 0.2423697,
  0.2532677, 0.3544867, 0.3158791, 0.5872202, 0.3819738, 0.2788328, 
    0.2106652, 0.2363785, 0.05720509, 0.173264, 0.1611964, 0.1089739, 
    0.08599643, 0.05505871, 0.271847, 0.3662895, 0.277354, 0.14742, 
    0.09579751, 0.4003947, 0.1677983, 0.195157, 0.2396794, 0.4927946, 
    0.3452128, 0.174783, 0.1622091, 0.158832, 0.2004489,
  0.1086822, 0.4073681, 0.5450824, 0.5634169, 0.6265302, 0.5459539, 
    0.6428558, 0.7711727, 0.6551042, 0.6654674, 0.7679568, 0.3787071, 
    0.3952834, 0.1802903, 0.4106165, 0.3898535, 0.5034795, 0.1975199, 
    0.3825078, 0.2583806, 0.7638082, 0.4039072, 0.4575391, 0.3152599, 
    0.2931722, 0.02486357, 0.07377063, 0.09888443, 0.1514303,
  0.2187676, 0.2347317, 0.3420016, 0.2060833, 0.4885031, 0.6763076, 
    0.7796678, 0.5268064, 0.3231072, 0.5111326, 0.4147753, 0.568942, 
    0.6763239, 0.6898463, 0.4997528, 0.2527753, 0.3552568, 0.3419772, 
    0.4869844, 0.644676, 0.4104216, 0.5152307, 0.4905282, 0.2918752, 
    0.1806656, 0.4226441, 0.5961329, 0.2554574, 0.3377195,
  0.3838598, 0.1574054, 0.3476948, 0.2893218, 0.3892764, 0.5696724, 
    0.5566589, 0.551356, 0.471912, 0.5373279, 0.5755804, 0.6211079, 
    0.6971186, 0.6748452, 0.5723839, 0.5775915, 0.5413892, 0.5307474, 
    0.6177455, 0.5396904, 0.5723886, 0.4709461, 0.4428477, 0.2280712, 
    0.1085853, 0.04922092, 0.1542486, 0.3643622, 0.66197,
  0.2736285, 0.2775607, 0.2814929, 0.285425, 0.2893572, 0.2932894, 0.2972216, 
    0.2569009, 0.2608455, 0.2647901, 0.2687347, 0.2726793, 0.2766239, 
    0.2805685, 0.3659922, 0.3679372, 0.3698822, 0.3718272, 0.3737721, 
    0.3757171, 0.377662, 0.3322157, 0.3223939, 0.3125722, 0.3027504, 
    0.2929287, 0.283107, 0.2732852, 0.2704827,
  0.1516945, 0.1765874, 0.1493648, 0.1649658, 0.1105111, 0.03672484, 
    0.06342629, 0.1831083, 0.2739534, 0.227652, 0.192617, 0.1325723, 
    0.150309, -0.001438049, 0.0907087, 0.1794816, 0.1034727, 0.1864313, 
    0.126364, 0.07798779, 0.138804, 0.2224634, 0.2876948, 0.1839366, 
    0.1336068, 0.1884205, 0.09257313, 0.04486627, 0.0827252,
  0.1427379, 0.1369161, 0.2082799, 0.1241636, 0.05624159, 0.2456754, 
    0.09491417, 0.05964746, 0.06311285, 0.06233777, 0.0744651, 0.10944, 
    0.04383465, 0.222178, 0.4320515, 0.3374864, 0.3989398, 0.3424414, 
    0.3217572, 0.3225268, 0.3593823, 0.4843914, 0.5428815, 0.599174, 
    0.1040952, 0.3155382, 0.3287732, 0.3585872, 0.2768202,
  0.3845668, 0.4109573, 0.4856548, 0.453976, 0.4366787, 0.443515, 0.4313289, 
    0.2435324, 0.2326154, 0.2673212, 0.2753128, 0.3215415, 0.4697237, 
    0.3697305, 0.2543399, 0.3277611, 0.3294678, 0.408861, 0.3528282, 
    0.2596991, 0.2668248, 0.2920398, 0.3376267, 0.3176161, 0.3479038, 
    0.460867, 0.5291284, 0.5468906, 0.5382604,
  0.3291747, 0.3076281, 0.327654, 0.3406712, 0.3528844, 0.3693774, 0.3866777, 
    0.366232, 0.3720143, 0.333722, 0.2560454, 0.2890863, 0.2439872, 
    0.2704673, 0.1296758, 0.2103132, 0.257216, 0.279628, 0.2206149, 
    0.1900275, 0.1971117, 0.2601773, 0.2206399, 0.1107501, 0.04619027, 
    0.1258511, 0.2993831, 0.3229018, 0.3362905,
  0.1018983, 0.05050637, 0.03400311, 0.1798995, 0.1932087, 0.1538377, 
    0.2115376, 0.1473652, 0.1218393, 0.09899861, 0.1145303, 0.04576647, 
    0.0320155, 0.106492, 0.2466336, 0.1740612, 0.1267954, 0.1202533, 
    0.2225882, 0.2290401, 0.2134228, 0.1914363, 0.1246715, 0.09436459, 
    0.1026896, 0.1632986, 0.2268108, 0.1976457, 0.1123365,
  0.04155581, 0.03544429, 0.01635719, 0.06742373, 0.03627497, 0.03711449, 
    0.05629623, 0.01777121, 0.02359042, 0.008916333, 0.008705634, 
    0.0003186711, 0.0003605589, 0.01014726, 0.1145897, 0.03030085, 
    0.05350367, 0.1561038, 0.1530799, 0.04469575, 0.03639243, 0.01156934, 
    0.02845309, 0.01174585, 0.0005973195, 0.03802846, 0.05891495, 
    0.005804229, 0.009353325,
  0.04154225, 0.09322146, 0.01411915, 0.008575481, -0.003498661, 0.003617924, 
    0.004795783, 0.001757089, 0.05142686, 0.01768159, 0.006651307, 
    0.0002410413, 0.004695059, 0.01015933, 0.03897994, 0.009515059, 
    0.01079159, 0.005589331, 0.0007283993, 1.885792e-05, 0.0001317381, 
    0.003556437, 0.05366697, 0.1712211, 0.02836792, 0.0989892, 0.00013249, 
    0.001576435, 0.01257611,
  0.05769842, 0.0243062, 0.0281535, 0.06555305, 0.00899271, 0.002278402, 
    0.00869602, 0.009349156, 0.004098325, 0.0016245, 0.005322148, 
    0.001441152, 0.004788246, 0.003769334, 0.0006839348, 0.0005478502, 
    8.865289e-05, 0.0001057031, 5.810008e-05, 0.0001411983, 0.006059109, 
    0.02917313, 0.1262306, 0.02571342, 0.02787876, 0.01221543, -0.0008954172, 
    0.001449525, 0.01840927,
  0.0620007, 0.0003726309, 0.009482395, 0.0623761, 0.00913647, 0.001973062, 
    0.02496668, 0.005187331, 0.06140106, 0.08340404, 0.01232197, 0.007373847, 
    0.000647377, 0.001266497, 0.001101362, 0.00174337, 0.003740041, 
    0.003070623, 0.0007490008, 0.00102748, 0.02551517, 0.2012808, 0.1753149, 
    0.03354934, 0.007950963, 0.0003189907, 0.006239448, 0.01238742, 0.00675367,
  6.298536e-10, 3.361431e-10, 3.345543e-09, 0.0118992, 0.1498199, 
    0.002173875, -0.002350142, 0.002056419, 0.01544348, 0.002098915, 
    0.007166451, 0.002893937, 0.005774042, 0.001811997, 0.008298939, 
    0.006047116, 0.009512131, 0.01299923, 0.03539779, 0.02351422, 
    0.006006735, 0.002748409, 0.2472305, 0.07744235, 0.005002226, 
    0.0002779005, 0.004708558, -1.155644e-05, -5.969128e-07,
  1.000065e-08, 5.532725e-09, -3.634146e-09, -0.0002102913, 0.001244822, 
    0.002090347, 0.003230298, 0.0005117402, 0.03481696, 0.1411954, 
    0.01369833, 0.01249134, 0.001607749, 0.0007057296, 0.00136334, 
    0.0007942665, 0.007210285, 0.03648538, 0.0190749, 0.09126756, 
    0.007223485, 0.1833885, 0.0003806704, -0.002435244, 0.01042136, 
    0.0001675455, 0.001442469, 7.693568e-05, 4.05248e-08,
  -3.244084e-05, 0.02257203, 0.0002758593, 0.01127608, 0.09579278, 
    0.07413419, -0.003038991, 0.001565845, 0.01508333, 0.1991929, 0.04797422, 
    0.007365749, 0.01637242, 0.01522001, 0.02639354, 0.08844393, 0.1189441, 
    0.02433014, 0.06400003, 0.07769432, 0.1108494, 0.2063922, 0.1106144, 
    0.04505691, 0.06211125, 0.04204626, 0.004729497, 0.01771985, 0.001550447,
  0.01675142, 0.02042383, 0.1095007, 0.3043347, 0.01678361, 0.04999303, 
    0.1693811, 0.0002297109, 0.001136188, 0.06517798, 0.2274184, 0.02880623, 
    0.01927369, 0.05308807, 0.19316, 0.1892333, 0.2281996, 0.08741685, 
    0.05377369, 0.2945206, 0.1681519, 0.07941251, 0.3261544, 0.2348884, 
    0.1437089, 0.1597725, 0.1646479, 0.1050789, 0.1974837,
  0.1843323, 0.3532776, 0.3428235, 0.5528722, 0.3755283, 0.2559796, 
    0.1483205, 0.2265021, 0.06275325, 0.1640352, 0.1266124, 0.1394185, 
    0.05687797, 0.04395998, 0.2608696, 0.3235376, 0.2054801, 0.1006159, 
    0.08081259, 0.3918476, 0.1450959, 0.1465372, 0.2186162, 0.4969615, 
    0.2851985, 0.1470005, 0.1379983, 0.1209132, 0.180397,
  0.08166735, 0.4268506, 0.5354043, 0.565362, 0.6300862, 0.5480488, 
    0.6520243, 0.7643415, 0.6933846, 0.6866419, 0.7559795, 0.436496, 
    0.3212694, 0.16493, 0.3627166, 0.3567386, 0.5233384, 0.1731346, 
    0.3863843, 0.2733412, 0.8215871, 0.365727, 0.4822747, 0.3088825, 
    0.259667, 0.01843636, 0.06064121, 0.07551335, 0.122204,
  0.1944223, 0.185519, 0.3396705, 0.1319346, 0.4142314, 0.5724294, 0.7622488, 
    0.4532003, 0.4045819, 0.5261785, 0.4801393, 0.6427424, 0.754226, 
    0.6280092, 0.4614213, 0.2874015, 0.3651246, 0.2845102, 0.4328572, 
    0.5483965, 0.4453613, 0.6206664, 0.5530642, 0.3600232, 0.2766542, 
    0.3422059, 0.6158329, 0.175159, 0.3085575,
  0.4070839, 0.1373739, 0.3757792, 0.3517095, 0.4953892, 0.6660557, 
    0.6412817, 0.6215737, 0.5269803, 0.6137348, 0.6626629, 0.7157784, 
    0.769787, 0.7283004, 0.6032678, 0.6079236, 0.5815032, 0.5696045, 
    0.6527678, 0.5815802, 0.6168533, 0.4650547, 0.4654334, 0.2941182, 
    0.1082698, 0.04315129, 0.1560731, 0.3302009, 0.6402186,
  0.2197597, 0.2236073, 0.227455, 0.2313026, 0.2351503, 0.2389979, 0.2428456, 
    0.1988875, 0.2022018, 0.2055161, 0.2088304, 0.2121447, 0.215459, 
    0.2187734, 0.306343, 0.3060291, 0.3057151, 0.3054012, 0.3050872, 
    0.3047733, 0.3044593, 0.2534021, 0.2465541, 0.2397061, 0.2328581, 
    0.22601, 0.219162, 0.212314, 0.2166816,
  0.1146186, 0.1284907, 0.1177746, 0.126821, 0.0732173, 0.02580007, 
    0.04524288, 0.1401114, 0.2075213, 0.1565291, 0.1172496, 0.07857912, 
    0.09253548, -0.002782742, 0.07837933, 0.1353868, 0.07187439, 0.1235004, 
    0.08571154, 0.05348791, 0.09619158, 0.1608513, 0.2483869, 0.1408415, 
    0.08602706, 0.1343498, 0.07069183, 0.02757743, 0.04922357,
  0.1248149, 0.1000308, 0.1302564, 0.0770907, 0.03345878, 0.2130416, 
    0.08001107, 0.04425711, 0.0434425, 0.04876079, 0.04797063, 0.07267674, 
    0.03164532, 0.2060515, 0.3799014, 0.2734511, 0.3469403, 0.2911069, 
    0.2552262, 0.2581716, 0.2849813, 0.4203677, 0.5374444, 0.5523872, 
    0.1099074, 0.2977823, 0.3043162, 0.3026924, 0.2035836,
  0.3183392, 0.3385198, 0.4012362, 0.332545, 0.3661131, 0.3543535, 0.3356058, 
    0.1690702, 0.1676906, 0.2352895, 0.2310193, 0.2865351, 0.370885, 
    0.3123128, 0.1935507, 0.2641643, 0.2900154, 0.3321202, 0.2864821, 
    0.2134016, 0.2033444, 0.238044, 0.2715356, 0.2116082, 0.3002822, 
    0.442745, 0.4448765, 0.4424136, 0.4461473,
  0.2698845, 0.2362637, 0.2683093, 0.3093374, 0.3246185, 0.3135601, 
    0.3142661, 0.2761507, 0.2999685, 0.2646016, 0.2100688, 0.2256886, 
    0.1997449, 0.2039768, 0.1101647, 0.1502762, 0.1654688, 0.2231793, 
    0.1607261, 0.1332332, 0.151781, 0.2198963, 0.1717294, 0.08544292, 
    0.0396691, 0.107459, 0.2586707, 0.2586147, 0.2800333,
  0.06839982, 0.02697717, 0.01621218, 0.1600079, 0.1487772, 0.1157605, 
    0.1652032, 0.09912771, 0.08094915, 0.05878267, 0.08436481, 0.0249037, 
    0.01710806, 0.08103358, 0.2222221, 0.1172629, 0.09250128, 0.07983574, 
    0.1770351, 0.1923654, 0.1584867, 0.155929, 0.09783239, 0.09089383, 
    0.1033535, 0.1358691, 0.1920531, 0.1592273, 0.08149652,
  0.02382354, 0.01694392, 0.0152114, 0.04043527, 0.01779838, 0.01701917, 
    0.03727822, 0.009499709, 0.01271419, 0.01222864, 0.004131594, 
    0.0003065492, -0.0006508284, 0.004170104, 0.08578291, 0.01903891, 
    0.03742742, 0.1393752, 0.1029323, 0.0198944, 0.01601769, 0.006766508, 
    0.01450579, 0.006752243, 0.0002577662, 0.01762223, 0.03225233, 
    0.002811179, 0.003706026,
  0.01977022, 0.06681245, 0.00845428, 0.004131013, -0.002821814, 0.001305026, 
    0.001440244, 0.0009145332, 0.02867009, 0.003348247, 0.006019989, 
    7.042741e-05, 0.002123945, 0.004408603, 0.01090632, 0.001560779, 
    0.002879031, 0.001106794, 0.0003388744, 5.160435e-06, 7.235903e-05, 
    0.001847396, 0.02234893, 0.09806586, 0.02082673, 0.08572907, 
    6.423298e-05, 0.0009124114, 0.005458268,
  0.02887822, 0.004799722, 0.02263247, 0.06096717, 0.006443006, 0.0005551523, 
    0.002953272, 0.003472487, 0.001610404, 0.0008114229, 0.002295491, 
    0.000757163, 0.0005865198, 0.001187675, 0.0002436855, 0.0001487894, 
    3.445787e-05, 3.382552e-05, 2.82408e-05, 7.269898e-05, 0.003328037, 
    0.0142343, 0.05977743, 0.02251836, 0.02841539, 0.01215921, -0.0003932146, 
    0.0007892605, 0.009514472,
  0.02623323, 0.0004242743, 0.02525011, 0.05165325, 0.003045841, 
    0.0007616279, 0.01555501, 0.00263568, 0.04582117, 0.0874657, 0.007635543, 
    0.003856364, 0.0001500307, 0.0005671979, 0.000585736, 0.0008510026, 
    0.001794218, 0.0007804569, 0.0004365985, 0.0003761274, 0.003630399, 
    0.06796817, 0.0755235, 0.02904053, 0.008066191, 1.621263e-05, 
    0.002395238, 0.004699985, 0.001961594,
  6.357377e-10, 3.206079e-10, 3.39727e-09, 0.01196809, 0.09922738, 
    0.001195242, -0.002274492, 0.001230899, 0.006844297, 0.0005800684, 
    0.001704156, 0.0009636761, 0.00275066, 0.0003413826, 0.001939117, 
    0.002010345, 0.004112564, 0.004009036, 0.01170371, 0.01012834, 
    0.002636782, 0.0009733956, 0.1657404, 0.06266516, 0.002034357, 
    9.272827e-05, 0.002849119, -9.223128e-06, -2.058771e-07,
  9.170079e-09, 5.243048e-09, -6.978937e-09, -3.432919e-05, 0.0005133845, 
    0.00131592, 0.004804558, 0.0003374809, 0.03266509, 0.07342558, 
    0.004981223, 0.005869118, 0.0007511526, 0.0003583149, 0.0004955949, 
    0.0003266513, 0.002320687, 0.01830827, 0.008164681, 0.02899371, 
    0.003308816, 0.1112745, 0.0002078934, -0.001624754, 0.006820839, 
    9.296618e-05, 0.0008846314, 5.269532e-05, 4.336294e-08,
  -2.907999e-05, 0.01981209, 0.0001038486, 0.007738368, 0.08880068, 
    0.07103667, -0.0001505667, 0.0009848468, 0.01220657, 0.1564143, 
    0.03512747, 0.00415787, 0.0103475, 0.007897031, 0.01327891, 0.04886137, 
    0.06011336, 0.01212741, 0.04070367, 0.0445756, 0.09074248, 0.1748621, 
    0.0982812, 0.02357704, 0.04801749, 0.01525447, 0.001971321, 0.009545542, 
    0.0006970291,
  0.01095742, 0.01408159, 0.07743782, 0.2907879, 0.008771637, 0.03648115, 
    0.1575817, 0.001176026, 0.0007641072, 0.0579069, 0.1981697, 0.02115089, 
    0.0143286, 0.03789997, 0.1506018, 0.1382326, 0.1581036, 0.0546307, 
    0.03838543, 0.2842418, 0.1398666, 0.06691703, 0.2873552, 0.2074543, 
    0.1012121, 0.1068998, 0.1154609, 0.08042843, 0.148028,
  0.1289006, 0.3361846, 0.2931724, 0.4815644, 0.3214075, 0.1920601, 
    0.1179624, 0.2107194, 0.07014212, 0.1730934, 0.1005889, 0.1531154, 
    0.03569808, 0.03402314, 0.2344799, 0.2517578, 0.1564963, 0.06957145, 
    0.06595683, 0.368562, 0.1023868, 0.1029508, 0.192373, 0.4688374, 
    0.2141456, 0.1209113, 0.1104992, 0.08086465, 0.1266036,
  0.05347754, 0.4409231, 0.4677756, 0.5160118, 0.5946575, 0.4789514, 
    0.6199799, 0.7171469, 0.6860762, 0.6904086, 0.7399483, 0.4784839, 
    0.2745566, 0.1664428, 0.3046936, 0.2852509, 0.5030259, 0.1541535, 
    0.3609797, 0.2844015, 0.8442355, 0.3413652, 0.4457892, 0.3111065, 
    0.2341442, 0.01275596, 0.04798883, 0.06127756, 0.08728772,
  0.1612624, 0.1428543, 0.3282816, 0.08641474, 0.332321, 0.4403739, 
    0.6546895, 0.4158417, 0.4391582, 0.5279835, 0.6012326, 0.6087556, 
    0.8624506, 0.4680522, 0.4014866, 0.3587798, 0.3158477, 0.2317692, 
    0.3696155, 0.44975, 0.4169958, 0.672973, 0.6898192, 0.4139554, 0.4337173, 
    0.2688977, 0.6224231, 0.1040364, 0.2722846,
  0.3870505, 0.1150383, 0.385956, 0.4793539, 0.6762186, 0.7064464, 0.6371492, 
    0.6757209, 0.5982763, 0.6125499, 0.7465674, 0.7407264, 0.7177554, 
    0.6910635, 0.6080844, 0.6206171, 0.5752296, 0.5875629, 0.6311842, 
    0.6073447, 0.6799302, 0.4264209, 0.4840902, 0.4044915, 0.07721376, 
    0.02840046, 0.1506779, 0.2584805, 0.5794922,
  0.1388423, 0.1424826, 0.1461229, 0.1497632, 0.1534036, 0.1570439, 
    0.1606842, 0.1288067, 0.1318213, 0.1348359, 0.1378505, 0.1408652, 
    0.1438798, 0.1468944, 0.1935527, 0.1920101, 0.1904675, 0.188925, 
    0.1873824, 0.1858398, 0.1842972, 0.1575058, 0.1523935, 0.1472811, 
    0.1421688, 0.1370564, 0.1319441, 0.1268317, 0.13593,
  0.08461437, 0.09215746, 0.09054419, 0.1008403, 0.04521523, 0.02080829, 
    0.0287591, 0.09828699, 0.1488397, 0.1067655, 0.07730694, 0.05180975, 
    0.06167487, -0.002385885, 0.0592066, 0.09839453, 0.04637785, 0.08918928, 
    0.06016706, 0.03790886, 0.06301703, 0.116111, 0.2157486, 0.1047583, 
    0.05862179, 0.1018009, 0.04797516, 0.01695215, 0.02792582,
  0.1009953, 0.06937667, 0.08313335, 0.05264259, 0.02082388, 0.1798804, 
    0.06563154, 0.03407142, 0.03300519, 0.03631461, 0.03208151, 0.05176358, 
    0.02253566, 0.178511, 0.3091242, 0.2093628, 0.2746352, 0.2400895, 
    0.2008051, 0.1985098, 0.2138352, 0.3298542, 0.447781, 0.469368, 
    0.1380289, 0.2611684, 0.25346, 0.2311581, 0.155996,
  0.24624, 0.248758, 0.2962911, 0.2397178, 0.277449, 0.2791018, 0.2589393, 
    0.1138065, 0.1116376, 0.183291, 0.1777096, 0.2361067, 0.2902021, 
    0.2460363, 0.1385277, 0.1872662, 0.2318292, 0.2632401, 0.2175674, 
    0.1639773, 0.146729, 0.1610256, 0.1859753, 0.1317321, 0.2340461, 
    0.3774364, 0.3779345, 0.3401237, 0.3220482,
  0.2033948, 0.1731042, 0.195456, 0.2583814, 0.2670555, 0.2502501, 0.2441025, 
    0.1907856, 0.2201603, 0.1907911, 0.1538848, 0.1570179, 0.1404405, 
    0.1412772, 0.08276931, 0.09707692, 0.09639353, 0.1511018, 0.1060772, 
    0.09611107, 0.1048059, 0.1669528, 0.1236398, 0.06436223, 0.02868807, 
    0.08521228, 0.2056739, 0.1888673, 0.215721,
  0.04427152, 0.01489632, 0.009580793, 0.126097, 0.09806512, 0.07685585, 
    0.1116804, 0.06307843, 0.0484934, 0.03021092, 0.05239752, 0.01743621, 
    0.007505825, 0.05888617, 0.1948074, 0.07248136, 0.0624817, 0.04986759, 
    0.124185, 0.1249457, 0.09785379, 0.1039446, 0.06337099, 0.08177798, 
    0.09079047, 0.09103683, 0.1403784, 0.1040051, 0.04886856,
  0.01614586, 0.01002595, 0.01076806, 0.01610666, 0.007249649, 0.007055183, 
    0.02520779, 0.00649855, 0.008541154, 0.009811479, 0.00243611, 
    0.0001279066, -0.001394102, 0.002629699, 0.05714449, 0.01116001, 
    0.02252706, 0.09012507, 0.03617043, 0.007614377, 0.007589648, 
    0.004700769, 0.009254964, 0.004570132, 4.080325e-05, 0.007782765, 
    0.01440115, 0.001838687, 0.002367807,
  0.01186056, 0.04332205, 0.004107036, 0.001914286, -0.001906133, 
    0.0008073805, 0.0005580047, 0.0005757757, 0.01834844, 0.001432849, 
    0.004921415, 2.315719e-05, 0.001214523, 0.001217931, 0.004687066, 
    0.0005518707, 0.00117866, 0.0003403397, 0.0002130868, 2.791868e-06, 
    4.669583e-05, 0.001175403, 0.01200935, 0.0647916, 0.01249032, 0.06873951, 
    4.190267e-05, 0.000613008, 0.00311982,
  0.01827384, 0.0002082767, 0.01651542, 0.04858993, 0.003328769, 
    0.0002943988, 0.001174656, 0.001407013, 0.001010752, 0.0007682592, 
    0.0005970722, 0.0005058149, 8.526058e-05, 0.0004329936, 7.309971e-05, 
    6.205609e-05, 2.006848e-05, 1.828399e-05, 1.859603e-05, 4.681314e-05, 
    0.002155197, 0.008716208, 0.03701421, 0.01986589, 0.02668069, 
    0.009364333, -7.787883e-05, 0.0005160412, 0.006097923,
  0.01105662, 0.002274967, 0.01964918, 0.04351794, 0.001212068, 0.0004391043, 
    0.007405464, 0.0012601, 0.0359934, 0.0895395, 0.003711313, 0.002406828, 
    8.267301e-05, 0.0002876224, 0.0003846726, 0.000507076, 0.001075126, 
    0.0004564174, 0.0002937409, 0.0002182295, 0.001423728, 0.03338859, 
    0.03632516, 0.02523292, 0.006891882, 1.675718e-05, 0.0009041346, 
    0.002651174, 0.00104794,
  6.387736e-10, 3.169223e-10, 3.353526e-09, 0.01842306, 0.05454435, 
    0.0007865812, -0.002033475, 0.0008485912, 0.00289725, 0.0002984656, 
    0.0007855259, 0.0003886648, 0.001098714, 0.0001373709, 0.0006697893, 
    0.000966137, 0.001784091, 0.001304456, 0.004379684, 0.004479795, 
    0.001278055, 0.0006597938, 0.128982, 0.04945103, 0.0006903919, 
    5.094632e-05, 0.001958262, -7.157953e-06, -5.066197e-08,
  8.896377e-09, 5.140318e-09, -5.801272e-09, 1.559057e-05, 0.0002993756, 
    0.0009713719, 0.005962452, 0.0002416271, 0.03324633, 0.03770377, 
    0.001710377, 0.002578237, 0.0005138094, 0.0002324218, 0.0003194996, 
    0.0002096454, 0.000997014, 0.007999288, 0.004163412, 0.01101408, 
    0.001347534, 0.07362361, 0.0001379791, -0.001182726, 0.003651923, 
    6.1815e-05, 0.0006212111, 3.976332e-05, 4.339567e-08,
  -2.291166e-05, 0.01477411, 6.819289e-05, 0.005110168, 0.07515921, 
    0.06535993, 0.00670587, 0.0007315393, 0.01208804, 0.1134519, 0.02539393, 
    0.002989372, 0.006068999, 0.003911424, 0.006061377, 0.02646603, 
    0.0375958, 0.005216396, 0.02587125, 0.02447738, 0.07080712, 0.1405621, 
    0.08270616, 0.01695981, 0.028782, 0.005620804, 0.001137438, 0.006491886, 
    0.0003466991,
  0.008559017, 0.01093283, 0.0587602, 0.2682458, 0.005351979, 0.02667577, 
    0.1412199, 0.002568329, 0.0005933272, 0.05102696, 0.1692228, 0.01566383, 
    0.007852301, 0.02617971, 0.1073715, 0.08980642, 0.09970608, 0.03578865, 
    0.0236077, 0.2618805, 0.1158204, 0.05557529, 0.2355352, 0.1811764, 
    0.06489638, 0.05852288, 0.07041516, 0.0525681, 0.1009686,
  0.08119579, 0.2957265, 0.2466336, 0.3953352, 0.2571037, 0.1447462, 
    0.09032059, 0.1967542, 0.08836897, 0.1802414, 0.08267233, 0.1893987, 
    0.02495263, 0.02635475, 0.1874447, 0.1908432, 0.1145397, 0.05186329, 
    0.04764841, 0.3676628, 0.07682306, 0.07529259, 0.1640829, 0.4238921, 
    0.1756412, 0.1018377, 0.08082184, 0.05117659, 0.07674395,
  0.03052642, 0.4607167, 0.3973078, 0.4587223, 0.5299191, 0.3953719, 
    0.5705792, 0.6215802, 0.5962116, 0.6437774, 0.7071898, 0.5499614, 
    0.2602432, 0.1901468, 0.2489488, 0.2109352, 0.4829552, 0.1410232, 
    0.3116858, 0.2652649, 0.8443052, 0.3257589, 0.3158561, 0.3430129, 
    0.2181959, 0.008925777, 0.03625064, 0.04744774, 0.05601493,
  0.1249964, 0.09892668, 0.3094972, 0.06427006, 0.2608288, 0.3234767, 
    0.5298651, 0.4302699, 0.4793988, 0.5746469, 0.7202016, 0.5374492, 
    0.8408923, 0.3135099, 0.3590341, 0.360331, 0.2762237, 0.1769698, 
    0.3391041, 0.338382, 0.3337844, 0.6840536, 0.6590533, 0.5294213, 
    0.3449177, 0.1973104, 0.6081221, 0.07156266, 0.2242621,
  0.3706939, 0.1055124, 0.4504075, 0.5644404, 0.6889284, 0.6917335, 
    0.6012367, 0.6115847, 0.5658116, 0.5522311, 0.6869158, 0.6313943, 
    0.6455308, 0.5960052, 0.5497047, 0.5663873, 0.5094029, 0.5027248, 
    0.5257382, 0.5483465, 0.6094024, 0.355054, 0.4611598, 0.4993505, 
    0.05606395, 0.01537589, 0.1171229, 0.2106903, 0.50757,
  0.1068983, 0.1095244, 0.1121504, 0.1147765, 0.1174025, 0.1200286, 
    0.1226546, 0.08894544, 0.09012629, 0.09130715, 0.09248801, 0.09366886, 
    0.09484972, 0.09603058, 0.1247563, 0.1245304, 0.1243044, 0.1240784, 
    0.1238525, 0.1236265, 0.1234006, 0.1071914, 0.1036104, 0.1000295, 
    0.09644853, 0.09286759, 0.08928664, 0.08570569, 0.1047975,
  0.06781885, 0.06706832, 0.06922375, 0.0766318, 0.02685393, 0.01533536, 
    0.01377148, 0.07099236, 0.09859196, 0.08277003, 0.05052856, 0.03545106, 
    0.0441127, -0.001215999, 0.04544992, 0.07466652, 0.02969102, 0.07043893, 
    0.04789005, 0.0306829, 0.04511005, 0.08939567, 0.1933099, 0.08197133, 
    0.03978054, 0.08402179, 0.03847676, 0.01098308, 0.01518753,
  0.09437893, 0.05435951, 0.06330728, 0.03806744, 0.01600567, 0.1528724, 
    0.05400231, 0.02855963, 0.02627641, 0.03053001, 0.02507479, 0.0471129, 
    0.01635631, 0.1578218, 0.2504427, 0.1704572, 0.2152713, 0.1965088, 
    0.1560327, 0.1530483, 0.1650436, 0.2608011, 0.3574877, 0.3971983, 
    0.134196, 0.2074055, 0.2072593, 0.1829214, 0.1280096,
  0.1889821, 0.1965541, 0.2268727, 0.1880687, 0.2202416, 0.22992, 0.2043889, 
    0.08400235, 0.08487815, 0.1413837, 0.1424897, 0.187554, 0.2397018, 
    0.1909629, 0.1058691, 0.1437921, 0.1882583, 0.2179752, 0.1734667, 
    0.1270389, 0.1109722, 0.1130674, 0.1301722, 0.09017873, 0.192635, 
    0.3072181, 0.3084048, 0.2759837, 0.2506917,
  0.1600469, 0.1346749, 0.1497232, 0.2176537, 0.2212986, 0.2087663, 0.201379, 
    0.1429395, 0.1715786, 0.1437786, 0.1176624, 0.112935, 0.09511561, 
    0.1024725, 0.05414949, 0.06474618, 0.05983736, 0.1028864, 0.06998312, 
    0.06787151, 0.07088216, 0.1260681, 0.08919749, 0.0531977, 0.01821484, 
    0.06485487, 0.162634, 0.1483671, 0.1733997,
  0.03055969, 0.009927686, 0.004649966, 0.09253747, 0.05773507, 0.05273506, 
    0.07487261, 0.04259037, 0.03197759, 0.01645324, 0.02713827, 0.01343148, 
    0.003232556, 0.04258604, 0.1728879, 0.04387994, 0.03361332, 0.03216473, 
    0.07857814, 0.08306085, 0.06316721, 0.06882679, 0.04000195, 0.07552601, 
    0.07503088, 0.06010918, 0.09637601, 0.06846432, 0.03064363,
  0.01030097, 0.007186933, 0.007175323, 0.007036475, 0.003390611, 
    0.003584234, 0.01748107, 0.004936019, 0.006531569, 0.007447935, 
    0.001613749, 6.315735e-05, -0.0006959985, 0.001944017, 0.03411904, 
    0.007355911, 0.01419459, 0.05165527, 0.01568238, 0.004608043, 
    0.003601409, 0.003641114, 0.006794741, 0.003363339, -1.1243e-05, 
    0.004245403, 0.005862468, 0.001353247, 0.001705829,
  0.008367741, 0.03245163, 0.001433607, 0.001204541, -0.001218757, 
    0.0005960616, 0.0003711398, 0.0004171893, 0.01340571, 0.0008658117, 
    0.002306513, 5.983215e-06, 0.0008420155, 0.0004867684, 0.002358359, 
    0.0003408609, 0.0007276176, 0.0001850125, 0.0001553101, 1.758552e-06, 
    3.467707e-05, 0.0008553111, 0.007838369, 0.04917852, 0.008755966, 
    0.05452817, 3.160164e-05, 0.0004619691, 0.00213353,
  0.01333337, -0.001173137, 0.01712781, 0.05532675, 0.001675403, 
    0.0001992212, 0.0005593669, 0.0007572943, 0.0007516085, 0.0007453786, 
    0.0003045377, 0.0003792699, 0.0001097006, 0.0002625955, 7.796343e-05, 
    4.17884e-05, 1.383044e-05, 1.251812e-05, 1.415375e-05, 3.480088e-05, 
    0.001594777, 0.00622263, 0.02656145, 0.01911323, 0.02024108, 0.005880263, 
    2.066168e-05, 0.0003839585, 0.004480435,
  0.005087976, 0.006857761, 0.01194821, 0.03879691, 0.0007091252, 
    0.0003173912, 0.003781819, 0.0007326869, 0.0300687, 0.1053887, 
    0.001635374, 0.001721403, 5.885521e-05, 0.0001918263, 0.0002874524, 
    0.0003510374, 0.0007485985, 0.0003279694, 0.0002215837, 0.0001510679, 
    0.0008633666, 0.02181349, 0.02238841, 0.01543026, 0.0065207, 
    2.943181e-05, 0.0002987918, 0.00183422, 0.0007130549,
  6.546933e-10, 3.208254e-10, 3.264196e-09, 0.01954712, 0.03248666, 
    0.0005716453, -0.001480983, 0.0006523286, 0.001552797, 0.0002166095, 
    0.000460099, 0.0002168238, 0.0004596041, 0.0001281798, 0.0004500762, 
    0.0005860443, 0.0008579211, 0.0005529858, 0.001936152, 0.001928113, 
    0.0006467726, 0.000522966, 0.08195183, 0.03460731, 0.0002184967, 
    3.624584e-05, 0.001496291, -6.036331e-06, 1.206781e-08,
  8.838087e-09, 5.045771e-09, -4.063522e-09, 2.262681e-05, 0.0001988943, 
    0.0007750968, 0.005155456, 0.0001904872, 0.03188147, 0.02285378, 
    0.000939131, 0.001376696, 0.0004001043, 0.0001724064, 0.0002456689, 
    0.0001545569, 0.000710485, 0.003811003, 0.002502129, 0.006028164, 
    0.0006867645, 0.05249433, 0.000104011, -0.0007968471, 0.001960024, 
    4.681875e-05, 0.0004830242, 3.255531e-05, 4.308657e-08,
  -1.867683e-05, 0.01122605, 5.092595e-05, 0.003648916, 0.06437065, 
    0.05664359, 0.01088192, 0.0002447577, 0.01542915, 0.09142019, 0.01946761, 
    0.002407769, 0.003618139, 0.002077974, 0.002669727, 0.01340683, 
    0.02344206, 0.00275369, 0.01613629, 0.01515858, 0.05620989, 0.1108261, 
    0.07028487, 0.009757637, 0.01646812, 0.002747079, 0.0008312146, 
    0.005018502, 0.0002302993,
  0.008250573, 0.009044491, 0.04876592, 0.2500696, 0.003792148, 0.02092732, 
    0.133777, 0.004477574, 0.0003840476, 0.04992442, 0.1468535, 0.01255968, 
    0.003911532, 0.01944863, 0.08108856, 0.05924969, 0.06517062, 0.02414235, 
    0.01384116, 0.2448632, 0.1013977, 0.05170854, 0.1999248, 0.1569646, 
    0.04331892, 0.03534609, 0.04340848, 0.03411292, 0.07179525,
  0.05487958, 0.2867033, 0.2224255, 0.3502561, 0.2203029, 0.1179461, 
    0.07328204, 0.2035869, 0.1493099, 0.174034, 0.07671633, 0.2110758, 
    0.01964542, 0.02101177, 0.1495645, 0.1527796, 0.08672116, 0.04115367, 
    0.03590506, 0.3620184, 0.06260189, 0.06000391, 0.1436986, 0.3752517, 
    0.1532274, 0.08788028, 0.05914137, 0.03359388, 0.0495141,
  0.01997785, 0.5092049, 0.3440805, 0.4180834, 0.4869859, 0.3266208, 
    0.4999299, 0.4987333, 0.5243056, 0.5631057, 0.6244596, 0.6257026, 
    0.2845632, 0.289715, 0.2090321, 0.1735325, 0.4582275, 0.1485776, 0.29687, 
    0.2506572, 0.7897447, 0.3578326, 0.2619477, 0.3536008, 0.2088606, 
    0.007575982, 0.02935046, 0.03851498, 0.0382737,
  0.09987211, 0.07290423, 0.3193627, 0.05259838, 0.2204651, 0.2558531, 
    0.4667277, 0.4804469, 0.5535048, 0.6407728, 0.7366098, 0.4703106, 
    0.7392492, 0.2160285, 0.3076313, 0.3202086, 0.2661932, 0.1375283, 
    0.296437, 0.2350844, 0.2500409, 0.5894023, 0.463488, 0.5731692, 
    0.3092496, 0.1358172, 0.6077848, 0.05817036, 0.1873264,
  0.3237495, 0.1082196, 0.4518302, 0.5184644, 0.5931779, 0.5912575, 
    0.4740221, 0.4989811, 0.4676973, 0.3847705, 0.5255852, 0.4849478, 
    0.4822357, 0.4535227, 0.4109171, 0.3996141, 0.3517148, 0.3779091, 
    0.4128006, 0.4287177, 0.494171, 0.323704, 0.4191294, 0.6301517, 
    0.04926851, -0.009757184, 0.08763441, 0.2031645, 0.4461834,
  0.07674241, 0.07860156, 0.08046072, 0.08231987, 0.08417903, 0.08603818, 
    0.08789734, 0.07315909, 0.07404946, 0.07493982, 0.07583018, 0.07672054, 
    0.0776109, 0.07850127, 0.09775186, 0.09836602, 0.09898017, 0.09959433, 
    0.1002085, 0.1008226, 0.1014368, 0.08943492, 0.08607125, 0.08270758, 
    0.07934391, 0.07598023, 0.07261656, 0.06925289, 0.07525509,
  0.06298608, 0.05691301, 0.06131209, 0.07717377, 0.02421139, 0.01288224, 
    0.01071117, 0.0513334, 0.07735418, 0.08503043, 0.03960858, 0.02685577, 
    0.03522391, -0.0003264539, 0.04931224, 0.06398478, 0.02408099, 
    0.06036206, 0.04154532, 0.02708734, 0.03657857, 0.07589931, 0.1796639, 
    0.07000879, 0.03314331, 0.07509608, 0.03463275, 0.008714728, 0.01701164,
  0.08944723, 0.04869654, 0.06148015, 0.03286271, 0.01641401, 0.1420805, 
    0.04803126, 0.02436183, 0.02420384, 0.03217957, 0.026016, 0.04801219, 
    0.01031661, 0.1516435, 0.2191216, 0.1416121, 0.1817938, 0.1675168, 
    0.1331052, 0.13077, 0.1443812, 0.227842, 0.3173442, 0.3520614, 0.1319073, 
    0.1844665, 0.1825645, 0.1551737, 0.1148332,
  0.1599243, 0.173311, 0.1943768, 0.1643429, 0.1895636, 0.1981373, 0.1700947, 
    0.06910387, 0.07189347, 0.1166461, 0.1236738, 0.1600865, 0.2070978, 
    0.1587655, 0.08798613, 0.1217403, 0.1612822, 0.1878079, 0.1501958, 
    0.105462, 0.08959421, 0.09118524, 0.102213, 0.07341953, 0.1559036, 
    0.2573506, 0.2714084, 0.2390753, 0.2129272,
  0.1365836, 0.1156082, 0.1280543, 0.1667462, 0.1807948, 0.1706742, 
    0.1644632, 0.1160077, 0.1365421, 0.1155751, 0.0901473, 0.08907103, 
    0.07266884, 0.0780775, 0.04109372, 0.05092181, 0.0443731, 0.0719841, 
    0.04652427, 0.04938143, 0.05186573, 0.09672961, 0.06950966, 0.05409445, 
    0.01409558, 0.05160355, 0.1320976, 0.1256752, 0.1486487,
  0.02395922, 0.007925856, 0.002534769, 0.07134633, 0.0389872, 0.03886246, 
    0.05482458, 0.03311899, 0.02346515, 0.0117758, 0.01642733, 0.008884153, 
    0.001886934, 0.03258637, 0.1771589, 0.02612763, 0.02192899, 0.02405998, 
    0.05582446, 0.05971741, 0.04387022, 0.04834355, 0.02734996, 0.07451446, 
    0.06196548, 0.04259945, 0.07385412, 0.05011481, 0.02289991,
  0.006818268, 0.005820801, 0.00643782, 0.004423468, 0.00209278, 0.002379149, 
    0.0100331, 0.004154751, 0.005516865, 0.00662024, 0.001162897, 
    4.003219e-05, 0.004708822, 0.001621096, 0.02154372, 0.003682056, 
    0.009281944, 0.03205293, 0.01000405, 0.003560235, 0.002373256, 
    0.003057508, 0.005642797, 0.002892237, 0.0100522, 0.00285833, 
    0.003086736, 0.001126897, 0.001461668,
  0.006828115, 0.02480517, 0.0004614274, 0.0009445757, -0.001005346, 
    0.0004534765, 0.0002834828, 0.0003469134, 0.01102244, 0.000639838, 
    0.00131702, 5.821051e-06, 0.000675337, 0.000324026, 0.001593403, 
    0.0002660459, 0.0005602469, 0.0001366207, 0.0001268914, 1.483935e-06, 
    2.909415e-05, 0.0007067056, 0.006098886, 0.04111865, 0.0172463, 
    0.1098819, 2.684812e-05, 0.0003895465, 0.001724789,
  0.01089286, -0.001869039, 0.09256234, 0.191107, 0.001127976, 0.0001566114, 
    0.0003638073, 0.0005573084, 0.000622359, 0.0006124122, 0.0002276764, 
    0.0003130456, 9.996715e-05, 0.0001964496, 7.387314e-05, 3.412627e-05, 
    1.143295e-05, 1.011609e-05, 1.216487e-05, 2.962744e-05, 0.001331517, 
    0.005062417, 0.02152426, 0.05277992, 0.06264275, 0.009073108, 
    2.764452e-05, 0.0003209124, 0.00369194,
  0.003335272, 0.01295085, 0.00919114, 0.04454828, 0.0005434659, 
    0.0002565994, 0.002572852, 0.0005290723, 0.05668129, 0.1521932, 
    0.0009777243, 0.001396345, 4.721121e-05, 0.0001376088, 0.0002399201, 
    0.0002832334, 0.0005943499, 0.0002674702, 0.0001868454, 0.0001229502, 
    0.0006546876, 0.01678299, 0.01668819, 0.04693228, 0.04875861, 
    2.750041e-05, 0.0001625545, 0.001456656, 0.0005591787,
  6.914107e-10, 3.285214e-10, 3.025128e-09, 0.02643722, 0.02367212, 
    0.0004789266, -0.000873705, 0.0005568506, 0.0004506271, 0.0001788941, 
    0.0003432938, 0.0001563284, 0.0002450678, 0.0001195556, 0.0003819347, 
    0.0004441373, 0.000555128, 0.0003731927, 0.001213144, 0.001148088, 
    0.0004344675, 0.0002348514, 0.1153457, 0.03198906, 0.0001300501, 
    3.080647e-05, 0.001291966, -5.523569e-06, 4.289295e-08,
  8.910463e-09, 4.972332e-09, -2.631327e-09, 2.787722e-05, 0.0001479652, 
    0.0006610234, 0.00579881, 0.0001258209, 0.03526179, 0.01674386, 
    0.0007029538, 0.001044984, 0.0003496009, 0.0001443953, 0.0002096087, 
    0.0001276977, 0.0005891845, 0.002378242, 0.001997446, 0.004469979, 
    0.0004431653, 0.04344125, 8.700753e-05, -0.001107169, 0.001317861, 
    4.000215e-05, 0.000413544, 2.932824e-05, 4.310581e-08,
  -2.180679e-05, 0.009896423, -4.305858e-05, 0.003069621, 0.05867095, 
    0.0506773, 0.013424, 0.003519346, 0.03486427, 0.09126625, 0.01668287, 
    0.002111509, 0.002426771, 0.001457845, 0.001680818, 0.00845421, 
    0.01400048, 0.001955152, 0.01110636, 0.01031984, 0.04686815, 0.1015164, 
    0.07005238, 0.006401517, 0.01023549, 0.002040638, 0.00071583, 
    0.004249352, 0.0001918742,
  0.01375003, 0.007672369, 0.04366863, 0.243953, 0.003013764, 0.01754756, 
    0.1393087, 0.004312834, 0.0003136816, 0.05495225, 0.1580715, 0.01102558, 
    0.002882826, 0.01503551, 0.06678531, 0.04455733, 0.04684991, 0.01863032, 
    0.01000336, 0.2403723, 0.09655289, 0.05770707, 0.1994929, 0.1326907, 
    0.03366568, 0.02501314, 0.02850168, 0.02246423, 0.0593882,
  0.04225862, 0.2823487, 0.2178942, 0.3525177, 0.2011126, 0.1102139, 
    0.06833063, 0.2897291, 0.224319, 0.1911865, 0.08888017, 0.2421172, 
    0.01717811, 0.0190027, 0.1221795, 0.130416, 0.07169749, 0.03529044, 
    0.02914676, 0.3617601, 0.06949889, 0.05903922, 0.1791056, 0.3680743, 
    0.1476838, 0.07942633, 0.04856845, 0.02547696, 0.03601222,
  0.01535123, 0.6309308, 0.3512247, 0.4046215, 0.4978404, 0.3227935, 
    0.4809228, 0.4705833, 0.5063029, 0.5177954, 0.5925896, 0.668733, 
    0.3132243, 0.3571957, 0.1894073, 0.1574477, 0.4971336, 0.1706808, 
    0.3278597, 0.2964301, 0.7360989, 0.3437091, 0.2351655, 0.3438397, 
    0.2066546, 0.01125126, 0.02656389, 0.03422096, 0.03016223,
  0.08413054, 0.06074178, 0.3998737, 0.04626688, 0.2009985, 0.2117355, 
    0.4299994, 0.4914602, 0.6142505, 0.6261711, 0.7084478, 0.5391309, 
    0.636575, 0.1672683, 0.2684707, 0.3049728, 0.2902068, 0.1152548, 
    0.2664709, 0.2138121, 0.2116181, 0.5238129, 0.3692279, 0.5976136, 
    0.4011057, 0.1210185, 0.5426702, 0.05293959, 0.1647524,
  0.2961468, 0.120839, 0.4273916, 0.4435375, 0.50322, 0.5030227, 0.3562856, 
    0.3711035, 0.3763838, 0.3186927, 0.4227129, 0.3846642, 0.3544313, 
    0.3495493, 0.3309602, 0.3178602, 0.2630677, 0.2987846, 0.3151607, 
    0.3400934, 0.359919, 0.2849385, 0.4308001, 0.7030888, 0.04058774, 
    -0.007929325, 0.07648811, 0.2188214, 0.40944 ;

 lat = -89.5, -79.5, -69.5, -59.5, -49.5, -39.5, -29.5, -19.5, -9.5, 0.5, 
    10.5, 20.5, 30.5, 40.5, 50.5, 60.5, 70.5, 80.5 ;

 lat_bnds =
  -90, -89,
  -80, -79,
  -70, -69,
  -60, -59,
  -50, -49,
  -40, -39,
  -30, -29,
  -20, -19,
  -10, -9,
  0, 1,
  10, 11,
  20, 21,
  30, 31,
  40, 41,
  50, 51,
  60, 61,
  70, 71,
  80, 81 ;

 lon = 0.625, 13.125, 25.625, 38.125, 50.625, 63.125, 75.625, 88.125, 
    100.625, 113.125, 125.625, 138.125, 150.625, 163.125, 175.625, 188.125, 
    200.625, 213.125, 225.625, 238.125, 250.625, 263.125, 275.625, 288.125, 
    300.625, 313.125, 325.625, 338.125, 350.625 ;

 lon_bnds =
  0, 1.25,
  12.5, 13.75,
  25, 26.25,
  37.5, 38.75,
  50, 51.25,
  62.5, 63.75,
  75, 76.25,
  87.5, 88.75,
  100, 101.25,
  112.5, 113.75,
  125, 126.25,
  137.5, 138.75,
  150, 151.25,
  162.5, 163.75,
  175, 176.25,
  187.5, 188.75,
  200, 201.25,
  212.5, 213.75,
  225, 226.25,
  237.5, 238.75,
  250, 251.25,
  262.5, 263.75,
  275, 276.25,
  287.5, 288.75,
  300, 301.25,
  312.5, 313.75,
  325, 326.25,
  337.5, 338.75,
  350, 351.25 ;

 pfull = 0.0252729048206747, 0.0885404738757409, 0.213072411383256, 
    0.41190537807884, 0.671080828691593, 0.987471468515016, 1.36790961365676, 
    1.82562112064242, 2.38097588033244, 3.06218961364243, 3.90121721567151, 
    4.9296281825995, 6.18008131929323, 7.68875807563375, 9.49537809361575, 
    11.643153995098, 14.1786857151188, 17.1517875598959, 20.6152476986609, 
    24.6245259348741, 29.237386591333, 34.5134757786445, 40.5138467378254, 
    47.3004421634272, 54.9355325495126, 63.4811392623337, 72.9984371159701, 
    83.5471442618119, 95.1849171805989, 107.966767294215, 121.944503506415, 
    137.166169497631, 153.675572970355, 171.511834307961, 190.708985325578, 
    211.295632932361, 233.294677858721, 256.723099608772, 281.591803639405, 
    307.905555737256, 335.66293113824, 364.856338389786, 395.47216160598, 
    427.490864234311, 460.887168786725, 495.630391513078, 531.761718445649, 
    569.289185351388, 607.768705103107, 646.445374671436, 684.792067788697, 
    722.468679913451, 759.124006783627, 794.401045766566, 827.769968639223, 
    858.597822486016, 886.389109609622, 910.841030891388, 931.860653469283, 
    949.549679924174, 964.159924710431, 976.012345333387, 985.470174132691, 
    992.77226220014, 997.948601287575 ;

 time = 380.5, 410.5, 440.5, 471, 501.5, 532, 562.5, 593.5, 624, 654.5, 685, 
    715.5 ;

 time_bnds =
  365, 396,
  396, 425,
  425, 456,
  456, 486,
  486, 517,
  517, 547,
  547, 578,
  578, 609,
  609, 639,
  639, 670,
  670, 700,
  700, 731 ;
}
