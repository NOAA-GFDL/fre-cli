netcdf ocean_daily_cmip.19150101-19191231.tos {
dimensions:
	time = UNLIMITED ; // (1825 currently)
	nv = 2 ;
	yh = 576 ;
	xh = 720 ;
variables:
	double average_DT(time) ;
		average_DT:long_name = "Length of average period" ;
		average_DT:units = "days" ;
		average_DT:missing_value = 1.e+20 ;
		average_DT:_FillValue = 1.e+20 ;
	double average_T1(time) ;
		average_T1:long_name = "Start time for average period" ;
		average_T1:units = "days since 1850-01-01 00:00:00" ;
		average_T1:missing_value = 1.e+20 ;
		average_T1:_FillValue = 1.e+20 ;
	double average_T2(time) ;
		average_T2:long_name = "End time for average period" ;
		average_T2:units = "days since 1850-01-01 00:00:00" ;
		average_T2:missing_value = 1.e+20 ;
		average_T2:_FillValue = 1.e+20 ;
	double nv(nv) ;
		nv:long_name = "vertex number" ;
	double time(time) ;
		time:long_name = "time" ;
		time:units = "days since 1850-01-01 00:00:00" ;
		time:axis = "T" ;
		time:calendar_type = "NOLEAP" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bnds" ;
	double time_bnds(time, nv) ;
		time_bnds:long_name = "time axis boundaries" ;
		time_bnds:units = "days since 1850-01-01 00:00:00" ;
		time_bnds:missing_value = 1.e+20 ;
		time_bnds:_FillValue = 1.e+20 ;
	float tos(time, yh, xh) ;
		tos:long_name = "Sea Surface Temperature" ;
		tos:units = "degC" ;
		tos:missing_value = 1.e+20f ;
		tos:_FillValue = 1.e+20f ;
		tos:cell_methods = "area:mean yh:mean xh:mean time: mean" ;
		tos:cell_measures = "area: areacello" ;
		tos:time_avg_info = "average_T1,average_T2,average_DT" ;
		tos:standard_name = "sea_surface_temperature" ;
	double xh(xh) ;
		xh:long_name = "h point nominal longitude" ;
		xh:units = "degrees_east" ;
		xh:axis = "X" ;
	double yh(yh) ;
		yh:long_name = "h point nominal latitude" ;
		yh:units = "degrees_north" ;
		yh:axis = "Y" ;

// global attributes:
		:filename = "ocean_daily_cmip.19150101-19191231.tos.nc" ;
		:title = "ESM4_historical_D151" ;
		:associated_files = "areacello: 19150101.ocean_static.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:external_variables = "areacello" ;
data:

 nv = 1, 2 ;

 time = 23725.5, 23726.5, 23727.5, 23728.5, 23729.5, 23730.5, 23731.5, 
    23732.5, 23733.5, 23734.5, 23735.5, 23736.5, 23737.5, 23738.5, 23739.5, 
    23740.5, 23741.5, 23742.5, 23743.5, 23744.5, 23745.5, 23746.5, 23747.5, 
    23748.5, 23749.5, 23750.5, 23751.5, 23752.5, 23753.5, 23754.5, 23755.5, 
    23756.5, 23757.5, 23758.5, 23759.5, 23760.5, 23761.5, 23762.5, 23763.5, 
    23764.5, 23765.5, 23766.5, 23767.5, 23768.5, 23769.5, 23770.5, 23771.5, 
    23772.5, 23773.5, 23774.5, 23775.5, 23776.5, 23777.5, 23778.5, 23779.5, 
    23780.5, 23781.5, 23782.5, 23783.5, 23784.5, 23785.5, 23786.5, 23787.5, 
    23788.5, 23789.5, 23790.5, 23791.5, 23792.5, 23793.5, 23794.5, 23795.5, 
    23796.5, 23797.5, 23798.5, 23799.5, 23800.5, 23801.5, 23802.5, 23803.5, 
    23804.5, 23805.5, 23806.5, 23807.5, 23808.5, 23809.5, 23810.5, 23811.5, 
    23812.5, 23813.5, 23814.5, 23815.5, 23816.5, 23817.5, 23818.5, 23819.5, 
    23820.5, 23821.5, 23822.5, 23823.5, 23824.5, 23825.5, 23826.5, 23827.5, 
    23828.5, 23829.5, 23830.5, 23831.5, 23832.5, 23833.5, 23834.5, 23835.5, 
    23836.5, 23837.5, 23838.5, 23839.5, 23840.5, 23841.5, 23842.5, 23843.5, 
    23844.5, 23845.5, 23846.5, 23847.5, 23848.5, 23849.5, 23850.5, 23851.5, 
    23852.5, 23853.5, 23854.5, 23855.5, 23856.5, 23857.5, 23858.5, 23859.5, 
    23860.5, 23861.5, 23862.5, 23863.5, 23864.5, 23865.5, 23866.5, 23867.5, 
    23868.5, 23869.5, 23870.5, 23871.5, 23872.5, 23873.5, 23874.5, 23875.5, 
    23876.5, 23877.5, 23878.5, 23879.5, 23880.5, 23881.5, 23882.5, 23883.5, 
    23884.5, 23885.5, 23886.5, 23887.5, 23888.5, 23889.5, 23890.5, 23891.5, 
    23892.5, 23893.5, 23894.5, 23895.5, 23896.5, 23897.5, 23898.5, 23899.5, 
    23900.5, 23901.5, 23902.5, 23903.5, 23904.5, 23905.5, 23906.5, 23907.5, 
    23908.5, 23909.5, 23910.5, 23911.5, 23912.5, 23913.5, 23914.5, 23915.5, 
    23916.5, 23917.5, 23918.5, 23919.5, 23920.5, 23921.5, 23922.5, 23923.5, 
    23924.5, 23925.5, 23926.5, 23927.5, 23928.5, 23929.5, 23930.5, 23931.5, 
    23932.5, 23933.5, 23934.5, 23935.5, 23936.5, 23937.5, 23938.5, 23939.5, 
    23940.5, 23941.5, 23942.5, 23943.5, 23944.5, 23945.5, 23946.5, 23947.5, 
    23948.5, 23949.5, 23950.5, 23951.5, 23952.5, 23953.5, 23954.5, 23955.5, 
    23956.5, 23957.5, 23958.5, 23959.5, 23960.5, 23961.5, 23962.5, 23963.5, 
    23964.5, 23965.5, 23966.5, 23967.5, 23968.5, 23969.5, 23970.5, 23971.5, 
    23972.5, 23973.5, 23974.5, 23975.5, 23976.5, 23977.5, 23978.5, 23979.5, 
    23980.5, 23981.5, 23982.5, 23983.5, 23984.5, 23985.5, 23986.5, 23987.5, 
    23988.5, 23989.5, 23990.5, 23991.5, 23992.5, 23993.5, 23994.5, 23995.5, 
    23996.5, 23997.5, 23998.5, 23999.5, 24000.5, 24001.5, 24002.5, 24003.5, 
    24004.5, 24005.5, 24006.5, 24007.5, 24008.5, 24009.5, 24010.5, 24011.5, 
    24012.5, 24013.5, 24014.5, 24015.5, 24016.5, 24017.5, 24018.5, 24019.5, 
    24020.5, 24021.5, 24022.5, 24023.5, 24024.5, 24025.5, 24026.5, 24027.5, 
    24028.5, 24029.5, 24030.5, 24031.5, 24032.5, 24033.5, 24034.5, 24035.5, 
    24036.5, 24037.5, 24038.5, 24039.5, 24040.5, 24041.5, 24042.5, 24043.5, 
    24044.5, 24045.5, 24046.5, 24047.5, 24048.5, 24049.5, 24050.5, 24051.5, 
    24052.5, 24053.5, 24054.5, 24055.5, 24056.5, 24057.5, 24058.5, 24059.5, 
    24060.5, 24061.5, 24062.5, 24063.5, 24064.5, 24065.5, 24066.5, 24067.5, 
    24068.5, 24069.5, 24070.5, 24071.5, 24072.5, 24073.5, 24074.5, 24075.5, 
    24076.5, 24077.5, 24078.5, 24079.5, 24080.5, 24081.5, 24082.5, 24083.5, 
    24084.5, 24085.5, 24086.5, 24087.5, 24088.5, 24089.5, 24090.5, 24091.5, 
    24092.5, 24093.5, 24094.5, 24095.5, 24096.5, 24097.5, 24098.5, 24099.5, 
    24100.5, 24101.5, 24102.5, 24103.5, 24104.5, 24105.5, 24106.5, 24107.5, 
    24108.5, 24109.5, 24110.5, 24111.5, 24112.5, 24113.5, 24114.5, 24115.5, 
    24116.5, 24117.5, 24118.5, 24119.5, 24120.5, 24121.5, 24122.5, 24123.5, 
    24124.5, 24125.5, 24126.5, 24127.5, 24128.5, 24129.5, 24130.5, 24131.5, 
    24132.5, 24133.5, 24134.5, 24135.5, 24136.5, 24137.5, 24138.5, 24139.5, 
    24140.5, 24141.5, 24142.5, 24143.5, 24144.5, 24145.5, 24146.5, 24147.5, 
    24148.5, 24149.5, 24150.5, 24151.5, 24152.5, 24153.5, 24154.5, 24155.5, 
    24156.5, 24157.5, 24158.5, 24159.5, 24160.5, 24161.5, 24162.5, 24163.5, 
    24164.5, 24165.5, 24166.5, 24167.5, 24168.5, 24169.5, 24170.5, 24171.5, 
    24172.5, 24173.5, 24174.5, 24175.5, 24176.5, 24177.5, 24178.5, 24179.5, 
    24180.5, 24181.5, 24182.5, 24183.5, 24184.5, 24185.5, 24186.5, 24187.5, 
    24188.5, 24189.5, 24190.5, 24191.5, 24192.5, 24193.5, 24194.5, 24195.5, 
    24196.5, 24197.5, 24198.5, 24199.5, 24200.5, 24201.5, 24202.5, 24203.5, 
    24204.5, 24205.5, 24206.5, 24207.5, 24208.5, 24209.5, 24210.5, 24211.5, 
    24212.5, 24213.5, 24214.5, 24215.5, 24216.5, 24217.5, 24218.5, 24219.5, 
    24220.5, 24221.5, 24222.5, 24223.5, 24224.5, 24225.5, 24226.5, 24227.5, 
    24228.5, 24229.5, 24230.5, 24231.5, 24232.5, 24233.5, 24234.5, 24235.5, 
    24236.5, 24237.5, 24238.5, 24239.5, 24240.5, 24241.5, 24242.5, 24243.5, 
    24244.5, 24245.5, 24246.5, 24247.5, 24248.5, 24249.5, 24250.5, 24251.5, 
    24252.5, 24253.5, 24254.5, 24255.5, 24256.5, 24257.5, 24258.5, 24259.5, 
    24260.5, 24261.5, 24262.5, 24263.5, 24264.5, 24265.5, 24266.5, 24267.5, 
    24268.5, 24269.5, 24270.5, 24271.5, 24272.5, 24273.5, 24274.5, 24275.5, 
    24276.5, 24277.5, 24278.5, 24279.5, 24280.5, 24281.5, 24282.5, 24283.5, 
    24284.5, 24285.5, 24286.5, 24287.5, 24288.5, 24289.5, 24290.5, 24291.5, 
    24292.5, 24293.5, 24294.5, 24295.5, 24296.5, 24297.5, 24298.5, 24299.5, 
    24300.5, 24301.5, 24302.5, 24303.5, 24304.5, 24305.5, 24306.5, 24307.5, 
    24308.5, 24309.5, 24310.5, 24311.5, 24312.5, 24313.5, 24314.5, 24315.5, 
    24316.5, 24317.5, 24318.5, 24319.5, 24320.5, 24321.5, 24322.5, 24323.5, 
    24324.5, 24325.5, 24326.5, 24327.5, 24328.5, 24329.5, 24330.5, 24331.5, 
    24332.5, 24333.5, 24334.5, 24335.5, 24336.5, 24337.5, 24338.5, 24339.5, 
    24340.5, 24341.5, 24342.5, 24343.5, 24344.5, 24345.5, 24346.5, 24347.5, 
    24348.5, 24349.5, 24350.5, 24351.5, 24352.5, 24353.5, 24354.5, 24355.5, 
    24356.5, 24357.5, 24358.5, 24359.5, 24360.5, 24361.5, 24362.5, 24363.5, 
    24364.5, 24365.5, 24366.5, 24367.5, 24368.5, 24369.5, 24370.5, 24371.5, 
    24372.5, 24373.5, 24374.5, 24375.5, 24376.5, 24377.5, 24378.5, 24379.5, 
    24380.5, 24381.5, 24382.5, 24383.5, 24384.5, 24385.5, 24386.5, 24387.5, 
    24388.5, 24389.5, 24390.5, 24391.5, 24392.5, 24393.5, 24394.5, 24395.5, 
    24396.5, 24397.5, 24398.5, 24399.5, 24400.5, 24401.5, 24402.5, 24403.5, 
    24404.5, 24405.5, 24406.5, 24407.5, 24408.5, 24409.5, 24410.5, 24411.5, 
    24412.5, 24413.5, 24414.5, 24415.5, 24416.5, 24417.5, 24418.5, 24419.5, 
    24420.5, 24421.5, 24422.5, 24423.5, 24424.5, 24425.5, 24426.5, 24427.5, 
    24428.5, 24429.5, 24430.5, 24431.5, 24432.5, 24433.5, 24434.5, 24435.5, 
    24436.5, 24437.5, 24438.5, 24439.5, 24440.5, 24441.5, 24442.5, 24443.5, 
    24444.5, 24445.5, 24446.5, 24447.5, 24448.5, 24449.5, 24450.5, 24451.5, 
    24452.5, 24453.5, 24454.5, 24455.5, 24456.5, 24457.5, 24458.5, 24459.5, 
    24460.5, 24461.5, 24462.5, 24463.5, 24464.5, 24465.5, 24466.5, 24467.5, 
    24468.5, 24469.5, 24470.5, 24471.5, 24472.5, 24473.5, 24474.5, 24475.5, 
    24476.5, 24477.5, 24478.5, 24479.5, 24480.5, 24481.5, 24482.5, 24483.5, 
    24484.5, 24485.5, 24486.5, 24487.5, 24488.5, 24489.5, 24490.5, 24491.5, 
    24492.5, 24493.5, 24494.5, 24495.5, 24496.5, 24497.5, 24498.5, 24499.5, 
    24500.5, 24501.5, 24502.5, 24503.5, 24504.5, 24505.5, 24506.5, 24507.5, 
    24508.5, 24509.5, 24510.5, 24511.5, 24512.5, 24513.5, 24514.5, 24515.5, 
    24516.5, 24517.5, 24518.5, 24519.5, 24520.5, 24521.5, 24522.5, 24523.5, 
    24524.5, 24525.5, 24526.5, 24527.5, 24528.5, 24529.5, 24530.5, 24531.5, 
    24532.5, 24533.5, 24534.5, 24535.5, 24536.5, 24537.5, 24538.5, 24539.5, 
    24540.5, 24541.5, 24542.5, 24543.5, 24544.5, 24545.5, 24546.5, 24547.5, 
    24548.5, 24549.5, 24550.5, 24551.5, 24552.5, 24553.5, 24554.5, 24555.5, 
    24556.5, 24557.5, 24558.5, 24559.5, 24560.5, 24561.5, 24562.5, 24563.5, 
    24564.5, 24565.5, 24566.5, 24567.5, 24568.5, 24569.5, 24570.5, 24571.5, 
    24572.5, 24573.5, 24574.5, 24575.5, 24576.5, 24577.5, 24578.5, 24579.5, 
    24580.5, 24581.5, 24582.5, 24583.5, 24584.5, 24585.5, 24586.5, 24587.5, 
    24588.5, 24589.5, 24590.5, 24591.5, 24592.5, 24593.5, 24594.5, 24595.5, 
    24596.5, 24597.5, 24598.5, 24599.5, 24600.5, 24601.5, 24602.5, 24603.5, 
    24604.5, 24605.5, 24606.5, 24607.5, 24608.5, 24609.5, 24610.5, 24611.5, 
    24612.5, 24613.5, 24614.5, 24615.5, 24616.5, 24617.5, 24618.5, 24619.5, 
    24620.5, 24621.5, 24622.5, 24623.5, 24624.5, 24625.5, 24626.5, 24627.5, 
    24628.5, 24629.5, 24630.5, 24631.5, 24632.5, 24633.5, 24634.5, 24635.5, 
    24636.5, 24637.5, 24638.5, 24639.5, 24640.5, 24641.5, 24642.5, 24643.5, 
    24644.5, 24645.5, 24646.5, 24647.5, 24648.5, 24649.5, 24650.5, 24651.5, 
    24652.5, 24653.5, 24654.5, 24655.5, 24656.5, 24657.5, 24658.5, 24659.5, 
    24660.5, 24661.5, 24662.5, 24663.5, 24664.5, 24665.5, 24666.5, 24667.5, 
    24668.5, 24669.5, 24670.5, 24671.5, 24672.5, 24673.5, 24674.5, 24675.5, 
    24676.5, 24677.5, 24678.5, 24679.5, 24680.5, 24681.5, 24682.5, 24683.5, 
    24684.5, 24685.5, 24686.5, 24687.5, 24688.5, 24689.5, 24690.5, 24691.5, 
    24692.5, 24693.5, 24694.5, 24695.5, 24696.5, 24697.5, 24698.5, 24699.5, 
    24700.5, 24701.5, 24702.5, 24703.5, 24704.5, 24705.5, 24706.5, 24707.5, 
    24708.5, 24709.5, 24710.5, 24711.5, 24712.5, 24713.5, 24714.5, 24715.5, 
    24716.5, 24717.5, 24718.5, 24719.5, 24720.5, 24721.5, 24722.5, 24723.5, 
    24724.5, 24725.5, 24726.5, 24727.5, 24728.5, 24729.5, 24730.5, 24731.5, 
    24732.5, 24733.5, 24734.5, 24735.5, 24736.5, 24737.5, 24738.5, 24739.5, 
    24740.5, 24741.5, 24742.5, 24743.5, 24744.5, 24745.5, 24746.5, 24747.5, 
    24748.5, 24749.5, 24750.5, 24751.5, 24752.5, 24753.5, 24754.5, 24755.5, 
    24756.5, 24757.5, 24758.5, 24759.5, 24760.5, 24761.5, 24762.5, 24763.5, 
    24764.5, 24765.5, 24766.5, 24767.5, 24768.5, 24769.5, 24770.5, 24771.5, 
    24772.5, 24773.5, 24774.5, 24775.5, 24776.5, 24777.5, 24778.5, 24779.5, 
    24780.5, 24781.5, 24782.5, 24783.5, 24784.5, 24785.5, 24786.5, 24787.5, 
    24788.5, 24789.5, 24790.5, 24791.5, 24792.5, 24793.5, 24794.5, 24795.5, 
    24796.5, 24797.5, 24798.5, 24799.5, 24800.5, 24801.5, 24802.5, 24803.5, 
    24804.5, 24805.5, 24806.5, 24807.5, 24808.5, 24809.5, 24810.5, 24811.5, 
    24812.5, 24813.5, 24814.5, 24815.5, 24816.5, 24817.5, 24818.5, 24819.5, 
    24820.5, 24821.5, 24822.5, 24823.5, 24824.5, 24825.5, 24826.5, 24827.5, 
    24828.5, 24829.5, 24830.5, 24831.5, 24832.5, 24833.5, 24834.5, 24835.5, 
    24836.5, 24837.5, 24838.5, 24839.5, 24840.5, 24841.5, 24842.5, 24843.5, 
    24844.5, 24845.5, 24846.5, 24847.5, 24848.5, 24849.5, 24850.5, 24851.5, 
    24852.5, 24853.5, 24854.5, 24855.5, 24856.5, 24857.5, 24858.5, 24859.5, 
    24860.5, 24861.5, 24862.5, 24863.5, 24864.5, 24865.5, 24866.5, 24867.5, 
    24868.5, 24869.5, 24870.5, 24871.5, 24872.5, 24873.5, 24874.5, 24875.5, 
    24876.5, 24877.5, 24878.5, 24879.5, 24880.5, 24881.5, 24882.5, 24883.5, 
    24884.5, 24885.5, 24886.5, 24887.5, 24888.5, 24889.5, 24890.5, 24891.5, 
    24892.5, 24893.5, 24894.5, 24895.5, 24896.5, 24897.5, 24898.5, 24899.5, 
    24900.5, 24901.5, 24902.5, 24903.5, 24904.5, 24905.5, 24906.5, 24907.5, 
    24908.5, 24909.5, 24910.5, 24911.5, 24912.5, 24913.5, 24914.5, 24915.5, 
    24916.5, 24917.5, 24918.5, 24919.5, 24920.5, 24921.5, 24922.5, 24923.5, 
    24924.5, 24925.5, 24926.5, 24927.5, 24928.5, 24929.5, 24930.5, 24931.5, 
    24932.5, 24933.5, 24934.5, 24935.5, 24936.5, 24937.5, 24938.5, 24939.5, 
    24940.5, 24941.5, 24942.5, 24943.5, 24944.5, 24945.5, 24946.5, 24947.5, 
    24948.5, 24949.5, 24950.5, 24951.5, 24952.5, 24953.5, 24954.5, 24955.5, 
    24956.5, 24957.5, 24958.5, 24959.5, 24960.5, 24961.5, 24962.5, 24963.5, 
    24964.5, 24965.5, 24966.5, 24967.5, 24968.5, 24969.5, 24970.5, 24971.5, 
    24972.5, 24973.5, 24974.5, 24975.5, 24976.5, 24977.5, 24978.5, 24979.5, 
    24980.5, 24981.5, 24982.5, 24983.5, 24984.5, 24985.5, 24986.5, 24987.5, 
    24988.5, 24989.5, 24990.5, 24991.5, 24992.5, 24993.5, 24994.5, 24995.5, 
    24996.5, 24997.5, 24998.5, 24999.5, 25000.5, 25001.5, 25002.5, 25003.5, 
    25004.5, 25005.5, 25006.5, 25007.5, 25008.5, 25009.5, 25010.5, 25011.5, 
    25012.5, 25013.5, 25014.5, 25015.5, 25016.5, 25017.5, 25018.5, 25019.5, 
    25020.5, 25021.5, 25022.5, 25023.5, 25024.5, 25025.5, 25026.5, 25027.5, 
    25028.5, 25029.5, 25030.5, 25031.5, 25032.5, 25033.5, 25034.5, 25035.5, 
    25036.5, 25037.5, 25038.5, 25039.5, 25040.5, 25041.5, 25042.5, 25043.5, 
    25044.5, 25045.5, 25046.5, 25047.5, 25048.5, 25049.5, 25050.5, 25051.5, 
    25052.5, 25053.5, 25054.5, 25055.5, 25056.5, 25057.5, 25058.5, 25059.5, 
    25060.5, 25061.5, 25062.5, 25063.5, 25064.5, 25065.5, 25066.5, 25067.5, 
    25068.5, 25069.5, 25070.5, 25071.5, 25072.5, 25073.5, 25074.5, 25075.5, 
    25076.5, 25077.5, 25078.5, 25079.5, 25080.5, 25081.5, 25082.5, 25083.5, 
    25084.5, 25085.5, 25086.5, 25087.5, 25088.5, 25089.5, 25090.5, 25091.5, 
    25092.5, 25093.5, 25094.5, 25095.5, 25096.5, 25097.5, 25098.5, 25099.5, 
    25100.5, 25101.5, 25102.5, 25103.5, 25104.5, 25105.5, 25106.5, 25107.5, 
    25108.5, 25109.5, 25110.5, 25111.5, 25112.5, 25113.5, 25114.5, 25115.5, 
    25116.5, 25117.5, 25118.5, 25119.5, 25120.5, 25121.5, 25122.5, 25123.5, 
    25124.5, 25125.5, 25126.5, 25127.5, 25128.5, 25129.5, 25130.5, 25131.5, 
    25132.5, 25133.5, 25134.5, 25135.5, 25136.5, 25137.5, 25138.5, 25139.5, 
    25140.5, 25141.5, 25142.5, 25143.5, 25144.5, 25145.5, 25146.5, 25147.5, 
    25148.5, 25149.5, 25150.5, 25151.5, 25152.5, 25153.5, 25154.5, 25155.5, 
    25156.5, 25157.5, 25158.5, 25159.5, 25160.5, 25161.5, 25162.5, 25163.5, 
    25164.5, 25165.5, 25166.5, 25167.5, 25168.5, 25169.5, 25170.5, 25171.5, 
    25172.5, 25173.5, 25174.5, 25175.5, 25176.5, 25177.5, 25178.5, 25179.5, 
    25180.5, 25181.5, 25182.5, 25183.5, 25184.5, 25185.5, 25186.5, 25187.5, 
    25188.5, 25189.5, 25190.5, 25191.5, 25192.5, 25193.5, 25194.5, 25195.5, 
    25196.5, 25197.5, 25198.5, 25199.5, 25200.5, 25201.5, 25202.5, 25203.5, 
    25204.5, 25205.5, 25206.5, 25207.5, 25208.5, 25209.5, 25210.5, 25211.5, 
    25212.5, 25213.5, 25214.5, 25215.5, 25216.5, 25217.5, 25218.5, 25219.5, 
    25220.5, 25221.5, 25222.5, 25223.5, 25224.5, 25225.5, 25226.5, 25227.5, 
    25228.5, 25229.5, 25230.5, 25231.5, 25232.5, 25233.5, 25234.5, 25235.5, 
    25236.5, 25237.5, 25238.5, 25239.5, 25240.5, 25241.5, 25242.5, 25243.5, 
    25244.5, 25245.5, 25246.5, 25247.5, 25248.5, 25249.5, 25250.5, 25251.5, 
    25252.5, 25253.5, 25254.5, 25255.5, 25256.5, 25257.5, 25258.5, 25259.5, 
    25260.5, 25261.5, 25262.5, 25263.5, 25264.5, 25265.5, 25266.5, 25267.5, 
    25268.5, 25269.5, 25270.5, 25271.5, 25272.5, 25273.5, 25274.5, 25275.5, 
    25276.5, 25277.5, 25278.5, 25279.5, 25280.5, 25281.5, 25282.5, 25283.5, 
    25284.5, 25285.5, 25286.5, 25287.5, 25288.5, 25289.5, 25290.5, 25291.5, 
    25292.5, 25293.5, 25294.5, 25295.5, 25296.5, 25297.5, 25298.5, 25299.5, 
    25300.5, 25301.5, 25302.5, 25303.5, 25304.5, 25305.5, 25306.5, 25307.5, 
    25308.5, 25309.5, 25310.5, 25311.5, 25312.5, 25313.5, 25314.5, 25315.5, 
    25316.5, 25317.5, 25318.5, 25319.5, 25320.5, 25321.5, 25322.5, 25323.5, 
    25324.5, 25325.5, 25326.5, 25327.5, 25328.5, 25329.5, 25330.5, 25331.5, 
    25332.5, 25333.5, 25334.5, 25335.5, 25336.5, 25337.5, 25338.5, 25339.5, 
    25340.5, 25341.5, 25342.5, 25343.5, 25344.5, 25345.5, 25346.5, 25347.5, 
    25348.5, 25349.5, 25350.5, 25351.5, 25352.5, 25353.5, 25354.5, 25355.5, 
    25356.5, 25357.5, 25358.5, 25359.5, 25360.5, 25361.5, 25362.5, 25363.5, 
    25364.5, 25365.5, 25366.5, 25367.5, 25368.5, 25369.5, 25370.5, 25371.5, 
    25372.5, 25373.5, 25374.5, 25375.5, 25376.5, 25377.5, 25378.5, 25379.5, 
    25380.5, 25381.5, 25382.5, 25383.5, 25384.5, 25385.5, 25386.5, 25387.5, 
    25388.5, 25389.5, 25390.5, 25391.5, 25392.5, 25393.5, 25394.5, 25395.5, 
    25396.5, 25397.5, 25398.5, 25399.5, 25400.5, 25401.5, 25402.5, 25403.5, 
    25404.5, 25405.5, 25406.5, 25407.5, 25408.5, 25409.5, 25410.5, 25411.5, 
    25412.5, 25413.5, 25414.5, 25415.5, 25416.5, 25417.5, 25418.5, 25419.5, 
    25420.5, 25421.5, 25422.5, 25423.5, 25424.5, 25425.5, 25426.5, 25427.5, 
    25428.5, 25429.5, 25430.5, 25431.5, 25432.5, 25433.5, 25434.5, 25435.5, 
    25436.5, 25437.5, 25438.5, 25439.5, 25440.5, 25441.5, 25442.5, 25443.5, 
    25444.5, 25445.5, 25446.5, 25447.5, 25448.5, 25449.5, 25450.5, 25451.5, 
    25452.5, 25453.5, 25454.5, 25455.5, 25456.5, 25457.5, 25458.5, 25459.5, 
    25460.5, 25461.5, 25462.5, 25463.5, 25464.5, 25465.5, 25466.5, 25467.5, 
    25468.5, 25469.5, 25470.5, 25471.5, 25472.5, 25473.5, 25474.5, 25475.5, 
    25476.5, 25477.5, 25478.5, 25479.5, 25480.5, 25481.5, 25482.5, 25483.5, 
    25484.5, 25485.5, 25486.5, 25487.5, 25488.5, 25489.5, 25490.5, 25491.5, 
    25492.5, 25493.5, 25494.5, 25495.5, 25496.5, 25497.5, 25498.5, 25499.5, 
    25500.5, 25501.5, 25502.5, 25503.5, 25504.5, 25505.5, 25506.5, 25507.5, 
    25508.5, 25509.5, 25510.5, 25511.5, 25512.5, 25513.5, 25514.5, 25515.5, 
    25516.5, 25517.5, 25518.5, 25519.5, 25520.5, 25521.5, 25522.5, 25523.5, 
    25524.5, 25525.5, 25526.5, 25527.5, 25528.5, 25529.5, 25530.5, 25531.5, 
    25532.5, 25533.5, 25534.5, 25535.5, 25536.5, 25537.5, 25538.5, 25539.5, 
    25540.5, 25541.5, 25542.5, 25543.5, 25544.5, 25545.5, 25546.5, 25547.5, 
    25548.5, 25549.5 ;

 xh = -299.75, -299.25, -298.75, -298.25, -297.75, -297.25, -296.75, -296.25, 
    -295.75, -295.25, -294.75, -294.25, -293.75, -293.25, -292.75, -292.25, 
    -291.75, -291.25, -290.75, -290.25, -289.75, -289.25, -288.75, -288.25, 
    -287.75, -287.25, -286.75, -286.25, -285.75, -285.25, -284.75, -284.25, 
    -283.75, -283.25, -282.75, -282.25, -281.75, -281.25, -280.75, -280.25, 
    -279.75, -279.25, -278.75, -278.25, -277.75, -277.25, -276.75, -276.25, 
    -275.75, -275.25, -274.75, -274.25, -273.75, -273.25, -272.75, -272.25, 
    -271.75, -271.25, -270.75, -270.25, -269.75, -269.25, -268.75, -268.25, 
    -267.75, -267.25, -266.75, -266.25, -265.75, -265.25, -264.75, -264.25, 
    -263.75, -263.25, -262.75, -262.25, -261.75, -261.25, -260.75, -260.25, 
    -259.75, -259.25, -258.75, -258.25, -257.75, -257.25, -256.75, -256.25, 
    -255.75, -255.25, -254.75, -254.25, -253.75, -253.25, -252.75, -252.25, 
    -251.75, -251.25, -250.75, -250.25, -249.75, -249.25, -248.75, -248.25, 
    -247.75, -247.25, -246.75, -246.25, -245.75, -245.25, -244.75, -244.25, 
    -243.75, -243.25, -242.75, -242.25, -241.75, -241.25, -240.75, -240.25, 
    -239.75, -239.25, -238.75, -238.25, -237.75, -237.25, -236.75, -236.25, 
    -235.75, -235.25, -234.75, -234.25, -233.75, -233.25, -232.75, -232.25, 
    -231.75, -231.25, -230.75, -230.25, -229.75, -229.25, -228.75, -228.25, 
    -227.75, -227.25, -226.75, -226.25, -225.75, -225.25, -224.75, -224.25, 
    -223.75, -223.25, -222.75, -222.25, -221.75, -221.25, -220.75, -220.25, 
    -219.75, -219.25, -218.75, -218.25, -217.75, -217.25, -216.75, -216.25, 
    -215.75, -215.25, -214.75, -214.25, -213.75, -213.25, -212.75, -212.25, 
    -211.75, -211.25, -210.75, -210.25, -209.75, -209.25, -208.75, -208.25, 
    -207.75, -207.25, -206.75, -206.25, -205.75, -205.25, -204.75, -204.25, 
    -203.75, -203.25, -202.75, -202.25, -201.75, -201.25, -200.75, -200.25, 
    -199.75, -199.25, -198.75, -198.25, -197.75, -197.25, -196.75, -196.25, 
    -195.75, -195.25, -194.75, -194.25, -193.75, -193.25, -192.75, -192.25, 
    -191.75, -191.25, -190.75, -190.25, -189.75, -189.25, -188.75, -188.25, 
    -187.75, -187.25, -186.75, -186.25, -185.75, -185.25, -184.75, -184.25, 
    -183.75, -183.25, -182.75, -182.25, -181.75, -181.25, -180.75, -180.25, 
    -179.75, -179.25, -178.75, -178.25, -177.75, -177.25, -176.75, -176.25, 
    -175.75, -175.25, -174.75, -174.25, -173.75, -173.25, -172.75, -172.25, 
    -171.75, -171.25, -170.75, -170.25, -169.75, -169.25, -168.75, -168.25, 
    -167.75, -167.25, -166.75, -166.25, -165.75, -165.25, -164.75, -164.25, 
    -163.75, -163.25, -162.75, -162.25, -161.75, -161.25, -160.75, -160.25, 
    -159.75, -159.25, -158.75, -158.25, -157.75, -157.25, -156.75, -156.25, 
    -155.75, -155.25, -154.75, -154.25, -153.75, -153.25, -152.75, -152.25, 
    -151.75, -151.25, -150.75, -150.25, -149.75, -149.25, -148.75, -148.25, 
    -147.75, -147.25, -146.75, -146.25, -145.75, -145.25, -144.75, -144.25, 
    -143.75, -143.25, -142.75, -142.25, -141.75, -141.25, -140.75, -140.25, 
    -139.75, -139.25, -138.75, -138.25, -137.75, -137.25, -136.75, -136.25, 
    -135.75, -135.25, -134.75, -134.25, -133.75, -133.25, -132.75, -132.25, 
    -131.75, -131.25, -130.75, -130.25, -129.75, -129.25, -128.75, -128.25, 
    -127.75, -127.25, -126.75, -126.25, -125.75, -125.25, -124.75, -124.25, 
    -123.75, -123.25, -122.75, -122.25, -121.75, -121.25, -120.75, -120.25, 
    -119.75, -119.25, -118.75, -118.25, -117.75, -117.25, -116.75, -116.25, 
    -115.75, -115.25, -114.75, -114.25, -113.75, -113.25, -112.75, -112.25, 
    -111.75, -111.25, -110.75, -110.25, -109.75, -109.25, -108.75, -108.25, 
    -107.75, -107.25, -106.75, -106.25, -105.75, -105.25, -104.75, -104.25, 
    -103.75, -103.25, -102.75, -102.25, -101.75, -101.25, -100.75, -100.25, 
    -99.75, -99.25, -98.75, -98.25, -97.75, -97.25, -96.75, -96.25, -95.75, 
    -95.25, -94.75, -94.25, -93.75, -93.25, -92.75, -92.25, -91.75, -91.25, 
    -90.75, -90.25, -89.75, -89.25, -88.75, -88.25, -87.75, -87.25, -86.75, 
    -86.25, -85.75, -85.25, -84.75, -84.25, -83.75, -83.25, -82.75, -82.25, 
    -81.75, -81.25, -80.75, -80.25, -79.75, -79.25, -78.75, -78.25, -77.75, 
    -77.25, -76.75, -76.25, -75.75, -75.25, -74.75, -74.25, -73.75, -73.25, 
    -72.75, -72.25, -71.75, -71.25, -70.75, -70.25, -69.75, -69.25, -68.75, 
    -68.25, -67.75, -67.25, -66.75, -66.25, -65.75, -65.25, -64.75, -64.25, 
    -63.75, -63.25, -62.75, -62.25, -61.75, -61.25, -60.75, -60.25, -59.75, 
    -59.25, -58.75, -58.25, -57.75, -57.25, -56.75, -56.25, -55.75, -55.25, 
    -54.75, -54.25, -53.75, -53.25, -52.75, -52.25, -51.75, -51.25, -50.75, 
    -50.25, -49.75, -49.25, -48.75, -48.25, -47.75, -47.25, -46.75, -46.25, 
    -45.75, -45.25, -44.75, -44.25, -43.75, -43.25, -42.75, -42.25, -41.75, 
    -41.25, -40.75, -40.25, -39.75, -39.25, -38.75, -38.25, -37.75, -37.25, 
    -36.75, -36.25, -35.75, -35.25, -34.75, -34.25, -33.75, -33.25, -32.75, 
    -32.25, -31.75, -31.25, -30.75, -30.25, -29.75, -29.25, -28.75, -28.25, 
    -27.75, -27.25, -26.75, -26.25, -25.75, -25.25, -24.75, -24.25, -23.75, 
    -23.25, -22.75, -22.25, -21.75, -21.25, -20.75, -20.25, -19.75, -19.25, 
    -18.75, -18.25, -17.75, -17.25, -16.75, -16.25, -15.75, -15.25, -14.75, 
    -14.25, -13.75, -13.25, -12.75, -12.25, -11.75, -11.25, -10.75, -10.25, 
    -9.75, -9.25, -8.75, -8.25, -7.75, -7.25, -6.75, -6.25, -5.75, -5.25, 
    -4.75, -4.25, -3.75, -3.25, -2.75, -2.25, -1.75, -1.25, -0.75, -0.25, 
    0.25, 0.75, 1.25, 1.75, 2.25, 2.75, 3.25, 3.75, 4.25, 4.75, 5.25, 5.75, 
    6.25, 6.75, 7.25, 7.75, 8.25, 8.75, 9.25, 9.75, 10.25, 10.75, 11.25, 
    11.75, 12.25, 12.75, 13.25, 13.75, 14.25, 14.75, 15.25, 15.75, 16.25, 
    16.75, 17.25, 17.75, 18.25, 18.75, 19.25, 19.75, 20.25, 20.75, 21.25, 
    21.75, 22.25, 22.75, 23.25, 23.75, 24.25, 24.75, 25.25, 25.75, 26.25, 
    26.75, 27.25, 27.75, 28.25, 28.75, 29.25, 29.75, 30.25, 30.75, 31.25, 
    31.75, 32.25, 32.75, 33.25, 33.75, 34.25, 34.75, 35.25, 35.75, 36.25, 
    36.75, 37.25, 37.75, 38.25, 38.75, 39.25, 39.75, 40.25, 40.75, 41.25, 
    41.75, 42.25, 42.75, 43.25, 43.75, 44.25, 44.75, 45.25, 45.75, 46.25, 
    46.75, 47.25, 47.75, 48.25, 48.75, 49.25, 49.75, 50.25, 50.75, 51.25, 
    51.75, 52.25, 52.75, 53.25, 53.75, 54.25, 54.75, 55.25, 55.75, 56.25, 
    56.75, 57.25, 57.75, 58.25, 58.75, 59.25, 59.75 ;

 yh = -77.9079375348705, -77.7238126046114, -77.5396876743523, 
    -77.3555627440933, -77.1714378138342, -76.9873128835751, 
    -76.8031879533161, -76.619063023057, -76.4349380927979, 
    -76.2508131625389, -76.0666882322798, -75.8825633020207, 
    -75.6984383717617, -75.5143134415026, -75.3301885112435, 
    -75.1460635809845, -74.9619386507254, -74.7778137204664, 
    -74.5936887902073, -74.4095638599482, -74.2254389296892, 
    -74.0413139994301, -73.857189069171, -73.673064138912, -73.4889392086529, 
    -73.3048142783938, -73.1206893481348, -72.9365644178757, 
    -72.7524394876166, -72.5683145573576, -72.3841896270985, 
    -72.2000646968394, -72.0159397665804, -71.8318148363213, 
    -71.6476899060622, -71.4635649758032, -71.2794400455441, 
    -71.095315115285, -70.911190185026, -70.7270652547669, -70.5429403245078, 
    -70.3588153942488, -70.1746904639897, -69.9905655337306, 
    -69.8064406034716, -69.6223156732125, -69.4381907429535, 
    -69.2540658126944, -69.0699408824353, -68.8858159521763, 
    -68.7016910219172, -68.5175660916581, -68.3334411613991, -68.14931623114, 
    -67.9636445304209, -67.7752866505205, -67.5854009965385, 
    -67.3939772792524, -67.2010051944971, -67.0064744247379, 
    -66.8103746406885, -66.6126955029787, -66.4134266638701, 
    -66.2125577690213, -66.0100784593041, -65.8059783726705, 
    -65.6002471460721, -65.3928744174328, -65.1838498276744, 
    -64.9731630227985, -64.760803656022, -64.5467613899703, 
    -64.3310258989275, -64.1135868711439, -63.894434011203, 
    -63.6735570424482, -63.4509457094688, -63.2265897806486, 
    -63.0004790507758, -62.7726033437149, -62.5429525151436, 
    -62.3115164553525, -62.0782850921101, -61.8432483935938, 
    -61.6063963713863, -61.3677190835396, -61.1272066377062, 
    -60.884849194338, -60.6406369699546, -60.3945602404801, -60.14660934465, 
    -59.8967746874882, -59.6450467438542, -59.3914160620619, 
    -59.1358732675693, -58.8784090667402, -58.6190142506776, 
    -58.3576796991292, -58.0943963844658, -57.8291553757318, 
    -57.5619478427679, -57.2927650604075, -57.0215984127446, 
    -56.7484393974749, -56.4732796303085, -56.1961108494559, 
    -55.9169249201846, -55.6357138394475, -55.3524697405834, 
    -55.0671848980862, -54.7798517324457, -54.4904628150566, 
    -54.199010873197, -53.9054887950733, -53.6098896349336, 
    -53.3122066182453, -53.0124331469381, -52.7105628047106, 
    -52.4065893623985, -52.1005067834039, -51.7923092291839, 
    -51.4819910647963, -51.1695468645014, -50.8549714174182, 
    -50.5382597332318, -50.2194070479511, -49.8984088297146, 
    -49.5752607846407, -49.2499588627218, -48.9224992637582, 
    -48.5928784433296, -48.2610931188013, -47.9271402753627, 
    -47.5910171720938, -47.2527213480571, -46.9122506284122, 
    -46.5696031305474, -46.2247772702279, -45.8777717677532, 
    -45.5285856541224, -45.1772182772023, -44.8236693078935, 
    -44.4679387462917, -44.1100269278373, -43.7499345294513, 
    -43.3876625756504, -43.0232124446377, -42.6565858743633, 
    -42.2877849685499, -41.9168122026777, -41.5436704299229, 
    -41.1683628870455, -40.790893200218, -40.4112653907925, 
    -40.0294838809968, -39.6455534995561, -39.2594794872318, 
    -38.8712675022735, -38.4809236257751, -38.0884543669302, 
    -37.6938666681796, -37.2971679102448, -36.8983659170386, 
    -36.4974689604493, -36.0944857649878, -35.6894255122942, 
    -35.2822978454935, -34.8731128733961, -34.461881174534, 
    -34.0486138010269, -33.6333222822699, -33.2160186284369, 
    -32.7967153337909, -32.3754253797966, -31.952162238025, 
    -31.5269398728455, -31.0997727438981, -30.6706758083373, 
    -30.2396645228428, -29.8067548453888, -29.3722350905309, 
    -28.9369844818468, -28.5011135682704, -28.0647328987354, 
    -27.6279530221758, -27.1908844875253, -26.7536378437177, 
    -26.316323639687, -25.8790524243669, -25.4419347466912, 
    -25.0050811555939, -24.5686022000086, -24.1326084288694, 
    -23.6972103911098, -23.2625186356639, -22.8286437114655, 
    -22.3956961674483, -21.9637865525462, -21.533025415693, 
    -21.1035233058226, -20.6753907718688, -20.2487383627654, 
    -19.8236766274463, -19.4003161148452, -18.9787673738961, 
    -18.5591409535327, -18.1415474026888, -17.7260972702984, 
    -17.3129011052952, -16.9020694566131, -16.4937128731858, 
    -16.0879419039473, -15.6848670978313, -15.2845990037717, 
    -14.8872481707024, -14.492925147557, -14.1017404832696, 
    -13.7138047267738, -13.3292284270036, -12.9481221328927, 
    -12.5705963933751, -12.1967617573844, -11.8267287738547, 
    -11.4606079917196, -11.098509959913, -10.7405452273687, 
    -10.3868243430207, -10.0374578558026, -9.6925563146484, 
    -9.35223026849184, -9.01659026626678, -8.68574685690705, 
    -8.35981058934647, -8.03889201251887, -7.7231016753581, 
    -7.41255012679797, -7.10734791577232, -6.80760559121498, 
    -6.51343370205977, -6.22494279724053, -5.94224342569109, 
    -5.66544613634527, -5.39466147813692, -5.12999999999985, 
    -4.87179487179475, -4.6153846153845, -4.35897435897425, -4.102564102564, 
    -3.84615384615375, -3.5897435897435, -3.33333333333325, -3.076923076923, 
    -2.82051282051275, -2.5641025641025, -2.30769230769225, -2.051282051282, 
    -1.79487179487175, -1.5384615384615, -1.28205128205125, -1.025641025641, 
    -0.76923076923075, -0.5128205128205, -0.25641025641025, -0, 
    0.25641025641025, 0.5128205128205, 0.76923076923075, 1.025641025641, 
    1.28205128205125, 1.5384615384615, 1.79487179487175, 2.051282051282, 
    2.30769230769225, 2.5641025641025, 2.82051282051275, 3.076923076923, 
    3.33333333333325, 3.5897435897435, 3.84615384615375, 4.102564102564, 
    4.35897435897425, 4.6153846153845, 4.87179487179475, 5.12999999999985, 
    5.39466147813692, 5.66544613634527, 5.94224342569109, 6.22494279724053, 
    6.51343370205977, 6.80760559121498, 7.10734791577232, 7.41255012679797, 
    7.7231016753581, 8.03889201251887, 8.35981058934647, 8.68574685690705, 
    9.01659026626678, 9.35223026849184, 9.6925563146484, 10.0374578558026, 
    10.3868243430207, 10.7405452273687, 11.098509959913, 11.4606079917196, 
    11.8267287738547, 12.1967617573844, 12.5705963933751, 12.9481221328927, 
    13.3292284270036, 13.7138047267738, 14.1017404832696, 14.492925147557, 
    14.8872481707024, 15.2845990037717, 15.6848670978313, 16.0879419039473, 
    16.4937128731858, 16.9020694566131, 17.3129011052952, 17.7260972702984, 
    18.1415474026888, 18.5591409535327, 18.9787673738961, 19.4003161148452, 
    19.8236766274463, 20.2487383627654, 20.6753907718688, 21.1035233058226, 
    21.533025415693, 21.9637865525462, 22.3956961674483, 22.8286437114655, 
    23.2625186356639, 23.6972103911098, 24.1326084288694, 24.5686022000086, 
    25.0050811555939, 25.4419347466912, 25.8790524243669, 26.316323639687, 
    26.7536378437177, 27.1908844875253, 27.6279530221758, 28.0647328987354, 
    28.5011135682704, 28.9369844818468, 29.3722350905309, 29.8067548453888, 
    30.2396645228428, 30.6706758083373, 31.0997727438981, 31.5269398728455, 
    31.952162238025, 32.3754253797966, 32.7967153337909, 33.2160186284369, 
    33.6333222822699, 34.0486138010269, 34.461881174534, 34.8731128733961, 
    35.2822978454935, 35.6894255122942, 36.0944857649878, 36.4974689604493, 
    36.8983659170386, 37.2971679102448, 37.6938666681796, 38.0884543669302, 
    38.4809236257751, 38.8712675022735, 39.2594794872318, 39.6455534995561, 
    40.0294838809968, 40.4112653907925, 40.790893200218, 41.1683628870455, 
    41.5436704299229, 41.9168122026777, 42.2877849685499, 42.6565858743633, 
    43.0232124446377, 43.3876625756504, 43.7499345294513, 44.1100269278373, 
    44.4679387462917, 44.8236693078935, 45.1772182772023, 45.5285856541224, 
    45.8777717677532, 46.2247772702279, 46.5696031305474, 46.9122506284122, 
    47.2527213480571, 47.5910171720938, 47.9271402753627, 48.2610931188013, 
    48.5928784433296, 48.9224992637582, 49.2499588627218, 49.5752607846407, 
    49.8984088297146, 50.2194070479511, 50.5382597332318, 50.8549714174182, 
    51.1695468645014, 51.4819910647963, 51.7923092291839, 52.1005067834039, 
    52.4065893623985, 52.7105628047106, 53.0124331469381, 53.3122066182453, 
    53.6098896349336, 53.9054887950733, 54.199010873197, 54.4904628150566, 
    54.7798517324457, 55.0671848980862, 55.3524697405834, 55.6357138394475, 
    55.9169249201846, 56.1961108494559, 56.4732796303085, 56.7484393974749, 
    57.0215984127446, 57.2927650604075, 57.5619478427679, 57.8291553757318, 
    58.0943963844658, 58.3576796991292, 58.6190142506776, 58.8784090667402, 
    59.1358732675693, 59.3914160620619, 59.6450467438542, 59.8967746874882, 
    60.14660934465, 60.3945602404801, 60.6406369699546, 60.884849194338, 
    61.1272066377062, 61.3677190835396, 61.6063963713863, 61.8432483935938, 
    62.0782850921101, 62.3115164553525, 62.5429525151436, 62.7726033437149, 
    63.0004790507758, 63.2265897806486, 63.4509457094688, 63.6735570424482, 
    63.894434011203, 64.1135868711439, 64.3310258989275, 64.5467613899703, 
    64.760803656022, 64.9727930851569, 65.18399314351, 65.3951932018631, 
    65.6063932602162, 65.8175933185693, 66.0287933769224, 66.2399934352755, 
    66.4511934936286, 66.6623935519817, 66.8735936103349, 67.084793668688, 
    67.2959937270411, 67.5071937853942, 67.7183938437473, 67.9295939021004, 
    68.1407939604535, 68.3519940188066, 68.5631940771597, 68.7743941355128, 
    68.9855941938659, 69.196794252219, 69.4079943105721, 69.6191943689252, 
    69.8303944272783, 70.0415944856315, 70.2527945439845, 70.4639946023377, 
    70.6751946606908, 70.8863947190439, 71.097594777397, 71.3087948357501, 
    71.5199948941032, 71.7311949524563, 71.9423950108094, 72.1535950691625, 
    72.3647951275156, 72.5759951858687, 72.7871952442218, 72.9983953025749, 
    73.209595360928, 73.4207954192811, 73.6319954776342, 73.8431955359874, 
    74.0543955943405, 74.2655956526936, 74.4767957110467, 74.6879957693998, 
    74.8991958277529, 75.110395886106, 75.3215959444591, 75.5327960028122, 
    75.7439960611653, 75.9551961195184, 76.1663961778715, 76.3775962362246, 
    76.5887962945777, 76.7999963529308, 77.011196411284, 77.2223964696371, 
    77.4335965279902, 77.6447965863433, 77.8559966446964, 78.0671967030495, 
    78.2783967614026, 78.4895968197557, 78.7007968781088, 78.9119969364619, 
    79.123196994815, 79.3343970531681, 79.5455971115212, 79.7567971698743, 
    79.9679972282274, 80.1791972865805, 80.3903973449337, 80.6015974032868, 
    80.8127974616399, 81.023997519993, 81.2351975783461, 81.4463976366992, 
    81.6575976950523, 81.8687977534054, 82.0799978117585, 82.2911978701116, 
    82.5023979284647, 82.7135979868178, 82.9247980451709, 83.135998103524, 
    83.3471981618771, 83.5583982202303, 83.7695982785834, 83.9807983369365, 
    84.1919983952896, 84.4031984536427, 84.6143985119958, 84.8255985703489, 
    85.036798628702, 85.2479986870551, 85.4591987454082, 85.6703988037613, 
    85.8815988621144, 86.0927989204675, 86.3039989788206, 86.5151990371737, 
    86.7263990955269, 86.93759915388, 87.1487992122331, 87.3599992705862, 
    87.5711993289393, 87.7823993872924, 87.9935994456455, 88.2047995039986, 
    88.4159995623517, 88.6271996207048, 88.8383996790579, 89.049599737411, 
    89.2607997957641, 89.4719998541172, 89.6831999124703, 89.8943999708235 ;
}
