netcdf \00010101.atmos_daily.zg500.tile3 {
dimensions:
	time = UNLIMITED ; // (182 currently)
	phalf = 66 ;
	grid_xt = 15 ;
	grid_yt = 10 ;
	scalar_axis = 1 ;
	nv = 2 ;
	pfull = 65 ;
variables:
	double average_DT(time) ;
		average_DT:_FillValue = 1.e+20 ;
		average_DT:missing_value = 1.e+20 ;
		average_DT:units = "days" ;
		average_DT:long_name = "Length of average period" ;
	double average_T1(time) ;
		average_T1:_FillValue = 1.e+20 ;
		average_T1:missing_value = 1.e+20 ;
		average_T1:units = "days since 0001-01-01 00:00:00" ;
		average_T1:long_name = "Start time for average period" ;
	double average_T2(time) ;
		average_T2:_FillValue = 1.e+20 ;
		average_T2:missing_value = 1.e+20 ;
		average_T2:units = "days since 0001-01-01 00:00:00" ;
		average_T2:long_name = "End time for average period" ;
	float bk(phalf) ;
		bk:_FillValue = 1.e+20f ;
		bk:missing_value = 1.e+20f ;
		bk:long_name = "vertical coordinate sigma value" ;
		bk:cell_methods = "time: point" ;
	double grid_xt(grid_xt) ;
		grid_xt:units = "degrees_E" ;
		grid_xt:long_name = "T-cell longitude" ;
		grid_xt:axis = "X" ;
	double grid_yt(grid_yt) ;
		grid_yt:units = "degrees_N" ;
		grid_yt:long_name = "T-cell latitude" ;
		grid_yt:axis = "Y" ;
	float height10m(scalar_axis) ;
		height10m:_FillValue = 1.e+20f ;
		height10m:missing_value = 1.e+20f ;
		height10m:units = "m" ;
		height10m:long_name = "Height" ;
		height10m:cell_methods = "time: point" ;
		height10m:axis = "Z" ;
		height10m:positive = "up" ;
		height10m:standard_name = "height" ;
	float height2m(scalar_axis) ;
		height2m:_FillValue = 1.e+20f ;
		height2m:missing_value = 1.e+20f ;
		height2m:units = "m" ;
		height2m:long_name = "Height" ;
		height2m:cell_methods = "time: point" ;
		height2m:axis = "Z" ;
		height2m:positive = "up" ;
		height2m:standard_name = "height" ;
	double nv(nv) ;
		nv:long_name = "vertex number" ;
	double pfull(pfull) ;
		pfull:units = "mb" ;
		pfull:long_name = "ref full pressure level" ;
		pfull:axis = "Z" ;
		pfull:positive = "down" ;
	double phalf(phalf) ;
		phalf:units = "mb" ;
		phalf:long_name = "ref half pressure level" ;
		phalf:axis = "Z" ;
		phalf:positive = "down" ;
	float pk(phalf) ;
		pk:_FillValue = 1.e+20f ;
		pk:missing_value = 1.e+20f ;
		pk:units = "pascal" ;
		pk:long_name = "pressure part of the hybrid coordinate" ;
		pk:cell_methods = "time: point" ;
	double scalar_axis(scalar_axis) ;
		scalar_axis:long_name = "none" ;
	double time(time) ;
		time:units = "days since 0001-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "NOLEAP" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bnds" ;
	double time_bnds(time, nv) ;
		time_bnds:long_name = "time axis boundaries" ;
	float zg500(time, grid_yt, grid_xt) ;
		zg500:_FillValue = 1.e+20f ;
		zg500:missing_value = 1.e+20f ;
		zg500:units = "m" ;
		zg500:long_name = "Geopotential Height at 500 hPa" ;
		zg500:cell_methods = "time: mean" ;
		zg500:cell_measures = "area: area" ;
		zg500:time_avg_info = "average_T1,average_T2,average_DT" ;
		zg500:standard_name = "geopotential_height" ;

// global attributes:
		:title = "cm5_c96_am5f7c1r0_b06_piC_galb_noiceinit_alb" ;
		:associated_files = "area: 00010101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:history = "Wed Apr 30 14:48:00 2025: ncks -d grid_xt,0,14 -d grid_yt,0,9 -d time,0,181 /home/cew/Code/cmip7-sprint/testfiles/input/00010101.atmos_daily.tile3.nc -O /home/cew/Code/cmip7-sprint/testfiles/00010101.atmos_daily.tile3.nc\nFri Apr 25 14:15:06 2025: ncks -x -v sphum,psl 00010101.atmos_daily.tile3.nc -o reduce/00010101.atmos_daily.tile3.nc\nFri Apr 25 13:47:12 2025: ncks -d grid_xt,35,55 -d grid_yt,30,45 00010101.atmos_daily.tile3.nc var_select/00010101.atmos_daily.tile3.nc" ;
		:NCO = "netCDF Operators version 5.1.9 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 average_DT = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 average_T1 = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 
    18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 
    36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 
    54, 55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 
    72, 73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 
    90, 91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 
    106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 
    120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 
    134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 
    148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 
    162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 
    176, 177, 178, 179, 180, 181 ;

 average_T2 = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 
    19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 
    37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 
    55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 
    73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 
    91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 106, 
    107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 
    121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 
    135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 
    149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 
    163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 
    177, 178, 179, 180, 181, 182 ;

 bk = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.00193294, 0.00749994, 0.01640714, 0.02841953, 
    0.04334756, 0.06103661, 0.0813586, 0.1042054, 0.1294836, 0.1571101, 
    0.1870091, 0.2191095, 0.2533426, 0.2896406, 0.3279357, 0.3681587, 
    0.4102391, 0.454293, 0.5001689, 0.5468886, 0.5935643, 0.6397641, 
    0.6851825, 0.729505, 0.7723162, 0.8125153, 0.8492141, 0.8817441, 
    0.909788, 0.9332725, 0.9524949, 0.9678352, 0.9798011, 0.9889621, 0.99575, 1 ;

 grid_xt = 36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50 ;

 grid_yt = 31, 32, 33, 34, 35, 36, 37, 38, 39, 40 ;

 height10m = 10 ;

 height2m = 2 ;

 nv = 1, 2 ;

 pfull = 0.0252729048206747, 0.0885404738757409, 0.213072411383256, 
    0.41190537807884, 0.671080828691593, 0.987471468515016, 1.36790961365676, 
    1.82562112064242, 2.38097588033244, 3.06218961364243, 3.90121721567151, 
    4.9296281825995, 6.18008131929323, 7.68875807563375, 9.49537809361575, 
    11.643153995098, 14.1786857151188, 17.1517875598959, 20.6152476986609, 
    24.6245259348741, 29.237386591333, 34.5134757786445, 40.5138467378254, 
    47.3004421634272, 54.9355325495126, 63.4811392623337, 72.9984371159701, 
    83.5471442618119, 95.1849171805989, 107.966767294215, 121.944503506415, 
    137.166169497631, 153.675572970355, 171.511834307961, 190.708985325578, 
    211.295632932361, 233.294677858721, 256.723099608772, 281.591803639405, 
    307.905555737256, 335.66293113824, 364.856338389786, 395.47216160598, 
    427.490864234311, 460.887168786725, 495.630391513078, 531.761718445649, 
    569.289185351388, 607.768705103107, 646.445374671436, 684.792067788697, 
    722.468679913451, 759.124006783627, 794.401045766566, 827.769968639223, 
    858.597822486016, 886.389109609622, 910.841030891388, 931.860653469283, 
    949.549679924174, 964.159924710431, 976.012345333387, 985.470174132691, 
    992.77226220014, 997.948601287575 ;

 phalf = 0.01, 0.0513470268, 0.1404240036, 0.3072783852, 0.5379505539, 
    0.8245489502, 1.170559845, 1.5862843323, 2.0879000854, 2.700272522, 
    3.4550848389, 4.3841940308, 5.5185266113, 6.8925054932, 8.5440936279, 
    10.5147802734, 12.8495031738, 15.5965148926, 18.8071691895, 
    22.5356542969, 26.8386547852, 31.7749560547, 37.4049951172, 
    43.7903613281, 50.9932617188, 59.0759326172, 68.100078125, 78.1262353516, 
    89.2131933594, 101.4173632812, 114.7922466406, 129.3878501562, 
    145.2501478125, 162.4206823438, 180.9360560938, 200.8276451562, 
    222.1212074219, 244.8367185938, 268.9881007812, 294.5831945312, 
    321.6236510156, 350.1049399219, 380.0163883594, 411.3414303125, 
    444.0575547656, 478.1367280469, 513.5456339062, 550.403556875, 
    588.6019571094, 627.3470909766, 665.9273852344, 704.0097012891, 
    741.2475327734, 777.2856108203, 811.7659041211, 843.9830114648, 
    873.3803854492, 899.5263707422, 922.2501762402, 941.5376650684, 
    957.6070185254, 970.7426572876, 981.30107, 989.65107, 995.9000099865, 1000 ;

 pk = 1, 5.134703, 14.0424, 30.72784, 53.79506, 82.4549, 117.056, 158.6284, 
    208.79, 270.0273, 345.5085, 438.4194, 551.8527, 689.2505, 854.4094, 
    1051.478, 1284.95, 1559.651, 1880.717, 2253.565, 2683.865, 3177.496, 
    3740.5, 4379.036, 5099.326, 5907.593, 6810.008, 7812.624, 8921.319, 
    10141.74, 11285.93, 12188.79, 12884.3, 13400.12, 13758.85, 13979.1, 
    14076.26, 14063.13, 13950.46, 13747.31, 13461.45, 13099.54, 12667.38, 
    12170.08, 11612.19, 10997.8, 10330.65, 9611.055, 8843.304, 8045.85, 
    7236.312, 6424.557, 5606.509, 4778.059, 3944.972, 3146.775, 2416.634, 
    1778.226, 1246.215, 826.5195, 511.2139, 290.7407, 150, 68.893, 14.999, 0 ;

 scalar_axis = 0 ;

 time = 0.5, 1.5, 2.5, 3.5, 4.5, 5.5, 6.5, 7.5, 8.5, 9.5, 10.5, 11.5, 12.5, 
    13.5, 14.5, 15.5, 16.5, 17.5, 18.5, 19.5, 20.5, 21.5, 22.5, 23.5, 24.5, 
    25.5, 26.5, 27.5, 28.5, 29.5, 30.5, 31.5, 32.5, 33.5, 34.5, 35.5, 36.5, 
    37.5, 38.5, 39.5, 40.5, 41.5, 42.5, 43.5, 44.5, 45.5, 46.5, 47.5, 48.5, 
    49.5, 50.5, 51.5, 52.5, 53.5, 54.5, 55.5, 56.5, 57.5, 58.5, 59.5, 60.5, 
    61.5, 62.5, 63.5, 64.5, 65.5, 66.5, 67.5, 68.5, 69.5, 70.5, 71.5, 72.5, 
    73.5, 74.5, 75.5, 76.5, 77.5, 78.5, 79.5, 80.5, 81.5, 82.5, 83.5, 84.5, 
    85.5, 86.5, 87.5, 88.5, 89.5, 90.5, 91.5, 92.5, 93.5, 94.5, 95.5, 96.5, 
    97.5, 98.5, 99.5, 100.5, 101.5, 102.5, 103.5, 104.5, 105.5, 106.5, 107.5, 
    108.5, 109.5, 110.5, 111.5, 112.5, 113.5, 114.5, 115.5, 116.5, 117.5, 
    118.5, 119.5, 120.5, 121.5, 122.5, 123.5, 124.5, 125.5, 126.5, 127.5, 
    128.5, 129.5, 130.5, 131.5, 132.5, 133.5, 134.5, 135.5, 136.5, 137.5, 
    138.5, 139.5, 140.5, 141.5, 142.5, 143.5, 144.5, 145.5, 146.5, 147.5, 
    148.5, 149.5, 150.5, 151.5, 152.5, 153.5, 154.5, 155.5, 156.5, 157.5, 
    158.5, 159.5, 160.5, 161.5, 162.5, 163.5, 164.5, 165.5, 166.5, 167.5, 
    168.5, 169.5, 170.5, 171.5, 172.5, 173.5, 174.5, 175.5, 176.5, 177.5, 
    178.5, 179.5, 180.5, 181.5 ;

 time_bnds =
  0, 1,
  1, 2,
  2, 3,
  3, 4,
  4, 5,
  5, 6,
  6, 7,
  7, 8,
  8, 9,
  9, 10,
  10, 11,
  11, 12,
  12, 13,
  13, 14,
  14, 15,
  15, 16,
  16, 17,
  17, 18,
  18, 19,
  19, 20,
  20, 21,
  21, 22,
  22, 23,
  23, 24,
  24, 25,
  25, 26,
  26, 27,
  27, 28,
  28, 29,
  29, 30,
  30, 31,
  31, 32,
  32, 33,
  33, 34,
  34, 35,
  35, 36,
  36, 37,
  37, 38,
  38, 39,
  39, 40,
  40, 41,
  41, 42,
  42, 43,
  43, 44,
  44, 45,
  45, 46,
  46, 47,
  47, 48,
  48, 49,
  49, 50,
  50, 51,
  51, 52,
  52, 53,
  53, 54,
  54, 55,
  55, 56,
  56, 57,
  57, 58,
  58, 59,
  59, 60,
  60, 61,
  61, 62,
  62, 63,
  63, 64,
  64, 65,
  65, 66,
  66, 67,
  67, 68,
  68, 69,
  69, 70,
  70, 71,
  71, 72,
  72, 73,
  73, 74,
  74, 75,
  75, 76,
  76, 77,
  77, 78,
  78, 79,
  79, 80,
  80, 81,
  81, 82,
  82, 83,
  83, 84,
  84, 85,
  85, 86,
  86, 87,
  87, 88,
  88, 89,
  89, 90,
  90, 91,
  91, 92,
  92, 93,
  93, 94,
  94, 95,
  95, 96,
  96, 97,
  97, 98,
  98, 99,
  99, 100,
  100, 101,
  101, 102,
  102, 103,
  103, 104,
  104, 105,
  105, 106,
  106, 107,
  107, 108,
  108, 109,
  109, 110,
  110, 111,
  111, 112,
  112, 113,
  113, 114,
  114, 115,
  115, 116,
  116, 117,
  117, 118,
  118, 119,
  119, 120,
  120, 121,
  121, 122,
  122, 123,
  123, 124,
  124, 125,
  125, 126,
  126, 127,
  127, 128,
  128, 129,
  129, 130,
  130, 131,
  131, 132,
  132, 133,
  133, 134,
  134, 135,
  135, 136,
  136, 137,
  137, 138,
  138, 139,
  139, 140,
  140, 141,
  141, 142,
  142, 143,
  143, 144,
  144, 145,
  145, 146,
  146, 147,
  147, 148,
  148, 149,
  149, 150,
  150, 151,
  151, 152,
  152, 153,
  153, 154,
  154, 155,
  155, 156,
  156, 157,
  157, 158,
  158, 159,
  159, 160,
  160, 161,
  161, 162,
  162, 163,
  163, 164,
  164, 165,
  165, 166,
  166, 167,
  167, 168,
  168, 169,
  169, 170,
  170, 171,
  171, 172,
  172, 173,
  173, 174,
  174, 175,
  175, 176,
  176, 177,
  177, 178,
  178, 179,
  179, 180,
  180, 181,
  181, 182 ;

 zg500 =
  5016.91, 5014.094, 5010.697, 5008.675, 5005.066, 5001.233, 4997.681, 
    4997.488, 4998.486, 4999.898, 5006.186, 5016.654, 5028.275, 5041.976, 
    5056.665,
  5016.206, 5011.117, 5006.529, 5002.919, 4996.127, 4988.95, 4984.727, 
    4978.8, 4975.673, 4977.88, 4981.002, 4991.537, 5003.511, 5020.288, 
    5035.089,
  5016.883, 5010.208, 5003.837, 4998.53, 4988.037, 4981.21, 4965.73, 
    4963.812, 4955.026, 4951.932, 4954.414, 4963.894, 4978.147, 4996.36, 
    5016.882,
  5019.993, 5010.633, 5002.139, 4992.454, 4982.087, 4964.761, 4957.208, 
    4939.52, 4934.744, 4930.263, 4931.304, 4938.6, 4954.128, 4975.777, 
    4999.714,
  5027.089, 5014.977, 5003.647, 4991.393, 4977.18, 4962.76, 4944.542, 
    4934.722, 4922.415, 4912.895, 4915.585, 4921.293, 4937.432, 4958.279, 
    4986.216,
  5036.703, 5023.073, 5008.766, 4994.757, 4977.094, 4960.743, 4944.885, 
    4928.109, 4915.823, 4911.226, 4908.43, 4915.216, 4929.794, 4952.054, 
    4979.129,
  5050.585, 5036.109, 5020.361, 5004.626, 4986.902, 4969.612, 4952.109, 
    4939.521, 4926.878, 4918.279, 4916.16, 4921.684, 4934.462, 4954.931, 
    4979.824,
  5068.113, 5052.827, 5036.68, 5020.674, 5001.375, 4984.267, 4967.755, 
    4953.129, 4942.083, 4936.523, 4934.627, 4938.709, 4950.445, 4968.409, 
    4990.536,
  5088.918, 5073, 5057.331, 5041.878, 5025.108, 5008.585, 4991.771, 4979.022, 
    4968.467, 4961.878, 4960.02, 4963.774, 4973.188, 4988.205, 5007.15,
  5113.09, 5094.551, 5078.841, 5064.938, 5048.704, 5034.159, 5020.718, 
    5007.645, 4997.554, 4991.007, 4990.138, 4993.506, 5001.812, 5014.681, 
    5031.246,
  4964.104, 4953.202, 4942.328, 4937.605, 4933.519, 4931.811, 4931.452, 
    4935.724, 4944.386, 4964.776, 4998.107, 5044.174, 5090.215, 5135.171, 
    5176.324,
  4966.034, 4951.333, 4938.549, 4930.847, 4927.159, 4929.619, 4933.533, 
    4937.159, 4945.868, 4968.191, 4998.967, 5042.122, 5085.641, 5128.601, 
    5164.531,
  4970.005, 4951.095, 4936.989, 4927.704, 4922.616, 4929.083, 4930.461, 
    4941.885, 4951.889, 4969.895, 4999.942, 5038.318, 5080.658, 5116.869, 
    5155.171,
  4978.435, 4955.083, 4938.616, 4924.114, 4920.709, 4917.529, 4931.375, 
    4933.136, 4948.755, 4968.777, 4997.368, 5032.902, 5072.035, 5109.239, 
    5144.242,
  4992.264, 4966.385, 4946.037, 4929.044, 4919.9, 4920.502, 4922.087, 
    4935.609, 4950.612, 4964.158, 4992.821, 5024.387, 5061.628, 5092.841, 
    5127.604,
  5011.583, 4985.819, 4960.647, 4941.922, 4925.928, 4919.717, 4923.883, 
    4927.897, 4938.792, 4961.302, 4983.667, 5014.085, 5048.043, 5081.281, 
    5112.135,
  5033.725, 5009.99, 4984.143, 4961.83, 4944.298, 4932.804, 4927.23, 
    4934.295, 4944.453, 4957.689, 4977.411, 5004.117, 5033.513, 5063.951, 
    5094.141,
  5056.603, 5035.175, 5011.28, 4988.604, 4966.053, 4950.838, 4941.718, 
    4938.495, 4942.396, 4956.289, 4973.072, 4994.976, 5022.196, 5051.031, 
    5079.662,
  5078.818, 5060.523, 5038.536, 5018.315, 4997.584, 4979.124, 4963.716, 
    4958.027, 4958.125, 4963.239, 4974.663, 4992.668, 5015.098, 5040.763, 
    5066.865,
  5101.377, 5084.47, 5065.735, 5046.689, 5025.541, 5007.605, 4991.872, 
    4978.499, 4972.05, 4973.283, 4982.025, 4995.739, 5015.118, 5037.717, 
    5061.255,
  4965.508, 4944.197, 4923.596, 4913.562, 4908.782, 4912.33, 4917.467, 
    4931.029, 4942.224, 4958.373, 4980.552, 5007.733, 5046.747, 5098.196, 
    5150.428,
  4968.215, 4941.938, 4923.159, 4914.503, 4911.2, 4913.987, 4919.35, 
    4928.817, 4938.674, 4961.417, 4987.802, 5021.46, 5068.485, 5125.148, 
    5172.837,
  4969.981, 4944.117, 4926.535, 4920.448, 4917.022, 4921.107, 4923.172, 
    4933.15, 4948.123, 4969.45, 4999.146, 5038.013, 5092.211, 5145.019, 
    5193.941,
  4976.406, 4948.28, 4932.371, 4924.872, 4926.513, 4922.168, 4930.667, 
    4933.588, 4949.201, 4977.421, 5013.403, 5057.654, 5114.255, 5169.787, 
    5215.858,
  4984.003, 4956.619, 4939.627, 4932.04, 4932.65, 4933.905, 4934.578, 
    4944.057, 4968.045, 4989.234, 5030.337, 5078.192, 5137.853, 5186.284, 
    5232.592,
  4995.375, 4966.984, 4948.457, 4940.18, 4938.078, 4939.297, 4945.333, 
    4953.818, 4970.108, 5007.158, 5046.791, 5099.585, 5157.061, 5208.498, 
    5249.951,
  5009.294, 4981.26, 4960.468, 4950.643, 4947.007, 4949.817, 4954.341, 
    4971.055, 4996.217, 5026.274, 5067.87, 5121.389, 5174.519, 5222.446, 
    5264.068,
  5026.051, 4998.171, 4975.44, 4963.4, 4956.414, 4958.649, 4967.528, 4982.09, 
    5004.496, 5041.886, 5086.996, 5139.354, 5192.006, 5238.196, 5278.934,
  5042.819, 5017.827, 4994.755, 4980.218, 4973.251, 4973.764, 4981.654, 
    5001.744, 5028.396, 5062.28, 5105.221, 5156.646, 5205.822, 5249.696, 
    5288.351,
  5060.666, 5037.698, 5016.102, 5000.58, 4990.569, 4989.736, 4998.146, 
    5014.641, 5039.758, 5075.888, 5121.016, 5170.665, 5217.324, 5259.624, 
    5295.835,
  5053.167, 5034.066, 5017.181, 5009.562, 5002.811, 4998.091, 5001.071, 
    5014.876, 5030.06, 5042.117, 5058.143, 5081.231, 5112.723, 5143.874, 
    5176.053,
  5046.434, 5026.462, 5013.63, 5007.519, 5001.949, 5002.713, 5010.118, 
    5021.775, 5033.044, 5050.947, 5070.96, 5100.558, 5134.02, 5168.096, 
    5195.719,
  5037.902, 5019.254, 5009.813, 5007.252, 5004.847, 5011.55, 5015.954, 
    5033.975, 5048.736, 5062.968, 5087.302, 5120.816, 5155.892, 5185.038, 
    5211.652,
  5029.856, 5012.571, 5007.586, 5006.389, 5010.77, 5010.862, 5030.393, 
    5034.533, 5049.026, 5074.232, 5106.404, 5142.636, 5176.698, 5205.834, 
    5229.465,
  5021.601, 5009.204, 5006.215, 5008.668, 5012.692, 5023.625, 5030.677, 
    5049.259, 5072.149, 5090.511, 5129.556, 5163.571, 5197.002, 5219.525, 
    5241.724,
  5016.2, 5005.823, 5005.415, 5009.868, 5015.449, 5027.671, 5044.927, 
    5056.488, 5074.915, 5116.541, 5152.265, 5185.941, 5214.141, 5236.432, 
    5254.701,
  5011.336, 5005.644, 5008.044, 5013.108, 5021.902, 5035.701, 5051.525, 
    5076.204, 5108.191, 5142.523, 5175.876, 5206.787, 5229.801, 5249.096, 
    5267.563,
  5009.104, 5006.202, 5009.635, 5016.567, 5026.64, 5043.299, 5064.335, 
    5088.217, 5123.378, 5164.26, 5197.128, 5224.087, 5246.213, 5265.849, 
    5286.25,
  5008.533, 5010.289, 5016.562, 5024.48, 5038.133, 5055.566, 5079.263, 
    5115.556, 5155.787, 5188.698, 5217.145, 5241.263, 5263.069, 5284.27, 
    5308.26,
  5013.157, 5015.617, 5023.226, 5034.171, 5049.35, 5071.506, 5101.128, 
    5136.22, 5173.045, 5207.396, 5235.589, 5260.025, 5284.029, 5309.16, 
    5336.947,
  5179.965, 5178.492, 5168.348, 5155.463, 5139.925, 5127.719, 5122.734, 
    5124.899, 5132.28, 5143.704, 5167.479, 5200.307, 5236.374, 5269.353, 
    5303.806,
  5170.919, 5168.969, 5160.629, 5150.466, 5135.013, 5128.077, 5126.967, 
    5128.158, 5136.224, 5157.32, 5186.104, 5224.292, 5258.864, 5296.95, 
    5325.595,
  5161.221, 5159.636, 5152.942, 5144.043, 5133.692, 5131.419, 5129.407, 
    5139.097, 5153.175, 5172.683, 5207.512, 5244.565, 5280.532, 5312.75, 
    5343.656,
  5150.37, 5148.356, 5143.239, 5136.951, 5133.415, 5130.764, 5138.978, 
    5140.056, 5155.931, 5189.007, 5226.767, 5263.86, 5300.461, 5333.773, 
    5363.617,
  5138.666, 5137.86, 5134.233, 5132.593, 5131.871, 5139.424, 5140.556, 
    5156.744, 5182.905, 5205.73, 5246.537, 5281.227, 5317.599, 5346.397, 
    5376.268,
  5125.947, 5125.923, 5123.713, 5126.611, 5131.405, 5140.32, 5153.741, 
    5163.222, 5184.769, 5227.385, 5263.923, 5299.275, 5332.004, 5361.696, 
    5388.354,
  5114.322, 5116.938, 5117.978, 5124.765, 5134.271, 5147.301, 5159.118, 
    5182.841, 5215.464, 5248.092, 5282.717, 5315.061, 5344.748, 5371.259, 
    5395.952,
  5104.532, 5108.853, 5112.482, 5123.481, 5136.456, 5152.312, 5169.974, 
    5191.905, 5223.057, 5262.836, 5296.661, 5327.369, 5355.673, 5381.037, 
    5404.72,
  5096.738, 5104.775, 5114.322, 5128.335, 5144.333, 5161.17, 5181.11, 
    5212.636, 5249.272, 5281.499, 5310.74, 5338.636, 5363.901, 5387.605, 
    5410.075,
  5091.924, 5102.128, 5115.279, 5132.816, 5151.35, 5172.238, 5196.762, 
    5226.804, 5260.731, 5293.474, 5322.507, 5347.812, 5371.587, 5394.847, 
    5417.328,
  5233.297, 5242.573, 5250.869, 5257.121, 5256.113, 5248.693, 5250.685, 
    5268.249, 5292.704, 5319.059, 5345.813, 5369.455, 5389.122, 5402.452, 
    5411.551,
  5225.122, 5234.228, 5244.375, 5252.137, 5251.38, 5246.3, 5250.322, 
    5267.345, 5293.993, 5328.791, 5358.56, 5385.494, 5404.92, 5420.778, 
    5428.75,
  5217.466, 5227.001, 5239.259, 5248.47, 5249.897, 5245.475, 5249.286, 
    5273.033, 5305.125, 5337.419, 5370.144, 5398.114, 5420.39, 5434.864, 
    5444.518,
  5210.694, 5220.647, 5233.517, 5243.054, 5247.887, 5241.056, 5251.527, 
    5265.611, 5300.106, 5342.21, 5379.124, 5408.378, 5432.768, 5448.653, 
    5459.307,
  5203.421, 5214.807, 5227.973, 5239.609, 5242.719, 5245.677, 5244.671, 
    5274.482, 5312.913, 5346.203, 5386.003, 5417.435, 5443.11, 5459.305, 
    5470.628,
  5195.087, 5208.192, 5220.829, 5232.602, 5236.883, 5238.519, 5248.397, 
    5265.25, 5300.565, 5352.047, 5390.25, 5425.393, 5450.791, 5469.892, 
    5480.67,
  5186.447, 5201.258, 5214.364, 5226.139, 5232.044, 5236.194, 5242.479, 
    5269.534, 5313.333, 5354.024, 5395.351, 5430.576, 5457.487, 5476.848, 
    5487.834,
  5178.374, 5194.044, 5205.89, 5217.756, 5223.616, 5230.45, 5239.363, 
    5258.304, 5300.479, 5353.015, 5396.491, 5433.473, 5461.814, 5481.93, 
    5493.266,
  5171.337, 5187.92, 5199.991, 5212.035, 5219.223, 5225.357, 5236.141, 
    5260.119, 5306.741, 5354.842, 5396.884, 5435.836, 5463.626, 5484.258, 
    5494.451,
  5165.549, 5181.38, 5192.499, 5204.688, 5212.793, 5220.438, 5232.735, 
    5251.987, 5297.253, 5350.659, 5396.982, 5436.067, 5464.341, 5484.622, 
    5494.305,
  5304.342, 5295.548, 5295.882, 5302.979, 5309.552, 5325.196, 5342.271, 
    5358.164, 5369.121, 5373.128, 5373.361, 5371.386, 5365.783, 5357.827, 
    5348.687,
  5302.169, 5294.971, 5295.469, 5302.486, 5307.183, 5324.304, 5345.019, 
    5361.892, 5373.83, 5384.091, 5386.797, 5387.224, 5382.823, 5378.602, 
    5371.389,
  5296.761, 5292.204, 5293.819, 5301.368, 5306.707, 5324.667, 5344.724, 
    5368.631, 5385.419, 5394, 5398.711, 5400.163, 5398.537, 5394.422, 5388.685,
  5286.5, 5286.844, 5289.351, 5296.836, 5305.753, 5317.615, 5348.11, 
    5365.288, 5386.204, 5400.51, 5409.357, 5410.796, 5411.138, 5407.304, 
    5403.961,
  5273.489, 5278.876, 5283.599, 5294.308, 5301.725, 5319.451, 5341.687, 
    5372.021, 5395.508, 5407.386, 5418.732, 5422.645, 5424.335, 5420.768, 
    5417.125,
  5254.693, 5265.227, 5273.691, 5286.361, 5295.998, 5309.705, 5342.491, 
    5365.466, 5390.757, 5413.823, 5426.14, 5434.199, 5437.083, 5435.911, 
    5431.647,
  5234.334, 5249.127, 5263.425, 5278.929, 5292.087, 5305.242, 5333.7, 
    5368.495, 5397.61, 5416.967, 5433.541, 5444.533, 5450.178, 5450.412, 
    5445.873,
  5216.446, 5233.226, 5249.754, 5268.624, 5283.405, 5297.624, 5326.244, 
    5357.964, 5388.279, 5416.993, 5437.504, 5451.803, 5460.655, 5463.021, 
    5460.061,
  5202.231, 5219.583, 5240.299, 5261.27, 5279.199, 5292.269, 5317.057, 
    5353.853, 5387.07, 5414.876, 5437.829, 5455.863, 5467.656, 5472.538, 
    5470.844,
  5192.268, 5208.158, 5228.499, 5250.641, 5270.745, 5286.146, 5308.207, 
    5340.504, 5373.452, 5406.508, 5434.354, 5455.415, 5470.299, 5477.965, 
    5478.793,
  5305.358, 5300.871, 5294.144, 5289.099, 5293.458, 5295.626, 5292.379, 
    5287.74, 5284.036, 5281.228, 5281.517, 5284.889, 5289.504, 5294.116, 
    5298.63,
  5286.63, 5287.205, 5287.807, 5285.776, 5291.618, 5298.938, 5302.233, 
    5300.458, 5296.928, 5297.403, 5298.584, 5302.704, 5306.599, 5312.124, 
    5317.446,
  5263.654, 5270.401, 5278.108, 5280.729, 5289.494, 5301.805, 5307.004, 
    5311.782, 5312.261, 5312.123, 5314.466, 5318.479, 5324.295, 5329.813, 
    5335.516,
  5242.844, 5254.558, 5267.319, 5273.342, 5284.738, 5298.534, 5312.775, 
    5315.891, 5319.169, 5322.978, 5327.643, 5332.045, 5338.673, 5344.876, 
    5352.235,
  5233.162, 5245.374, 5260.588, 5269.976, 5279.553, 5299.707, 5311.638, 
    5323.576, 5329.331, 5331.127, 5337.231, 5342.729, 5350.661, 5357.801, 
    5365.603,
  5226.101, 5239.761, 5254.969, 5265.957, 5274.018, 5293.788, 5313.596, 
    5324.348, 5330.586, 5338.459, 5344.56, 5352.694, 5361.12, 5370.716, 
    5378.206,
  5223.362, 5237.423, 5252.211, 5263.891, 5272.334, 5290.913, 5310.813, 
    5327.636, 5337.453, 5344.323, 5352.071, 5361.927, 5372.212, 5382.049, 
    5389.128,
  5227.12, 5233.905, 5246.946, 5259.743, 5267.698, 5285.156, 5308.469, 
    5325.439, 5337.292, 5348.973, 5358.99, 5370.699, 5382.082, 5392.369, 
    5399.688,
  5235.562, 5233.456, 5241.332, 5255.797, 5266.669, 5281.458, 5304.097, 
    5325.004, 5340.599, 5352.986, 5365.465, 5379.081, 5391.451, 5401.956, 
    5409.507,
  5236.447, 5235.798, 5235.167, 5246.569, 5260.008, 5274.4, 5297.864, 
    5320.193, 5337.777, 5354.221, 5370.062, 5385.445, 5399.146, 5411.028, 
    5419.344,
  5189.159, 5203.968, 5215.478, 5223.44, 5229.025, 5236.602, 5246.618, 
    5260.452, 5272.687, 5280.221, 5285.386, 5288.685, 5289.299, 5289.144, 
    5288.142,
  5178.89, 5194.617, 5210.849, 5222.227, 5228.845, 5236.762, 5248.552, 
    5261.236, 5274.012, 5286.897, 5294.02, 5298.26, 5299.556, 5300.271, 
    5301.036,
  5172.854, 5187.007, 5206.907, 5220.326, 5230.471, 5238.87, 5247.091, 
    5263.788, 5278.894, 5290.09, 5299.066, 5304.24, 5308.128, 5311.642, 
    5313.863,
  5170.753, 5182.937, 5203.995, 5218.175, 5232.72, 5237.202, 5249.517, 
    5257.836, 5274.701, 5289.965, 5301.91, 5308.493, 5315.835, 5322.102, 
    5325.923,
  5172.601, 5183.566, 5203.731, 5219.771, 5232.457, 5243.738, 5247.486, 
    5262.686, 5278.038, 5289.948, 5303.888, 5313.342, 5324.413, 5332.469, 
    5337.424,
  5178.046, 5187.582, 5205.437, 5220.679, 5233.58, 5242.775, 5252.994, 
    5260.569, 5273.249, 5292.228, 5305.4, 5319.125, 5331.617, 5342.624, 
    5348.202,
  5187.005, 5195.575, 5210.832, 5223.472, 5236.031, 5247.348, 5254.516, 
    5266.46, 5279.765, 5293.312, 5308.444, 5324.034, 5338.991, 5351.27, 
    5358.839,
  5199.008, 5205.745, 5215.714, 5226.112, 5235.663, 5248.203, 5258.082, 
    5266.497, 5277.391, 5294.585, 5310.23, 5327.639, 5344.357, 5358.208, 
    5368.391,
  5208.95, 5213.72, 5220.992, 5228.733, 5236.859, 5249.751, 5260.122, 
    5271.437, 5282.702, 5295.508, 5311.163, 5330.1, 5347.673, 5363.331, 
    5375.363,
  5217.959, 5216.681, 5220.942, 5227.639, 5233.813, 5246.147, 5260.129, 
    5269.937, 5280.294, 5294.26, 5311.1, 5330.016, 5348.852, 5365.774, 
    5380.043,
  5192.384, 5205.438, 5215.158, 5224.75, 5233.345, 5240.052, 5243.388, 
    5244.624, 5242.972, 5235.956, 5226.518, 5214.022, 5199.841, 5183.782, 
    5168.864,
  5199.021, 5212.179, 5223.279, 5235.164, 5244.153, 5251.625, 5257.303, 
    5257.88, 5253.743, 5248.113, 5237.729, 5225.554, 5209.609, 5194.519, 
    5178.134,
  5205.566, 5219.032, 5231.092, 5244.436, 5254.935, 5265.354, 5269.203, 
    5272.688, 5269.524, 5261.404, 5250.039, 5237.431, 5222.654, 5206.666, 
    5190.938,
  5213.3, 5226.396, 5239.056, 5251.309, 5264.364, 5271.541, 5279.899, 
    5280.945, 5279.647, 5273.201, 5263.478, 5250.427, 5237.452, 5222.321, 
    5207.994,
  5221.381, 5233.851, 5245.186, 5257.06, 5267.042, 5277.339, 5282.323, 
    5288.116, 5290.839, 5284.379, 5276.771, 5264.917, 5254.244, 5239.292, 
    5226.601,
  5229.981, 5240.3, 5248.925, 5259.097, 5266.519, 5272.774, 5279.607, 
    5284.469, 5289.961, 5293.032, 5288.383, 5280.828, 5272.388, 5261.104, 
    5249.101,
  5236.389, 5245.388, 5251.334, 5258.739, 5264.065, 5268.586, 5270.746, 
    5278.42, 5288.415, 5296.308, 5297.727, 5296.008, 5291.599, 5284.2, 5274.32,
  5245.249, 5248.621, 5251.905, 5257.456, 5260.324, 5262.636, 5263.725, 
    5266.707, 5278.134, 5294.647, 5303.193, 5309.187, 5311.121, 5309.617, 
    5303.824,
  5252.888, 5248.955, 5250.459, 5253.612, 5257.513, 5259.897, 5259.658, 
    5262.485, 5272.241, 5290.655, 5305.022, 5318.432, 5327.104, 5331.493, 
    5330.609,
  5256.843, 5248.46, 5245.545, 5247.674, 5250.773, 5254.899, 5256.134, 
    5257.296, 5265.06, 5284.442, 5303.331, 5321.813, 5336.14, 5345.407, 
    5349.899,
  5245.714, 5251.382, 5256.781, 5257.951, 5254.151, 5244.2, 5226.433, 
    5208.703, 5190.147, 5170.822, 5155.607, 5142.221, 5131.884, 5121.303, 
    5112.952,
  5254.055, 5259.832, 5265.454, 5267.5, 5264.291, 5252.561, 5240.485, 
    5219.061, 5199.003, 5183.482, 5169.865, 5158.667, 5147.72, 5139.366, 
    5130.569,
  5261.853, 5267.823, 5272.977, 5276.75, 5272.032, 5266.896, 5247.613, 
    5234.315, 5215.811, 5198.223, 5184.817, 5175.122, 5166.261, 5157.767, 
    5149.686,
  5271.296, 5275.298, 5280.504, 5281.731, 5281.186, 5270.293, 5261.3, 
    5242.014, 5225.578, 5211.481, 5200.654, 5191.027, 5184.255, 5176.478, 
    5169.761,
  5282.146, 5283.975, 5286.732, 5287.049, 5285.61, 5278.843, 5266.948, 
    5253.226, 5243.82, 5225.342, 5216.87, 5207.673, 5203.202, 5195.937, 
    5191.14,
  5295.458, 5293.977, 5291.349, 5290.221, 5285.975, 5279.778, 5273.031, 
    5260.479, 5249.489, 5241.138, 5232.531, 5226.289, 5221.931, 5217.487, 
    5212.709,
  5307.862, 5303.92, 5296.983, 5292.693, 5286.697, 5281.212, 5274.415, 
    5268.302, 5263.282, 5255.952, 5249.601, 5246.141, 5242.819, 5240.065, 
    5235.638,
  5318.601, 5309.989, 5300.093, 5293.664, 5285.965, 5279.844, 5275.907, 
    5270.552, 5268.465, 5268.531, 5266.382, 5265.468, 5264.399, 5262.895, 
    5259.472,
  5322.581, 5311.316, 5300.638, 5292.498, 5286.596, 5280.233, 5276.083, 
    5274.514, 5276.444, 5279.735, 5281.706, 5284.617, 5286.021, 5285.755, 
    5282.938,
  5326.018, 5306.965, 5292.997, 5285.806, 5280.672, 5275.892, 5273.604, 
    5272.65, 5276.351, 5285.532, 5292.944, 5299.606, 5303.709, 5305.986, 
    5304.857,
  5286.047, 5286.089, 5279.389, 5267.708, 5254.691, 5241.557, 5228.175, 
    5218.905, 5211.26, 5202.066, 5192.552, 5182.223, 5170.966, 5156.526, 
    5141.234,
  5289.386, 5288.774, 5282.357, 5272.01, 5260.885, 5247.267, 5240.012, 
    5231.692, 5224.035, 5217.88, 5209.976, 5201.14, 5188.545, 5174.721, 
    5157.427,
  5292.017, 5291.443, 5285.95, 5278.349, 5266.672, 5259.236, 5248.211, 
    5243.581, 5239.481, 5234.688, 5227.872, 5220.077, 5208.922, 5193.379, 
    5174.53,
  5297.159, 5295.493, 5290.867, 5282.344, 5274.546, 5263.611, 5259.703, 
    5255.35, 5251.355, 5249.138, 5245.415, 5237.917, 5227.746, 5213.396, 
    5193.997,
  5305.445, 5302.949, 5298.111, 5290.668, 5282.288, 5275.327, 5268.454, 
    5264.347, 5266.351, 5262.802, 5261.165, 5254.744, 5246.928, 5231.966, 
    5214.314,
  5313.308, 5309.233, 5304.083, 5298.103, 5288.793, 5280.884, 5278.292, 
    5275.923, 5274.303, 5275.287, 5274.153, 5269.817, 5263.15, 5251.22, 
    5234.606,
  5316.578, 5309.727, 5305.792, 5303.944, 5297.745, 5290.274, 5284.526, 
    5283.837, 5284.733, 5285.509, 5285.023, 5282.914, 5277.591, 5268.526, 
    5254.337,
  5325.146, 5310.465, 5302.66, 5302.361, 5299.668, 5294.714, 5290.134, 
    5290.118, 5289.909, 5292.245, 5293.321, 5292.599, 5289.583, 5283.279, 
    5272.602,
  5345.56, 5325.15, 5308.95, 5302.488, 5302.091, 5300.154, 5293.805, 
    5294.016, 5294.909, 5296.844, 5299.027, 5299.902, 5298.848, 5295.197, 
    5287.623,
  5368.561, 5349.22, 5329.172, 5313.71, 5305.136, 5302.057, 5297.365, 
    5295.704, 5296.79, 5298.334, 5301.667, 5303.881, 5304.86, 5304.163, 
    5300.296,
  5275.86, 5275.384, 5275.735, 5279.208, 5284.864, 5290.639, 5292.921, 
    5291.918, 5286.478, 5274.062, 5255.934, 5230.146, 5200.646, 5167.651, 
    5137.034,
  5275.185, 5275.539, 5277.714, 5283.134, 5289.435, 5295.869, 5300.306, 
    5300.674, 5294.598, 5285.352, 5268.713, 5246.341, 5215.927, 5183.788, 
    5151.195,
  5275.197, 5278.432, 5282.064, 5288.543, 5294.352, 5301.81, 5305.694, 
    5306.476, 5303.426, 5294.993, 5281.369, 5261.471, 5234.688, 5201.327, 
    5167.821,
  5278.212, 5281.469, 5286.967, 5291.425, 5300.312, 5304.396, 5311.317, 
    5312.213, 5309.131, 5302.297, 5292.229, 5275.17, 5251.996, 5222.582, 
    5189.093,
  5282.329, 5287.58, 5292.696, 5297.118, 5303.139, 5310.545, 5314.079, 
    5315.154, 5314.446, 5307.554, 5300.287, 5287.195, 5269.496, 5242.292, 
    5212.761,
  5287.925, 5292.833, 5296.567, 5301.736, 5306.422, 5311.949, 5317.114, 
    5318.34, 5316.495, 5311.881, 5305.566, 5295.944, 5283.022, 5262.489, 
    5236.214,
  5291.48, 5297.318, 5300.743, 5305.014, 5308.475, 5313.753, 5316.246, 
    5318.531, 5317.502, 5314.127, 5308.642, 5302.108, 5292.584, 5277.812, 
    5256.675,
  5304.238, 5301.531, 5302.307, 5307.157, 5310.125, 5314.201, 5316.881, 
    5318.322, 5317.405, 5315.392, 5310.933, 5305.636, 5299.094, 5289.758, 
    5274.126,
  5326.863, 5320.697, 5315.542, 5313.171, 5313.803, 5315.406, 5316.562, 
    5317.676, 5316.918, 5315.642, 5312.528, 5308.328, 5302.812, 5296.289, 
    5285.798,
  5343.165, 5339.347, 5334.811, 5330.228, 5326.192, 5324.682, 5323.792, 
    5323.016, 5321.83, 5319.787, 5316.542, 5312.122, 5306.634, 5301.155, 
    5293.827,
  5251.763, 5260.902, 5269.228, 5277.066, 5288.11, 5299.447, 5308.009, 
    5312.054, 5311.063, 5302.132, 5287.738, 5266.623, 5241.256, 5209.567, 
    5177.359,
  5245.167, 5253.845, 5262.583, 5272.606, 5283.858, 5297.001, 5307.873, 
    5312.179, 5310.284, 5304.662, 5291.986, 5274.888, 5250.978, 5222.822, 
    5189.547,
  5237.389, 5246.647, 5256.537, 5269.037, 5282.602, 5297.208, 5305.062, 
    5311.613, 5309.498, 5304.488, 5294.5, 5280.439, 5260.698, 5233.213, 
    5201.235,
  5231.418, 5240.75, 5252.066, 5265.605, 5281.539, 5294.546, 5306.271, 
    5309.15, 5308.941, 5303.489, 5295.796, 5284.629, 5268.727, 5246.38, 
    5215.193,
  5227.111, 5237.185, 5249.392, 5264.746, 5280.836, 5296.641, 5303.847, 
    5308.825, 5306.753, 5301.902, 5295.577, 5286.929, 5275.517, 5255.209, 
    5229.076,
  5226.634, 5237.727, 5249.69, 5265.203, 5280.812, 5294.471, 5304.35, 
    5306.834, 5305.433, 5300.988, 5295.566, 5289.091, 5281.166, 5266.29, 
    5243.177,
  5230.159, 5241.324, 5253.09, 5267.462, 5282.26, 5294.477, 5301.26, 
    5304.509, 5302.849, 5299.071, 5295.505, 5291.7, 5285.552, 5273.674, 
    5254.646,
  5238.441, 5248.674, 5258.529, 5270.674, 5281.673, 5291.904, 5298.268, 
    5300.674, 5299.402, 5297.773, 5296, 5295.317, 5291.324, 5282.569, 5267.492,
  5249.758, 5256.78, 5264.111, 5273.378, 5282.33, 5289.633, 5293.133, 
    5294.754, 5294.988, 5296.147, 5298.121, 5299.564, 5296.59, 5288.95, 
    5276.877,
  5267.415, 5270.023, 5273.588, 5278.202, 5282.481, 5287.09, 5290.784, 
    5293.849, 5296.225, 5299.109, 5302.018, 5303.542, 5301.007, 5295.648, 
    5286.039,
  5240.426, 5254.739, 5268.713, 5281.27, 5291.639, 5297.704, 5299.336, 
    5299.871, 5295.539, 5285.706, 5273.326, 5257.298, 5235.28, 5202.33, 
    5168.703,
  5240.312, 5254.481, 5267.333, 5279.488, 5287.854, 5294.535, 5299.804, 
    5296.642, 5293.093, 5287.196, 5275.797, 5263.014, 5240.735, 5211.92, 
    5177.46,
  5237.771, 5251.519, 5264.259, 5276.653, 5286.353, 5292.788, 5292.742, 
    5299.026, 5293.899, 5287.663, 5278.953, 5268.806, 5249.321, 5221.267, 
    5189.549,
  5234.522, 5246.917, 5259.569, 5270.955, 5279.865, 5288.01, 5292.064, 
    5289.479, 5291.29, 5288.074, 5282.417, 5274.755, 5259.305, 5236.167, 
    5207.143,
  5229.445, 5241.11, 5252.788, 5265.016, 5273.91, 5281.082, 5286.609, 
    5291.935, 5291.174, 5287.456, 5285.181, 5280.534, 5268.969, 5248.25, 
    5224.75,
  5223.088, 5234.341, 5244.505, 5255.168, 5264.914, 5273.135, 5280.833, 
    5284.704, 5287.8, 5287.855, 5286.32, 5285.467, 5277.979, 5262.88, 5242.982,
  5215.365, 5226.282, 5236.184, 5246.496, 5256.751, 5267.151, 5274.681, 
    5282.98, 5286.344, 5285.33, 5285.919, 5288.358, 5284.211, 5272.805, 
    5257.274,
  5208.197, 5218.368, 5227.299, 5237.239, 5246.843, 5258.285, 5268.209, 
    5275.191, 5280.447, 5282.688, 5283.761, 5288.683, 5288.849, 5282.636, 
    5270.78,
  5203.366, 5212.855, 5221.81, 5231.834, 5242.805, 5253.646, 5263.269, 
    5271.636, 5275.877, 5276.535, 5278.865, 5286.035, 5289.636, 5286.758, 
    5279.196,
  5203.491, 5211.044, 5218.999, 5228.037, 5238.06, 5248.763, 5258.043, 
    5264.233, 5268.178, 5270.687, 5274.191, 5282.211, 5287.81, 5288.456, 
    5284.163,
  5249.843, 5262.465, 5273.87, 5280.917, 5286.406, 5287.833, 5285.498, 
    5281.08, 5274.612, 5265.375, 5254.438, 5240.072, 5223.165, 5203.435, 
    5182.851,
  5257.386, 5268.612, 5278.341, 5284.423, 5288.618, 5290.567, 5291.464, 
    5285.134, 5278.958, 5273.957, 5265.377, 5254.501, 5238.778, 5223.438, 
    5203.328,
  5261.681, 5271.672, 5280.183, 5286.549, 5290.86, 5293.722, 5292.104, 
    5292.554, 5286.956, 5280.917, 5273.979, 5265.333, 5253.327, 5238.332, 
    5220.104,
  5265.013, 5272.916, 5280.274, 5285.881, 5289.485, 5293.253, 5293.625, 
    5289.188, 5284.924, 5285.052, 5280.288, 5273.648, 5264.075, 5252.712, 
    5236.466,
  5266.04, 5272.431, 5277.875, 5283.208, 5288.002, 5290.345, 5291.59, 
    5292.044, 5291.055, 5284.935, 5284.34, 5278.725, 5272.265, 5261.616, 
    5249.028,
  5265.087, 5269.762, 5273.923, 5277.268, 5281.295, 5284.855, 5286.717, 
    5285.57, 5284.653, 5283.909, 5284.239, 5282.19, 5277.583, 5270.851, 
    5260.545,
  5260.104, 5263.78, 5266.766, 5269.806, 5273.014, 5276.939, 5279.845, 
    5282.21, 5282.279, 5281.468, 5280.666, 5281.438, 5279.41, 5275.035, 
    5267.687,
  5251.095, 5254.042, 5256.635, 5259.331, 5261.796, 5265.104, 5269.352, 
    5271.485, 5273.175, 5275.083, 5275.451, 5277.851, 5279.462, 5278.201, 
    5274.269,
  5237.33, 5240.332, 5243.367, 5246.604, 5249.706, 5253.264, 5256.766, 
    5261.171, 5264.501, 5266.571, 5267.986, 5270.778, 5274.527, 5276.711, 
    5275.671,
  5223.299, 5225.555, 5228.62, 5231.765, 5234.328, 5237.743, 5241.48, 
    5245.518, 5250.028, 5255.177, 5258.867, 5261.993, 5267.755, 5273.376, 
    5275.691,
  5230.404, 5243.575, 5255.063, 5262.056, 5266.922, 5267.575, 5264.476, 
    5260.01, 5252.032, 5238.927, 5223.808, 5203.75, 5178.957, 5144.257, 
    5105.12,
  5243.954, 5255.89, 5265.736, 5271.428, 5274.795, 5273.187, 5271.795, 
    5263.397, 5253.788, 5243.789, 5228.844, 5211.086, 5186.249, 5156.041, 
    5117.616,
  5254.946, 5266.055, 5273.957, 5279.56, 5280.323, 5281.69, 5274.765, 
    5271.599, 5261.528, 5249.104, 5234.337, 5218.042, 5195.751, 5167.114, 
    5131.293,
  5264.501, 5272.295, 5278.662, 5282.755, 5284.705, 5282.484, 5279.51, 
    5270.829, 5260.393, 5251.915, 5239.11, 5224.241, 5205.673, 5181.847, 
    5149.819,
  5269.225, 5276.06, 5281.249, 5285.154, 5286.554, 5285.393, 5279.236, 
    5273.664, 5266.013, 5253.385, 5243.172, 5229.994, 5215.249, 5194.334, 
    5168.819,
  5272.328, 5277.868, 5281.47, 5284.384, 5283.585, 5281.51, 5276.477, 
    5268.299, 5259.315, 5252.089, 5243.99, 5234.518, 5223.216, 5209.158, 
    5189.492,
  5271.87, 5276.634, 5279.029, 5280.222, 5278.688, 5274.725, 5268.555, 
    5262.886, 5256.095, 5249.037, 5242.571, 5236.311, 5228.175, 5219.346, 
    5206.267,
  5270.124, 5272.065, 5272.264, 5271.16, 5267.238, 5262.519, 5256.353, 
    5249.937, 5243.675, 5239.693, 5236.817, 5234.186, 5230.928, 5226.879, 
    5220.396,
  5262.498, 5262.459, 5260.834, 5257.464, 5252.567, 5246.77, 5239.814, 
    5234.562, 5230.734, 5228.041, 5227.717, 5228.291, 5228.413, 5228.586, 
    5227.87,
  5250.296, 5246.404, 5241.75, 5237.071, 5230.811, 5225.419, 5220.595, 
    5216.823, 5214.113, 5213.78, 5214.985, 5218.611, 5222.401, 5226.681, 
    5231.1,
  5222.274, 5234.953, 5245.081, 5250.515, 5252.183, 5247.919, 5237.128, 
    5223.309, 5204.506, 5180.521, 5156.657, 5131.463, 5110.468, 5093.508, 
    5081.869,
  5235.162, 5246.94, 5256.185, 5260.949, 5261.344, 5255.113, 5246.755, 
    5228.175, 5208.709, 5190.274, 5169.125, 5147.171, 5126.549, 5112.619, 
    5102.437,
  5245.717, 5257.933, 5265.455, 5270.227, 5267.675, 5265.193, 5250.652, 
    5240.905, 5221.751, 5200.412, 5181.572, 5162.358, 5144.318, 5131.272, 
    5122.172,
  5255.834, 5266.132, 5272.458, 5275.31, 5274.72, 5266.23, 5258.266, 5238.84, 
    5221.31, 5206.992, 5192.018, 5176.338, 5161.025, 5149.257, 5142.932,
  5263.529, 5271.776, 5276.902, 5278.54, 5276.057, 5270.814, 5257.029, 
    5247.026, 5230.775, 5210.683, 5200.105, 5187.93, 5176.647, 5166.194, 
    5161.545,
  5268.829, 5275.124, 5277.886, 5278.572, 5274.548, 5267.062, 5256.038, 
    5238.822, 5222.29, 5211.791, 5204.07, 5197.014, 5188.88, 5181.646, 
    5178.469,
  5270.641, 5275.639, 5276.544, 5275.045, 5269.839, 5261.163, 5248.534, 
    5236.328, 5222.651, 5209.274, 5204.781, 5202.668, 5198.036, 5193.662, 
    5191.778,
  5269.952, 5272.006, 5270.795, 5267.774, 5260.67, 5251.322, 5238.916, 
    5224.552, 5210.896, 5203.725, 5202.7, 5204.753, 5204.977, 5203.439, 
    5204.232,
  5264.199, 5265.038, 5262.499, 5257.749, 5250.084, 5240.093, 5228.963, 
    5218.546, 5208.621, 5201.071, 5199.656, 5203.994, 5208.402, 5210.1, 
    5212.85,
  5255.861, 5254.3, 5250.144, 5245.59, 5238.142, 5230.783, 5222.93, 5213.558, 
    5204.57, 5199.004, 5197.291, 5202.19, 5208.414, 5213.464, 5218.468,
  5277.063, 5281.623, 5281.402, 5273.778, 5261.999, 5245.187, 5224.044, 
    5206.8, 5191.819, 5178.229, 5167.671, 5157.44, 5145.125, 5129.858, 
    5110.511,
  5283.711, 5288.588, 5287.582, 5281.045, 5269.045, 5249.729, 5235.595, 
    5211.227, 5193.445, 5183.919, 5174.413, 5165.69, 5154.127, 5140.584, 
    5122.132,
  5287.635, 5293.384, 5291.784, 5287.407, 5273.435, 5262.165, 5235.423, 
    5224.444, 5202.303, 5188.406, 5179.872, 5172.238, 5162.742, 5149.415, 
    5131.572,
  5290.22, 5295.183, 5294.816, 5289.693, 5279.297, 5260.547, 5247.322, 
    5222.165, 5204.003, 5190.932, 5183.684, 5176.924, 5169.633, 5159.382, 
    5143.321,
  5289.838, 5294.816, 5295.489, 5290.607, 5281.036, 5266.566, 5246.492, 
    5231.908, 5212.235, 5193.41, 5187.139, 5180.228, 5175.864, 5166.357, 
    5154.135,
  5287.228, 5292.712, 5293.447, 5289.764, 5279.272, 5265.126, 5249.59, 
    5230.333, 5211.146, 5197.455, 5189.414, 5182.762, 5180.04, 5174.433, 
    5165.018,
  5282.541, 5288.575, 5290.087, 5285.757, 5276.98, 5263.5, 5248.732, 5235.03, 
    5218.262, 5201.374, 5191.637, 5185.256, 5182.015, 5179.761, 5173.471,
  5277.21, 5282.81, 5284.044, 5279.927, 5270.523, 5258.872, 5247.412, 
    5233.127, 5217.542, 5203.209, 5193.06, 5186.591, 5183.612, 5183.452, 
    5181.321,
  5270.13, 5275.657, 5276.276, 5271.519, 5264.11, 5254.306, 5244.609, 
    5233.516, 5219.706, 5203.979, 5192.104, 5186.55, 5183.397, 5183.71, 
    5185.259,
  5263.209, 5266.496, 5265.813, 5261.985, 5254.349, 5247.114, 5238.283, 
    5225.708, 5212.393, 5200.115, 5189.35, 5184.226, 5182.164, 5182.617, 
    5186.999,
  5297.39, 5299.072, 5298.632, 5292.287, 5283.429, 5269.472, 5251.694, 
    5233.711, 5211.77, 5183.736, 5160.298, 5135.355, 5109.747, 5078.981, 
    5044.902,
  5292.872, 5295.721, 5295.68, 5291.195, 5283.158, 5267.958, 5256.326, 
    5230.514, 5208.009, 5186.792, 5162.396, 5136.788, 5109.464, 5080.505, 
    5044.776,
  5286.226, 5290.632, 5291.215, 5289.374, 5280.313, 5272.289, 5250.681, 
    5241.168, 5216.673, 5190.192, 5163.976, 5139.023, 5109.967, 5080.557, 
    5045.886,
  5279, 5283.245, 5284.94, 5283.233, 5277.321, 5264.646, 5254.709, 5230.601, 
    5211.128, 5193.036, 5165.814, 5140.262, 5112.07, 5084.418, 5051.19,
  5269.542, 5274.105, 5277.063, 5275.768, 5271.462, 5262.255, 5246.728, 
    5236.124, 5217.154, 5190.188, 5168.38, 5140.831, 5114.774, 5086.499, 
    5058.025,
  5259.606, 5263.637, 5265.977, 5265.659, 5260.8, 5252.811, 5241.84, 
    5223.377, 5206.114, 5189.341, 5167.309, 5142.13, 5117.213, 5092.311, 
    5066.38,
  5248.89, 5252.48, 5254.4, 5253.74, 5250.252, 5242.373, 5231.247, 5220.579, 
    5205.156, 5185.086, 5164.707, 5142.494, 5118.422, 5096.526, 5074.36,
  5239.938, 5241.177, 5241.049, 5240.421, 5235.396, 5228.815, 5219.092, 
    5205.978, 5191.792, 5177.982, 5160.158, 5140.05, 5119.759, 5101.509, 
    5084.487,
  5233.479, 5233.583, 5232.134, 5228.731, 5223.66, 5216.211, 5206.226, 
    5197.088, 5185.127, 5169.857, 5153.391, 5135.851, 5118.723, 5104.191, 
    5092.696,
  5232.644, 5228.138, 5223.251, 5218.662, 5210.997, 5201.925, 5192.3, 
    5180.915, 5169.313, 5158.424, 5144.38, 5128.977, 5115.912, 5106.584, 
    5101.105,
  5281.218, 5276.957, 5274.274, 5270.771, 5266.627, 5259.299, 5248.202, 
    5238.133, 5223.783, 5202.497, 5181.308, 5158.146, 5131.968, 5102.703, 
    5069.742,
  5272.461, 5268.619, 5265.436, 5260.644, 5254.925, 5245.54, 5239.006, 
    5220.961, 5206.686, 5193.804, 5172.432, 5150.396, 5124.207, 5099.736, 
    5063.798,
  5267.511, 5262.524, 5257.912, 5253.106, 5243.796, 5239.299, 5222.366, 
    5220.728, 5200.69, 5181.929, 5161.979, 5143.215, 5117.719, 5092.61, 
    5058.345,
  5263.383, 5256.81, 5250.697, 5243.867, 5236.521, 5224.765, 5219.056, 
    5197.066, 5186.51, 5173.692, 5152.502, 5134.622, 5112.194, 5088.606, 
    5055.298,
  5262.564, 5255.016, 5246.985, 5238.883, 5229.905, 5220.016, 5204.919, 
    5197.09, 5179.415, 5159.204, 5144.983, 5125.576, 5106.584, 5081.614, 
    5052.418,
  5264.369, 5254.986, 5244.132, 5234.44, 5221.906, 5210.218, 5196.701, 
    5177.756, 5162.499, 5149.641, 5132.457, 5116.648, 5098.705, 5077.008, 
    5049.225,
  5268.796, 5257.954, 5244.544, 5231.674, 5217.217, 5202.194, 5185.033, 
    5170.617, 5152.3, 5133.606, 5119.204, 5105.373, 5088.984, 5069.81, 5044.12,
  5272.726, 5258.862, 5242.577, 5227.142, 5208.681, 5191.682, 5171.856, 
    5151.656, 5132.134, 5117.073, 5102.187, 5090.486, 5077.882, 5062.541, 
    5040.222,
  5274.462, 5259.167, 5241.364, 5222.172, 5202.023, 5180.682, 5157.664, 
    5137.049, 5116.004, 5096.752, 5083.736, 5075.108, 5065.598, 5053.549, 
    5035.061,
  5272.007, 5252.312, 5232.415, 5211.758, 5187.965, 5164.478, 5139.969, 
    5114.888, 5093.181, 5077.172, 5066.243, 5059.666, 5053.277, 5044.931, 
    5030.801,
  5247.519, 5243.82, 5241.659, 5239.821, 5239.079, 5237.379, 5234.385, 
    5231.862, 5225.039, 5212.034, 5198.766, 5183.333, 5166.209, 5144.132, 
    5123.599,
  5251.107, 5246.157, 5243.507, 5240.976, 5239.461, 5235.875, 5234.764, 
    5224.654, 5216.943, 5209.376, 5193.226, 5175.771, 5154.658, 5134.603, 
    5110.349,
  5259.21, 5252.996, 5248.687, 5245.955, 5240.372, 5239.743, 5230.691, 
    5230.104, 5216.322, 5199.78, 5182.489, 5163.92, 5139.253, 5117.428, 
    5096.805,
  5266.31, 5259.05, 5253.973, 5248.732, 5245.336, 5236.464, 5233.163, 
    5216.752, 5206.383, 5195.471, 5170.09, 5146.867, 5121.932, 5099.578, 
    5083.744,
  5269.522, 5262.181, 5256.215, 5250.339, 5243.911, 5237.795, 5226.575, 
    5218.441, 5201.068, 5176.838, 5156.534, 5127.25, 5101.733, 5080.917, 
    5072.199,
  5265.218, 5258.143, 5252.126, 5246.533, 5239.203, 5230.821, 5219.742, 
    5204.613, 5186.06, 5165.899, 5137.382, 5108.891, 5081.611, 5067.738, 
    5063.258,
  5252.57, 5246.414, 5240.538, 5236.088, 5229.361, 5221.482, 5209.789, 
    5196.205, 5174.534, 5148.68, 5120.003, 5091.396, 5064.733, 5057.265, 
    5056.452,
  5234.598, 5228.083, 5222.224, 5219.892, 5213.878, 5207.544, 5194.776, 
    5179.185, 5158.178, 5136.101, 5105.225, 5076.898, 5054.043, 5051.324, 
    5053.683,
  5212.994, 5206.74, 5202.032, 5199.809, 5195.553, 5190.158, 5179.574, 
    5166.917, 5145.985, 5121.709, 5092.551, 5067.386, 5048.121, 5048.847, 
    5052.994,
  5191.191, 5183.183, 5178.706, 5177.079, 5174.043, 5169.965, 5161.11, 
    5148.43, 5130.38, 5109.844, 5083.407, 5061.424, 5047.13, 5049.788, 
    5053.629,
  5228.762, 5219.91, 5213.69, 5211.3, 5213.462, 5218.079, 5224.466, 5231.421, 
    5235.199, 5235.623, 5232.128, 5223.748, 5206.036, 5181.104, 5152.628,
  5229.608, 5221.052, 5215.69, 5212.356, 5211.71, 5215.639, 5221.391, 
    5225.83, 5229.629, 5232.643, 5226.058, 5217.139, 5196.6, 5172.952, 
    5137.749,
  5227.065, 5218.874, 5214.09, 5212.243, 5211.686, 5214.812, 5217.337, 
    5225.177, 5226.033, 5226.406, 5220.982, 5210.574, 5189.185, 5162.202, 
    5127.738,
  5216.752, 5208.862, 5204.678, 5203.743, 5205.179, 5206.741, 5212.173, 
    5211.077, 5218.542, 5218.343, 5213.337, 5202.43, 5182.8, 5156.345, 
    5123.846,
  5203.173, 5194.98, 5190.111, 5189.403, 5190.688, 5195.117, 5197.625, 
    5208.263, 5206.115, 5209.026, 5205.805, 5195.01, 5176.832, 5151.26, 
    5124.383,
  5188.243, 5177.935, 5170.313, 5168.432, 5168.362, 5172.822, 5179.837, 
    5183.616, 5192.658, 5196.154, 5193.617, 5186.845, 5171.25, 5149.233, 
    5126.139,
  5171.63, 5159.516, 5149.083, 5143.214, 5141.838, 5145.695, 5153.285, 
    5166.147, 5173.439, 5178.054, 5182.85, 5177.446, 5164.878, 5145.789, 
    5127.722,
  5153.96, 5137.848, 5122.715, 5114.1, 5109.513, 5113.082, 5121.546, 
    5132.843, 5147.247, 5160.629, 5166.372, 5165.381, 5158.175, 5142.865, 
    5128.719,
  5135.67, 5116.436, 5097.573, 5083.996, 5078.051, 5080.161, 5089.489, 
    5105.419, 5122.504, 5136.574, 5148.712, 5152.862, 5149.349, 5138.014, 
    5128.041,
  5121.864, 5096.868, 5073.785, 5060.333, 5054.359, 5055.15, 5063.233, 
    5076.412, 5096.176, 5116.088, 5131.388, 5138.76, 5140.424, 5132.794, 
    5126.378,
  5180.27, 5180.952, 5177.129, 5172.559, 5172.58, 5183.149, 5197.637, 
    5215.868, 5234.411, 5249.079, 5256.522, 5258.363, 5248.831, 5232.56, 
    5209.271,
  5172.116, 5177.03, 5176.242, 5174.681, 5172.105, 5181.821, 5195.746, 
    5213.041, 5229.958, 5247.419, 5254.252, 5257.508, 5247.605, 5236.352, 
    5212.226,
  5163.067, 5170.188, 5174.845, 5175.475, 5176.394, 5183.038, 5194.028, 
    5212.845, 5228.185, 5242.538, 5250.741, 5254.949, 5247.507, 5237.188, 
    5215.702,
  5151.46, 5158.931, 5166.773, 5171.909, 5177.58, 5180.779, 5192.875, 
    5200.865, 5219.801, 5234.077, 5244.963, 5249.585, 5246.373, 5238.924, 
    5220.384,
  5141.406, 5148.624, 5157.063, 5166.109, 5172.664, 5182.106, 5185.215, 
    5201.23, 5211.072, 5224.196, 5235.685, 5242.732, 5243.077, 5238.763, 
    5223.982,
  5130.844, 5137.687, 5145.703, 5155.798, 5164.518, 5172.625, 5182.724, 
    5189.285, 5200.297, 5214.075, 5222.927, 5233.956, 5237.591, 5238.259, 
    5227.188,
  5122.014, 5125.957, 5134.124, 5143.4, 5152.982, 5163.23, 5171.183, 
    5183.637, 5193.224, 5201.085, 5213.605, 5223.829, 5231.504, 5235.808, 
    5228.955,
  5117.701, 5115.094, 5119.305, 5129.424, 5136.968, 5146.696, 5155.675, 
    5164.331, 5175.485, 5189.914, 5201.139, 5212.643, 5224.438, 5232.405, 
    5230.726,
  5123.647, 5114.233, 5110.288, 5113.506, 5119.581, 5126.924, 5135.297, 
    5147.269, 5159.206, 5171.83, 5186.891, 5202.541, 5216.249, 5227.68, 
    5230.945,
  5136.955, 5121.29, 5111.661, 5107.243, 5105.218, 5107.121, 5111.968, 
    5118.871, 5131.402, 5150.116, 5170.308, 5189.357, 5207.038, 5222.521, 
    5230.135,
  5166.443, 5176.715, 5178.353, 5176.41, 5182.771, 5194.721, 5212.447, 
    5231.94, 5248.074, 5257.18, 5259.762, 5260.392, 5259.748, 5260.354, 
    5263.69,
  5163.791, 5175.647, 5177.819, 5176.208, 5179.634, 5194.903, 5214.743, 
    5233.191, 5249.041, 5262.979, 5267.715, 5269.73, 5269.513, 5271.801, 
    5275.119,
  5161.693, 5174.913, 5179.393, 5177.432, 5181.781, 5198.221, 5216.36, 5240, 
    5258.969, 5269.481, 5275.254, 5278.048, 5279.882, 5281.311, 5284.94,
  5159.071, 5172.783, 5180.298, 5179.492, 5187.15, 5196.544, 5224.451, 
    5237.845, 5258.786, 5271.999, 5281.903, 5284.327, 5287.055, 5289.771, 
    5293.886,
  5156.231, 5171.868, 5180.165, 5185.262, 5188.144, 5209.114, 5220.508, 
    5249.346, 5264.931, 5276.845, 5284.965, 5289.966, 5292.989, 5295.799, 
    5299.789,
  5154.062, 5170.16, 5179.967, 5187.712, 5193.326, 5205.876, 5229.537, 
    5243.235, 5259.282, 5278.263, 5285.14, 5292.569, 5294.583, 5300.783, 
    5303.697,
  5152.873, 5168.857, 5180.624, 5189.705, 5197.927, 5211.417, 5225.943, 
    5248.038, 5265, 5275.157, 5285.994, 5292.283, 5296.893, 5303.112, 5306.25,
  5152.22, 5166.289, 5177.784, 5189.44, 5197.204, 5210.453, 5225.708, 
    5238.613, 5252.886, 5270.271, 5281.322, 5289.789, 5296.69, 5304.356, 
    5308.57,
  5153.568, 5164.005, 5174.582, 5186.144, 5196.617, 5207.729, 5220.825, 
    5237.843, 5251.744, 5263.511, 5274.599, 5287.031, 5295.427, 5305.14, 
    5310.016,
  5158.061, 5160.572, 5166.67, 5176.67, 5187.219, 5199.875, 5212.606, 
    5225.595, 5238.556, 5255.227, 5269.112, 5282.754, 5293.333, 5305.479, 
    5311.778,
  5179.295, 5188.037, 5196.963, 5208.076, 5218.706, 5228.229, 5237.067, 
    5247.824, 5260.752, 5272.379, 5284.86, 5297.944, 5307.689, 5316.051, 
    5320.374,
  5185.59, 5194.024, 5203.247, 5214.847, 5224.227, 5234.959, 5246.198, 
    5256.984, 5268.495, 5284.483, 5298.092, 5311.296, 5320.621, 5328.816, 
    5333.195,
  5193.289, 5202.824, 5213.074, 5224.759, 5233.691, 5247.035, 5254.564, 
    5269.806, 5284.804, 5296.701, 5310.554, 5322.482, 5332.851, 5339.699, 
    5344.627,
  5203.27, 5212.369, 5222.948, 5231.547, 5246.359, 5250.931, 5269.289, 
    5276.313, 5291.164, 5306.269, 5320.969, 5331.632, 5342.029, 5348.989, 
    5354.71,
  5212.955, 5222.152, 5230.84, 5241.187, 5250.793, 5269.097, 5276.354, 
    5293.407, 5308.586, 5316.949, 5330.298, 5339.981, 5350.303, 5356.374, 
    5362.861,
  5222.059, 5230.933, 5236.054, 5246.409, 5259.292, 5274.052, 5293.525, 
    5302.729, 5312.585, 5327.398, 5337.792, 5347.687, 5356.513, 5363.904, 
    5370.292,
  5229.751, 5238.742, 5244.224, 5252.589, 5268.949, 5288.342, 5300.837, 
    5317.776, 5330.879, 5338.196, 5346.577, 5354.77, 5363.08, 5370.14, 
    5376.742,
  5237.109, 5245.096, 5250.399, 5259.516, 5275.738, 5296.598, 5313.774, 
    5325.61, 5334.976, 5345.603, 5353.358, 5360.771, 5368.437, 5375.666, 
    5382.921,
  5241.519, 5251.522, 5260.001, 5270.45, 5287.793, 5306.995, 5323.088, 
    5338.366, 5348.753, 5354.489, 5360.06, 5366.498, 5372.841, 5380.207, 
    5387.645,
  5245.331, 5256.347, 5265.812, 5278.788, 5296.194, 5316.149, 5332.591, 
    5343.944, 5351.257, 5358.526, 5364.104, 5370.071, 5376.392, 5384.041, 
    5392.186,
  5240.112, 5251.866, 5264.082, 5275.493, 5283.355, 5290.862, 5301.363, 
    5313.294, 5322.33, 5326.989, 5330.083, 5333.201, 5335, 5336.209, 5336.493,
  5236.513, 5250.23, 5264.1, 5277.718, 5284.743, 5296.09, 5311.351, 5324.758, 
    5333.318, 5343.018, 5348.009, 5352.631, 5354.023, 5356.1, 5356.787,
  5234.443, 5250.496, 5266.021, 5280.355, 5288.604, 5305.362, 5319.176, 
    5337.038, 5350.112, 5357.908, 5364.211, 5368.78, 5372.472, 5374.412, 
    5375.841,
  5235.08, 5251.203, 5269.1, 5280.727, 5297.417, 5307.25, 5332.784, 5343.915, 
    5359.016, 5369.288, 5378.347, 5382.692, 5387.702, 5390.472, 5394.226,
  5237.257, 5254.351, 5272.229, 5286.388, 5300.442, 5324.022, 5338.823, 
    5358.505, 5374.094, 5380.539, 5389.783, 5394.105, 5400.648, 5403.901, 
    5409.159,
  5242.277, 5259.454, 5274.413, 5290.629, 5307.614, 5327.57, 5353.244, 
    5365.849, 5378.468, 5390.997, 5397.628, 5403.643, 5409.771, 5415.724, 
    5422.324,
  5249.745, 5266.83, 5281.612, 5296.715, 5316.872, 5340.938, 5358.766, 
    5378.417, 5392.387, 5398.752, 5404.36, 5410.429, 5417.031, 5424.607, 
    5432.078,
  5258.803, 5274.22, 5288.839, 5306.271, 5325.439, 5348.852, 5369.22, 
    5383.07, 5393.34, 5402.842, 5409.252, 5415.251, 5422.207, 5430.904, 
    5440.074,
  5268.702, 5284.815, 5301.382, 5319.617, 5340.57, 5360.002, 5376.014, 
    5391.396, 5401.668, 5407.854, 5413.308, 5419.499, 5426.138, 5434.861, 
    5444.638,
  5280.459, 5296.537, 5314.03, 5333.296, 5352.585, 5370.551, 5384.717, 
    5394.314, 5401.911, 5409.703, 5416.377, 5422.738, 5429.174, 5437.596, 
    5447.791,
  5330.029, 5328.655, 5329.221, 5330.101, 5331.757, 5333.585, 5333.157, 
    5333.634, 5335.52, 5335.011, 5334.288, 5334.414, 5335.211, 5336.735, 
    5340.983,
  5336.923, 5337.289, 5339.112, 5342.858, 5346.072, 5347.898, 5351.479, 
    5353.715, 5352.224, 5353.489, 5351.961, 5351.56, 5349.957, 5351.81, 
    5356.164,
  5342.023, 5344.667, 5348.456, 5354.995, 5357.811, 5365.524, 5365.351, 
    5369.693, 5371.817, 5372.119, 5369.882, 5368, 5366.219, 5366.896, 5371.729,
  5345.73, 5348.854, 5356.612, 5362.163, 5372.425, 5374.582, 5382.62, 
    5385.477, 5387.398, 5388.186, 5388.392, 5384.527, 5383.495, 5384.616, 
    5392.208,
  5347.36, 5352.423, 5362.476, 5370.391, 5380.179, 5389.116, 5395.848, 
    5397.672, 5406.145, 5404.476, 5406.557, 5402.805, 5403.725, 5403.664, 
    5413.415,
  5346.623, 5354.695, 5364.813, 5375.607, 5387.092, 5396.442, 5406.806, 
    5413.74, 5416.429, 5420.37, 5422.393, 5422.06, 5422.988, 5425.92, 5434.16,
  5345.283, 5357.011, 5368.963, 5379.761, 5391.521, 5405.554, 5414.025, 
    5422.73, 5429.842, 5433.597, 5436.202, 5439.635, 5441.58, 5445.903, 
    5452.587,
  5343.806, 5357.442, 5370.459, 5382.831, 5394.913, 5408.944, 5421.311, 
    5431.363, 5436.557, 5442.243, 5447.418, 5452.591, 5457.292, 5462.771, 
    5469.189,
  5342.451, 5358.555, 5374.188, 5385.908, 5399.655, 5414.915, 5426.225, 
    5436.55, 5443.604, 5448.923, 5454.276, 5461.466, 5468.219, 5474.778, 
    5480.816,
  5340.567, 5357.616, 5373.945, 5387.463, 5402.642, 5418.813, 5432.26, 
    5441.774, 5446.193, 5451.213, 5457.654, 5465.47, 5473.582, 5482.157, 
    5489.213,
  5308.567, 5307.993, 5307.438, 5307.585, 5309.482, 5313.463, 5317.985, 
    5327.013, 5338.665, 5351.071, 5365.227, 5381.955, 5399.473, 5417.17, 
    5435.825,
  5321.622, 5322.442, 5322.452, 5323.44, 5324.514, 5326.498, 5332.784, 
    5339.43, 5348.021, 5362.765, 5377.605, 5396.707, 5414.904, 5436.91, 
    5455.023,
  5334.289, 5336.895, 5338.073, 5340.308, 5339.268, 5344.305, 5343.555, 
    5352.897, 5362.213, 5373.564, 5388.402, 5407.927, 5429.651, 5450.845, 
    5471.807,
  5346.87, 5350.065, 5353.643, 5353.938, 5357.297, 5353.641, 5359.184, 
    5359.632, 5366.71, 5379.569, 5396.732, 5416.889, 5441.496, 5465.637, 
    5487.698,
  5357.767, 5362.441, 5366.782, 5368.811, 5369.064, 5369.877, 5367.244, 
    5369.167, 5379.556, 5386.07, 5404.372, 5425.492, 5451.871, 5475.622, 
    5499.106,
  5367.805, 5374.092, 5378.4, 5381.888, 5381.823, 5379.473, 5379.174, 
    5378.653, 5380.857, 5395.732, 5412.343, 5435.769, 5461.423, 5487.547, 
    5509.473,
  5377.488, 5384.912, 5390.311, 5394.323, 5394.386, 5393.051, 5388.564, 
    5390.494, 5397.036, 5407.072, 5424.179, 5447.502, 5472.343, 5496.925, 
    5517.183,
  5386.709, 5394.104, 5400.108, 5405.257, 5406.381, 5405.174, 5403.431, 
    5403.086, 5406.742, 5419.931, 5438.236, 5460.414, 5484.071, 5506.762, 
    5524.926,
  5395.051, 5402.467, 5409.819, 5414.958, 5418.354, 5418.758, 5417.303, 
    5419.547, 5426.205, 5437.423, 5453.627, 5474.75, 5495.691, 5514.86, 
    5530.265,
  5401.742, 5408.901, 5416.579, 5422.427, 5427.395, 5430.342, 5432.068, 
    5434.104, 5439.867, 5452.176, 5468.638, 5487.137, 5505.513, 5522.314, 
    5534.759,
  5279.298, 5286.591, 5295.213, 5304.855, 5315.617, 5326.273, 5337.517, 
    5352.788, 5369.523, 5386.384, 5406.951, 5429.469, 5450.629, 5468.962, 
    5483.907,
  5290.241, 5297.826, 5306.131, 5316.768, 5326.522, 5337.798, 5353.895, 
    5368.445, 5385.037, 5409.106, 5431.485, 5455.73, 5474.913, 5492.955, 
    5505.776,
  5300.778, 5308.389, 5316.995, 5327.911, 5338.501, 5354.867, 5366.698, 
    5389.9, 5411.064, 5431.578, 5454.819, 5476.716, 5497.129, 5513.335, 
    5526.355,
  5311.77, 5318.31, 5328.252, 5336.947, 5352.915, 5361.221, 5386.413, 
    5398.915, 5422.468, 5448.724, 5473.572, 5495.023, 5515.861, 5531.625, 
    5542.831,
  5321.357, 5328.214, 5336.522, 5347.285, 5359.413, 5379.025, 5392.147, 
    5419.135, 5446.651, 5463.857, 5490.148, 5510.621, 5531.746, 5544.808, 
    5554.775,
  5330.958, 5337.195, 5343.128, 5353.465, 5365.763, 5381.445, 5405.524, 
    5424.273, 5447.057, 5478.646, 5501.419, 5524.323, 5543.007, 5556.592, 
    5563.439,
  5339.724, 5345.233, 5349.833, 5357.494, 5369.478, 5387.817, 5407.645, 
    5437.146, 5465.805, 5488.639, 5512.11, 5535.009, 5552.277, 5563.932, 
    5568.299,
  5349.897, 5353.183, 5355.746, 5361.493, 5369.593, 5386.55, 5411.099, 
    5435.627, 5462.479, 5493.392, 5519.265, 5541.524, 5558.438, 5568.862, 
    5571.742,
  5358.354, 5360.707, 5362.258, 5364.297, 5371.978, 5386.664, 5409.852, 
    5441.017, 5472.232, 5499.225, 5523.901, 5546.3, 5562.116, 5571.437, 
    5572.851,
  5365.575, 5366.852, 5367.214, 5367.032, 5371.168, 5385.274, 5409.361, 
    5437.675, 5468.193, 5499.396, 5526.64, 5548.671, 5564.164, 5572.535, 
    5573.733,
  5267.594, 5276.451, 5291.233, 5307.388, 5324.418, 5340.968, 5359.341, 
    5381.324, 5401.738, 5416.643, 5428.011, 5434.999, 5438.333, 5437.896, 
    5435.721,
  5275.511, 5283.5, 5296.978, 5313.73, 5328.585, 5346.414, 5369.282, 5390.49, 
    5411.058, 5432.181, 5443.959, 5452.105, 5453.753, 5453.732, 5450.938,
  5283.536, 5290.836, 5304.417, 5319.723, 5335.135, 5357.65, 5376.131, 
    5406.996, 5431.454, 5447.36, 5460.412, 5467.635, 5471.774, 5472.293, 
    5469.496,
  5291.305, 5298.598, 5311.652, 5324.512, 5344.465, 5357.863, 5392.897, 
    5411.026, 5438.492, 5460.639, 5475.711, 5483.43, 5488.941, 5489.429, 
    5490.085,
  5297.763, 5306.581, 5318.375, 5333.336, 5350.507, 5375.771, 5395.269, 
    5432.418, 5459.878, 5473.514, 5490.138, 5498.337, 5506.028, 5506.096, 
    5507.668,
  5303.944, 5313.674, 5324.489, 5339.671, 5357.611, 5378.525, 5411.629, 
    5434.645, 5460.386, 5487.373, 5501.825, 5513.129, 5519.083, 5522.421, 
    5523.543,
  5309.023, 5319.813, 5331.614, 5346.353, 5365.771, 5389.62, 5415.309, 
    5450.115, 5478.714, 5497.099, 5513.14, 5525.206, 5531.614, 5535.015, 
    5536.508,
  5313.595, 5324.687, 5336.052, 5351.188, 5368.278, 5392.532, 5422.557, 
    5449.264, 5475.316, 5502.05, 5520.532, 5533.356, 5541.278, 5545.411, 
    5547.707,
  5316.633, 5328.192, 5341.01, 5356.257, 5374.795, 5396.298, 5423.092, 
    5455.85, 5484.15, 5506.315, 5524.985, 5539.633, 5548.052, 5552.74, 
    5555.098,
  5319.625, 5329.859, 5341.792, 5355.881, 5372.961, 5395.261, 5421.981, 
    5449.811, 5476.74, 5504.114, 5526.209, 5542.617, 5552.357, 5557.637, 
    5560.056,
  5266.047, 5278.92, 5288.533, 5298.713, 5306.675, 5313.591, 5316.041, 
    5318.034, 5319.972, 5323.182, 5330.02, 5341.613, 5355.23, 5369.658, 5384.3,
  5267.557, 5280.482, 5291.515, 5303.717, 5313.095, 5320.568, 5324.916, 
    5326.18, 5325.99, 5330.513, 5337.711, 5350.259, 5363.874, 5379.547, 
    5394.832,
  5267.414, 5279.264, 5293.084, 5306.955, 5318.073, 5328.539, 5330.912, 
    5332.137, 5333.003, 5336.849, 5345.302, 5357.495, 5373.334, 5389.187, 
    5406.329,
  5266.899, 5275.6, 5292.317, 5306.052, 5322.02, 5329.694, 5338.16, 5335.969, 
    5337.445, 5342.065, 5352.495, 5365.758, 5382.997, 5402.043, 5423.591,
  5265.997, 5271.859, 5288.975, 5305.292, 5322.662, 5336.672, 5341.896, 
    5342.662, 5344.891, 5348.913, 5360.91, 5374.864, 5394.573, 5413.375, 
    5439.604,
  5264.137, 5267.497, 5282.471, 5301.211, 5319.118, 5335.525, 5346.438, 
    5349.484, 5350.878, 5358.023, 5369.466, 5385.167, 5404.517, 5428.06, 
    5454.667,
  5260.84, 5264.266, 5276.868, 5296.403, 5316.358, 5335.993, 5348.606, 
    5354.566, 5359.708, 5365.931, 5378.211, 5395.128, 5415.048, 5438.091, 
    5465.533,
  5257.59, 5261.637, 5270.86, 5289.046, 5308.896, 5330.922, 5348.506, 
    5358.054, 5363.58, 5372.667, 5385.458, 5402.247, 5423.977, 5447.534, 
    5474.274,
  5254.709, 5260.125, 5268.471, 5284.555, 5303.938, 5326.502, 5345.818, 
    5358.887, 5368.574, 5377.904, 5390.924, 5408.042, 5428.95, 5452.46, 
    5477.618,
  5252.738, 5258.986, 5265.464, 5277.861, 5295.649, 5317.532, 5340.149, 
    5356.701, 5368.471, 5381.058, 5394.704, 5410.959, 5431.066, 5453.944, 
    5477.543,
  5315.11, 5305.102, 5296.673, 5290.034, 5282.746, 5276.529, 5273.621, 
    5278.057, 5288.293, 5301.558, 5317.27, 5335.545, 5353.518, 5370.298, 
    5387.093,
  5316.386, 5306.143, 5299.322, 5294.845, 5290.203, 5284.372, 5281.185, 
    5282.692, 5289.389, 5303.734, 5320.164, 5339.523, 5358.249, 5377.173, 
    5395.257,
  5314.812, 5305.37, 5299.357, 5296.13, 5293.706, 5291.028, 5286.496, 
    5287.333, 5294.051, 5304.95, 5321.521, 5341.313, 5361.592, 5379.846, 
    5400.049,
  5308.545, 5301.551, 5296.49, 5294.078, 5294.228, 5293.303, 5290.221, 
    5288.039, 5291.621, 5303.33, 5320.805, 5340.483, 5362.455, 5382.625, 
    5405.301,
  5297.498, 5293.989, 5290.899, 5289.62, 5291.249, 5293.444, 5292.755, 
    5289.767, 5293.519, 5301.607, 5318.707, 5337.851, 5360.853, 5380.226, 
    5404.683,
  5282.547, 5282.472, 5281.582, 5281.96, 5284.411, 5288.837, 5291.632, 
    5290.412, 5290.817, 5300.03, 5313.125, 5333.914, 5356.017, 5378.055, 
    5401.386,
  5265.353, 5268.775, 5269.842, 5271.857, 5275.326, 5281.321, 5286.404, 
    5289.06, 5289.715, 5295.269, 5307.595, 5327.072, 5348.475, 5371.033, 
    5393.526,
  5248.078, 5252.782, 5255.043, 5258.312, 5262.711, 5270.284, 5277.544, 
    5282.936, 5283.566, 5288.948, 5299.355, 5317.112, 5338.908, 5361.957, 
    5384.577,
  5230.706, 5236.289, 5240.538, 5243.718, 5248.211, 5256.474, 5265.475, 
    5273.77, 5278.261, 5281.491, 5290.077, 5306.157, 5326.317, 5349.349, 
    5371.682,
  5213.73, 5219.636, 5223.929, 5227.738, 5232.574, 5240.2, 5250.979, 
    5261.003, 5268.646, 5274.078, 5280.892, 5293.557, 5312.488, 5334.751, 
    5358.052,
  5292.804, 5293.843, 5291.066, 5281.473, 5269.601, 5261.586, 5267.482, 
    5283.483, 5300.159, 5311.08, 5319.597, 5326.917, 5337.375, 5349.74, 
    5363.941,
  5271.646, 5278.762, 5283.24, 5280.612, 5273.066, 5263.755, 5269.541, 
    5281.583, 5297.887, 5313.455, 5322.417, 5331.132, 5342.246, 5356.457, 
    5370.444,
  5248.181, 5261.614, 5272.478, 5277.269, 5273.951, 5270.307, 5267.346, 
    5282.214, 5296.663, 5310.869, 5322.502, 5331.778, 5344.171, 5357.964, 
    5374.042,
  5223.605, 5241.424, 5258.222, 5270.542, 5273.271, 5270.008, 5270.186, 
    5273.689, 5288.684, 5305.06, 5318.441, 5329.314, 5342.365, 5357.271, 
    5374.928,
  5199.188, 5220.884, 5242.029, 5261.943, 5271.124, 5272.38, 5270.337, 
    5273.564, 5283.64, 5295.431, 5311.097, 5323.337, 5337.171, 5351.141, 
    5369.95,
  5175.072, 5199.45, 5224.675, 5248.686, 5264.563, 5270.211, 5270.833, 
    5272.281, 5277.423, 5289.019, 5300.345, 5314.676, 5328.862, 5343.638, 
    5361.15,
  5153.899, 5181.171, 5209.324, 5236.54, 5256.955, 5268.207, 5270.815, 
    5273.671, 5278.222, 5282.678, 5291.566, 5303.025, 5316.86, 5332.238, 
    5347.796,
  5136.969, 5164.893, 5194.574, 5223.575, 5246.134, 5261.51, 5268.953, 
    5271.977, 5274.874, 5280.003, 5285.372, 5291.993, 5303.569, 5318.021, 
    5333.613,
  5125.116, 5153.555, 5184.333, 5213.907, 5237.42, 5253.978, 5263.562, 
    5269.84, 5273.451, 5276.237, 5279.509, 5284.533, 5290.289, 5302.093, 
    5315.891,
  5119.539, 5145.96, 5174.749, 5202.398, 5225.472, 5242.883, 5254.088, 
    5261.268, 5265.834, 5270.296, 5273.403, 5276.43, 5280.198, 5287.531, 
    5299.018,
  5167.016, 5161.914, 5160.405, 5163.83, 5169.875, 5173.607, 5183.064, 
    5197.787, 5209.045, 5212.517, 5219.128, 5226.534, 5234.539, 5240.672, 
    5249.209,
  5156.191, 5150.679, 5149.7, 5154.202, 5162.06, 5167.629, 5179.987, 
    5193.339, 5205.378, 5214.872, 5223.599, 5233.404, 5242.848, 5252.047, 
    5262.035,
  5146.132, 5140.618, 5141.152, 5146.53, 5158.076, 5166.164, 5174.533, 
    5194.889, 5208.222, 5217.061, 5228.009, 5239.207, 5251.073, 5261.287, 
    5272.44,
  5136.317, 5131.203, 5131.891, 5138.403, 5152.992, 5160.058, 5174.341, 
    5184.523, 5203.375, 5217.664, 5231.396, 5243.433, 5257.495, 5269.512, 
    5283.454,
  5126.777, 5122.985, 5123.496, 5133.373, 5147.937, 5162.785, 5166.44, 
    5185.328, 5203.505, 5217.7, 5233.02, 5246.786, 5261.36, 5274.41, 5288.933,
  5116.944, 5113.329, 5114.212, 5123.693, 5141.38, 5155.195, 5166.963, 
    5174.706, 5193.658, 5216.923, 5232.721, 5248.967, 5262.709, 5277.712, 
    5291.783,
  5105.68, 5103.664, 5106.798, 5116.973, 5136.133, 5153.822, 5162.127, 
    5175.845, 5193.98, 5212.195, 5231.905, 5247.91, 5262.782, 5276.328, 
    5290.26,
  5093.209, 5091.921, 5097.228, 5108.931, 5127.932, 5147.847, 5160.92, 
    5168.394, 5182.814, 5206.421, 5226.388, 5243.693, 5259.565, 5273.043, 
    5286.386,
  5080.514, 5080.129, 5090.712, 5104.916, 5126.029, 5145.149, 5158.11, 
    5169.256, 5181.671, 5199.471, 5219.408, 5238.38, 5253.468, 5266.625, 
    5278.697,
  5071.25, 5069.561, 5081.988, 5098.258, 5120.943, 5142.161, 5157.231, 
    5165.92, 5176.339, 5194.555, 5215.471, 5232.681, 5247.519, 5259.852, 
    5270.255,
  5120.631, 5111.266, 5102.017, 5094.027, 5086.611, 5081.461, 5079.477, 
    5082.503, 5090.765, 5097.025, 5102.496, 5106.153, 5108.553, 5111.517, 
    5118.575,
  5114.728, 5103.945, 5095.146, 5087.284, 5080.731, 5076.784, 5075.572, 
    5077.145, 5085.056, 5094.032, 5099.682, 5103.618, 5105.949, 5108.998, 
    5116.424,
  5107.222, 5095.72, 5088.024, 5081.292, 5076.341, 5073.878, 5071.477, 
    5076.88, 5085.618, 5091.938, 5098.212, 5102.254, 5104.611, 5108.761, 
    5116.308,
  5096.622, 5086.12, 5079.254, 5074.095, 5071.953, 5069.818, 5071.128, 
    5071.368, 5081.736, 5089.793, 5097.773, 5101.417, 5105.374, 5110.352, 
    5120.288,
  5083.747, 5074.168, 5069.658, 5067.655, 5067.794, 5070.122, 5069.066, 
    5073.753, 5082.917, 5090.096, 5098.177, 5103.007, 5108.51, 5114.704, 
    5126.04,
  5068.66, 5060.645, 5057.737, 5058.301, 5060.118, 5064.673, 5067.797, 
    5070.899, 5079.699, 5091.904, 5100.144, 5106.575, 5113.21, 5122.689, 
    5134.433,
  5053.681, 5047.378, 5047.056, 5050.304, 5053.95, 5060.879, 5063.573, 
    5072.299, 5083.586, 5093.933, 5103.77, 5111.584, 5120.532, 5131.469, 
    5144.001,
  5041.194, 5035.311, 5035.488, 5041.99, 5046.655, 5055.939, 5061.714, 
    5068.885, 5081.357, 5095.521, 5106.795, 5117.399, 5128.736, 5141.142, 
    5155.088,
  5031.869, 5025.542, 5027.749, 5037.106, 5043.467, 5053.294, 5060.348, 
    5071.195, 5084.748, 5097.437, 5110.759, 5123.693, 5136.625, 5150.298, 
    5164.578,
  5026.285, 5017.734, 5023.104, 5032.618, 5039.347, 5051.131, 5060.253, 
    5069.147, 5083.426, 5099.283, 5114.627, 5128.856, 5143.628, 5158.505, 
    5173.359,
  5088.929, 5084.696, 5079.434, 5072.782, 5068.599, 5063.489, 5057.007, 
    5051.805, 5048.183, 5045.645, 5050.028, 5056.357, 5061.39, 5066.655, 
    5075.825,
  5071.022, 5066.466, 5063.085, 5056.914, 5054.698, 5049.742, 5048.78, 
    5042.288, 5039.011, 5040.17, 5044.633, 5052.438, 5058.555, 5064.313, 
    5072.37,
  5054.66, 5049.335, 5045.866, 5042.383, 5040.996, 5042.072, 5034.31, 
    5036.557, 5031.837, 5033.01, 5038.819, 5047.26, 5054.133, 5060.855, 
    5067.91,
  5037.585, 5031.555, 5028.173, 5026.96, 5027.565, 5027.722, 5031.257, 
    5022.536, 5025.347, 5026.27, 5032.969, 5040.438, 5048.801, 5055.418, 
    5063.881,
  5018.294, 5011.857, 5010.724, 5013.219, 5017.323, 5022.11, 5020.229, 
    5022.348, 5018.123, 5021.413, 5027.474, 5034.693, 5042.753, 5048.938, 
    5058.175,
  4996.848, 4989.711, 4992.167, 4999.695, 5006.082, 5011.399, 5015.91, 
    5014.562, 5015.573, 5019.312, 5022.89, 5029.972, 5036.118, 5043.089, 
    5051.72,
  4973.886, 4967.954, 4972.411, 4986.688, 4997.121, 5004.528, 5007.082, 
    5010.73, 5012.638, 5014.98, 5020.374, 5024.813, 5030.553, 5036.848, 
    5045.53,
  4959.478, 4957.303, 4964.509, 4979.318, 4989.455, 4997.699, 5001.839, 
    5004.041, 5007.186, 5012.198, 5015.885, 5019.977, 5025.624, 5031.96, 
    5041.436,
  4956.414, 4958.098, 4966.094, 4980.459, 4987.599, 4994.316, 4997.796, 
    5001.667, 5005.864, 5010.266, 5013.403, 5017.482, 5022.647, 5029.486, 
    5039.58,
  4960.883, 4963.455, 4972.548, 4982.541, 4987.175, 4993.793, 4996.528, 
    5000.243, 5006.171, 5011.543, 5013.239, 5017.073, 5023.116, 5030.83, 
    5041.985,
  5076.95, 5075.854, 5075.317, 5074.65, 5074.686, 5073.528, 5072.964, 
    5073.444, 5073.117, 5068.408, 5063.33, 5057.373, 5052.721, 5046.865, 
    5044.544,
  5061.723, 5058.688, 5057.326, 5055.68, 5055.002, 5054.448, 5056.201, 
    5054.765, 5055.2, 5056.177, 5052.046, 5048.536, 5044.815, 5042.31, 
    5040.804,
  5042.623, 5039.188, 5036.783, 5036.802, 5036.431, 5038.977, 5035.554, 
    5043.005, 5042.261, 5041.912, 5040.402, 5038.898, 5037.579, 5036.419, 
    5037.445,
  5021.683, 5018.449, 5017.747, 5018.354, 5020.036, 5021.806, 5027.029, 
    5021.835, 5029.529, 5030.361, 5030.577, 5028.762, 5031.114, 5031.426, 
    5035.808,
  4994.168, 4991.959, 4993.614, 4998.267, 5003.174, 5008.281, 5011.067, 
    5017.286, 5015.236, 5016.542, 5019.634, 5019.246, 5024.348, 5026.596, 
    5033.696,
  4971.346, 4969.044, 4971.399, 4978.526, 4987.51, 4995.513, 5001.981, 
    5003.187, 5007.285, 5010.493, 5010.802, 5013.129, 5018.329, 5024.125, 
    5031.51,
  4956.561, 4952.651, 4958.044, 4963.328, 4976.984, 4989.753, 4994.515, 
    4999.254, 4999.904, 5001.419, 5004.625, 5007.766, 5013.816, 5021.719, 
    5030.123,
  4954.983, 4950.01, 4955.121, 4959.153, 4973.29, 4987.836, 4992.892, 
    4992.528, 4992.476, 4996.172, 4998.17, 5002.935, 5010.438, 5019.963, 
    5029.61,
  4969.387, 4963.819, 4963.69, 4966.997, 4978.727, 4988.772, 4989.843, 
    4990.537, 4988.652, 4989.771, 4992.939, 4999.366, 5007.158, 5018.076, 
    5028.57,
  4978.798, 4974.665, 4974.474, 4977.106, 4982.198, 4986.666, 4986.056, 
    4983.813, 4982.514, 4985.991, 4989.743, 4995.733, 5004.363, 5015.863, 
    5027.585,
  5100.354, 5099.584, 5100.279, 5101.729, 5106.011, 5109.836, 5114.629, 
    5120.433, 5124.212, 5124.861, 5125.893, 5126.113, 5124.057, 5120.688, 
    5115.611,
  5079.938, 5079.788, 5082.914, 5086.222, 5089.196, 5093.654, 5099.239, 
    5100.411, 5103.824, 5108.664, 5108.201, 5109.14, 5107.129, 5105.252, 
    5099.139,
  5054.524, 5053.325, 5055.926, 5062.882, 5069.504, 5078.682, 5077.514, 
    5088.479, 5085.807, 5088.417, 5090.087, 5091.663, 5090.823, 5088.792, 
    5085.437,
  5034.188, 5028.625, 5030.017, 5034.338, 5044.358, 5050.962, 5065.508, 
    5060.344, 5071.298, 5072.877, 5075.022, 5075.347, 5076.336, 5075.094, 
    5072.191,
  5020.375, 5009.763, 5008.364, 5012.939, 5019.805, 5030.023, 5033.629, 
    5046.994, 5046.989, 5050.357, 5056.109, 5057.525, 5060.148, 5059.83, 
    5060.764,
  5013.727, 4999.768, 4994.874, 4997.584, 5002.323, 5008.082, 5016.706, 
    5019.394, 5028.232, 5035.652, 5038.344, 5042.092, 5045.794, 5048.192, 
    5050.202,
  5013.844, 4998.553, 4994.144, 4996.473, 4996.85, 4997.438, 5000.942, 
    5007.707, 5012.616, 5016.086, 5022.711, 5027.291, 5033.003, 5036.893, 
    5041.006,
  5019.212, 5002.743, 4991.275, 4986.277, 4985.427, 4990.072, 4993.552, 
    4996.073, 4999.423, 5005.483, 5010.664, 5016.958, 5023.245, 5028.406, 
    5033.722,
  5025.912, 5009.738, 4998.929, 4993.755, 4993.998, 4996.341, 4996.883, 
    4998.176, 4996.717, 4998.745, 5003.242, 5009.572, 5014.857, 5021.824, 
    5028.451,
  5034.897, 5018.513, 5005.983, 5001.292, 4999.439, 5000.465, 4998.735, 
    4995.57, 4992.862, 4994.843, 4998.02, 5003.552, 5009.305, 5017.834, 
    5025.604,
  5125.722, 5117.797, 5111.668, 5108.459, 5108.258, 5110.023, 5113.647, 
    5121.172, 5128.792, 5135.788, 5144.067, 5152.825, 5159.833, 5166.532, 
    5171.156,
  5115.079, 5103.31, 5091.895, 5085.634, 5083.325, 5086.282, 5092.509, 
    5097.057, 5104.675, 5115.406, 5122.464, 5131.939, 5139.174, 5148.129, 
    5152.182,
  5108.447, 5092.419, 5077.167, 5068.074, 5062.945, 5068.891, 5068.133, 
    5082.475, 5087.203, 5096.47, 5105.375, 5115.015, 5123.184, 5130.967, 
    5138.404,
  5101.512, 5082.447, 5066.301, 5054.508, 5050.048, 5047.042, 5059.477, 
    5058.403, 5073.999, 5083.973, 5094.208, 5102.317, 5111.807, 5120.041, 
    5126.852,
  5097.292, 5077.272, 5059.019, 5049.283, 5042.269, 5042.016, 5040.53, 
    5052.271, 5060.676, 5071.162, 5084.431, 5092.95, 5102.426, 5109.622, 
    5117.902,
  5094.398, 5074.299, 5056.145, 5044.597, 5036.792, 5034.112, 5035.575, 
    5036.29, 5045.668, 5061.583, 5072.423, 5084.619, 5093.771, 5102.865, 
    5110.141,
  5093.811, 5075.589, 5056.569, 5043.159, 5033.666, 5029.244, 5027.303, 
    5031.781, 5037.367, 5047.022, 5061.012, 5073.312, 5083.617, 5093.835, 
    5101.823,
  5094.181, 5076.896, 5057.554, 5041.75, 5028.997, 5022.525, 5020.317, 
    5019.783, 5023.972, 5034.795, 5047.14, 5059.668, 5072.918, 5084.799, 
    5093.683,
  5096.555, 5081.59, 5063.417, 5045.786, 5032.06, 5022.55, 5018.029, 
    5017.177, 5016.853, 5022.09, 5033.908, 5048.107, 5062.098, 5075.523, 
    5085.718,
  5098.792, 5084.155, 5066.617, 5048.86, 5031.66, 5020.556, 5017.009, 
    5014.624, 5013.461, 5016.57, 5025.661, 5038.73, 5053.618, 5068.055, 
    5079.489,
  5184.299, 5168.317, 5151.971, 5136.222, 5123.608, 5114.601, 5108.626, 
    5108.255, 5110.004, 5114.175, 5122.533, 5132.308, 5142.793, 5153.675, 
    5165.382,
  5181.928, 5163.775, 5145.43, 5127.885, 5113.475, 5101.583, 5096.912, 
    5090.444, 5090.77, 5095.424, 5101.337, 5112.323, 5122.027, 5134.328, 
    5142.701,
  5179.973, 5161.916, 5142.594, 5124.912, 5107.504, 5098.082, 5083.954, 
    5083.068, 5076.444, 5076.629, 5080.67, 5089.768, 5101.04, 5112.342, 
    5123.221,
  5178.342, 5160.767, 5142.888, 5124.007, 5106.617, 5091.058, 5084.074, 
    5070.202, 5067.719, 5065.351, 5066.12, 5072.048, 5081.545, 5094.025, 
    5104.955,
  5176.562, 5161.771, 5145.758, 5127.116, 5109.04, 5092.65, 5077.563, 
    5070.269, 5060.991, 5056.201, 5057.158, 5060.228, 5068.206, 5077.034, 
    5089.693,
  5175.259, 5163.27, 5148.498, 5130.927, 5110.94, 5093.117, 5077.667, 
    5063.186, 5054.19, 5050.602, 5050.909, 5055.131, 5061.625, 5069.585, 
    5080.477,
  5174.513, 5166.882, 5153.071, 5135.44, 5115.248, 5094.461, 5076.285, 
    5062.667, 5051.224, 5044.606, 5046.959, 5052.709, 5059.591, 5067.116, 
    5077.6,
  5176.395, 5168.82, 5154.59, 5137.531, 5115.329, 5094.142, 5074.979, 
    5058.087, 5045.588, 5040.01, 5043.06, 5051.731, 5059.934, 5068.552, 
    5079.693,
  5178.653, 5170.867, 5156.572, 5136.746, 5113.899, 5092.012, 5071.792, 5056, 
    5043.097, 5035.613, 5039.577, 5050.754, 5060.8, 5071.876, 5083.353,
  5181.353, 5168.173, 5150.66, 5129.621, 5105.924, 5085.091, 5066.343, 
    5048.903, 5037.091, 5031.061, 5035.994, 5049.161, 5062.251, 5075.827, 
    5086.946,
  5259.777, 5250.472, 5245.604, 5236.17, 5224.272, 5208.981, 5189.2, 
    5174.134, 5157.215, 5135.962, 5120.919, 5108.889, 5100.728, 5095.964, 
    5095.747,
  5258.22, 5252.359, 5247.334, 5237.155, 5223.109, 5203.147, 5190.41, 
    5161.955, 5141.872, 5127.601, 5110.115, 5097.576, 5088.78, 5086.248, 
    5085.244,
  5259.867, 5256.716, 5250.007, 5239.727, 5219.418, 5205.418, 5171.182, 
    5165.728, 5135.802, 5114.921, 5098.204, 5086.205, 5076.996, 5074.816, 
    5077.324,
  5263.501, 5259.422, 5251.534, 5236.451, 5216.924, 5190.941, 5172.312, 
    5132.8, 5119.832, 5101.838, 5086.108, 5073.602, 5066.183, 5063.843, 
    5068.669,
  5268.409, 5262.888, 5253.053, 5234.454, 5211.51, 5183.039, 5151.568, 
    5132.901, 5108.729, 5085.6, 5073.791, 5061.218, 5055.721, 5051.863, 
    5059.299,
  5273.339, 5265.887, 5251.297, 5229.256, 5199.239, 5167.065, 5135.039, 
    5106.021, 5086.3, 5073.733, 5060.5, 5051.551, 5046.202, 5043.572, 5048.718,
  5279.43, 5270.221, 5251.207, 5224.757, 5191.445, 5152.514, 5117.732, 
    5094.702, 5076.438, 5061.122, 5051.364, 5044.01, 5039.992, 5038.554, 
    5041.459,
  5286.12, 5271.718, 5248.826, 5219.323, 5179.461, 5139.834, 5102.747, 
    5076.208, 5060.58, 5052.51, 5044.037, 5038.167, 5036.541, 5036.291, 
    5038.639,
  5290.996, 5274.985, 5251.77, 5217.932, 5176.906, 5133.229, 5094.314, 
    5069.537, 5054.909, 5046, 5038.517, 5034.436, 5034.136, 5034.352, 5037.571,
  5295.632, 5275.861, 5249.011, 5213.736, 5170.94, 5127.734, 5089.229, 
    5059.978, 5045.739, 5041.083, 5034.44, 5032.105, 5033.217, 5035.202, 
    5039.409,
  5338.474, 5333.484, 5326.592, 5307.413, 5280.249, 5245.187, 5203.405, 
    5173.65, 5151.187, 5129.483, 5116.438, 5108.652, 5103.664, 5101.027, 
    5100.669,
  5340.541, 5339.309, 5327.779, 5304.542, 5273.26, 5227.386, 5192.047, 
    5146.794, 5120.932, 5107.901, 5097.75, 5092.893, 5089.188, 5089.177, 
    5087.601,
  5348.604, 5345.146, 5330.134, 5307.675, 5268.887, 5230.776, 5168.706, 
    5143.478, 5114.583, 5097.396, 5087.084, 5084.665, 5080.932, 5080.37, 
    5078.485,
  5356.327, 5350.316, 5335.491, 5308.692, 5273.867, 5222.467, 5179.667, 
    5130.218, 5104.767, 5092.942, 5083.38, 5077.042, 5073.149, 5070.731, 
    5069.425,
  5364.415, 5356.718, 5341.432, 5315.884, 5281.168, 5234.87, 5180.116, 
    5143.725, 5118.657, 5093.044, 5082.492, 5072.16, 5068.177, 5063.745, 
    5062.793,
  5371.086, 5363.438, 5346.66, 5323.238, 5288.533, 5245.495, 5198.775, 
    5151.789, 5120.765, 5101.515, 5085.087, 5073.69, 5066.68, 5061.421, 
    5058.762,
  5377.924, 5370.534, 5353.836, 5331.977, 5301.306, 5261.918, 5215.373, 
    5174.084, 5142.187, 5114.6, 5093.7, 5078.689, 5067.891, 5061.546, 5057.933,
  5384.884, 5376.434, 5360.667, 5339.562, 5309.894, 5275.012, 5235.744, 
    5191.017, 5154.884, 5128.057, 5104.864, 5085.795, 5072.444, 5064.729, 
    5061.66,
  5391.721, 5383.375, 5368.462, 5348.504, 5323.258, 5289.914, 5252.138, 
    5213.69, 5175.915, 5144.063, 5116.438, 5095.144, 5078.415, 5068.895, 
    5066.51,
  5396.308, 5387.213, 5374.254, 5355.427, 5329.307, 5299.145, 5265.853, 
    5227.463, 5189.579, 5157.286, 5129.304, 5105.208, 5086.042, 5073.516, 
    5071.403,
  5375.866, 5381.691, 5380.299, 5369.069, 5349.762, 5320.814, 5280.719, 
    5243.806, 5205.633, 5159.906, 5123.705, 5097.753, 5084.477, 5071.914, 
    5064.718,
  5383.135, 5388.782, 5386.651, 5377.186, 5360.035, 5330.22, 5302.663, 
    5256.349, 5215.071, 5178.188, 5139.08, 5108.422, 5090.63, 5081.557, 
    5073.642,
  5391.178, 5396.996, 5393.572, 5387.04, 5367.166, 5351.537, 5309.614, 
    5286.105, 5247.537, 5201.977, 5159.918, 5124.614, 5099.965, 5090.988, 
    5085.314,
  5399.917, 5403.598, 5402.37, 5393.313, 5381.644, 5354.971, 5336.443, 
    5297.405, 5259.074, 5223.985, 5182.899, 5144.888, 5114.438, 5098.059, 
    5093.998,
  5408.195, 5410.905, 5410.667, 5402.245, 5390.72, 5371.806, 5345.81, 
    5317.637, 5290.887, 5245.912, 5207.391, 5166.782, 5134.309, 5109.846, 
    5100.778,
  5415.235, 5419.21, 5417.497, 5411.308, 5397.886, 5379.287, 5359.232, 
    5330.109, 5297.093, 5266.78, 5230.646, 5190.406, 5155.017, 5126.176, 
    5110.791,
  5421.641, 5425.464, 5423.565, 5417.065, 5405.484, 5389.501, 5367.07, 
    5344.954, 5318.975, 5284.664, 5248.726, 5212.934, 5175.918, 5145.55, 
    5124.135,
  5426.075, 5429.092, 5427.489, 5421.471, 5408.69, 5393.215, 5374.68, 
    5350.491, 5322.615, 5295.624, 5264.256, 5229.903, 5195.407, 5162.696, 
    5139.615,
  5427.322, 5430.026, 5427.9, 5421.071, 5411.3, 5396.745, 5377.176, 5356.671, 
    5332.987, 5304.008, 5274.058, 5242.021, 5210.634, 5178.119, 5153.277,
  5424.265, 5425.65, 5424.45, 5418.813, 5406.823, 5391.959, 5374.296, 
    5351.877, 5327.973, 5304.337, 5278.03, 5248.951, 5219.309, 5189.664, 
    5163.714,
  5423.144, 5437.361, 5446.691, 5447.655, 5441.532, 5428.567, 5406.219, 
    5380.248, 5345.682, 5300.563, 5255.206, 5210.509, 5178.315, 5159.667, 
    5152.984,
  5423.698, 5439.086, 5448.154, 5449.993, 5445.507, 5432.71, 5418.354, 
    5388.472, 5355.995, 5322.413, 5282.808, 5242.71, 5205.289, 5185.17, 
    5174.906,
  5426.854, 5443.121, 5450.569, 5454.535, 5448.015, 5443.076, 5420.385, 
    5405.696, 5378.288, 5343.645, 5307.353, 5271.83, 5236.756, 5209.215, 
    5196.295,
  5432.209, 5446.289, 5454.32, 5455.835, 5452.82, 5441.915, 5431.729, 
    5408.938, 5382.231, 5359.114, 5327.165, 5295.507, 5264.209, 5235.198, 
    5216.841,
  5438.228, 5449.522, 5457.026, 5457.944, 5455.186, 5447.226, 5433.293, 
    5417.863, 5399.292, 5367.836, 5342.213, 5312.665, 5285.125, 5258.504, 
    5235.137,
  5442.683, 5451.844, 5456.931, 5457.934, 5453.4, 5445.005, 5433.633, 
    5414.613, 5393.361, 5372.792, 5348.981, 5323.05, 5298.187, 5273.837, 
    5252.517,
  5445.994, 5453.217, 5455.313, 5454.357, 5449.686, 5441.21, 5427.523, 
    5412.823, 5393.933, 5370.812, 5348.383, 5325.896, 5303.003, 5280.973, 
    5261.542,
  5447.698, 5451.003, 5450.417, 5447.982, 5440.213, 5430.162, 5416.767, 
    5399.395, 5380.355, 5361.993, 5341.677, 5320.599, 5300.024, 5280.385, 
    5263.358,
  5446.881, 5447.22, 5443.341, 5436.461, 5428, 5415.951, 5401.102, 5385.865, 
    5368.165, 5347.996, 5327.889, 5308.479, 5289.538, 5272.026, 5257.2,
  5442.322, 5437.282, 5430.582, 5422.033, 5409.269, 5394.877, 5380.18, 
    5362.539, 5344.964, 5327.931, 5309.364, 5290.54, 5273.059, 5257.657, 
    5245.05,
  5465.753, 5482.748, 5494.926, 5498.979, 5498.833, 5492.716, 5479.396, 
    5465.587, 5446.812, 5423.677, 5403.208, 5384.017, 5365.799, 5352.416, 
    5344.86,
  5473.21, 5489.752, 5500.086, 5504.989, 5504.279, 5497.042, 5488.245, 
    5469.708, 5452.171, 5435.875, 5415.348, 5396.19, 5376.832, 5360.41, 
    5347.087,
  5483.512, 5498.724, 5506.122, 5511.105, 5507.774, 5505.433, 5490.557, 
    5481.102, 5462.094, 5441.441, 5422.617, 5403.791, 5383.811, 5365.723, 
    5348.693,
  5493.903, 5505.37, 5513.012, 5514.817, 5513.795, 5502.818, 5496.143, 
    5477.219, 5461.046, 5444.836, 5423.561, 5405.504, 5385.307, 5367.117, 
    5348.126,
  5503.324, 5513.108, 5518.616, 5519.112, 5515.081, 5508.771, 5493.55, 
    5480.451, 5463.301, 5441.426, 5422.664, 5401.105, 5382.615, 5361.537, 
    5342.916,
  5510.885, 5518.87, 5521.29, 5521.111, 5514.528, 5504.074, 5491.918, 
    5473.853, 5454.558, 5435.648, 5415.283, 5393.228, 5373.023, 5351.742, 
    5331.787,
  5519.458, 5525.018, 5524.206, 5519.912, 5511.601, 5500.248, 5484.111, 
    5467.135, 5446.756, 5424.9, 5402.803, 5380.375, 5357.62, 5335.388, 
    5313.935,
  5526.258, 5526.866, 5523.117, 5516.534, 5504.188, 5489.787, 5472.782, 
    5453.354, 5431.429, 5409.535, 5385.813, 5361.686, 5337.435, 5313.794, 
    5291.088,
  5531.906, 5529.312, 5521.224, 5509.215, 5494.957, 5477.35, 5457.158, 
    5437.109, 5413.773, 5388.689, 5363.377, 5337.62, 5311.348, 5286.137, 
    5261.898,
  5531.69, 5522.692, 5511.431, 5498.745, 5480.064, 5459.172, 5437.06, 
    5411.828, 5387.042, 5361.963, 5335.368, 5307.507, 5279.5, 5253.507, 
    5228.207,
  5522.199, 5537.662, 5552.486, 5562.635, 5570.654, 5575.654, 5578.098, 
    5577.662, 5572.53, 5560.517, 5547.333, 5531.355, 5511.355, 5487.393, 
    5463.615,
  5514.332, 5533.665, 5552.437, 5566.089, 5575.141, 5579.453, 5580.354, 
    5576.144, 5570.471, 5562.486, 5546.156, 5526.125, 5503.285, 5477.667, 
    5449.536,
  5505.579, 5528.972, 5549.92, 5566.373, 5574.853, 5581.566, 5580.667, 
    5579.478, 5567.194, 5551.148, 5534.725, 5515.885, 5489.382, 5461.252, 
    5428.979,
  5497.282, 5522.042, 5546.068, 5562.919, 5575.382, 5575.866, 5576.859, 
    5567.555, 5561.686, 5548.628, 5522.563, 5499.749, 5471.675, 5439.912, 
    5402.37,
  5489.678, 5515.375, 5540.625, 5558.495, 5569.576, 5574.12, 5570.359, 
    5562.995, 5548.457, 5526.167, 5507.829, 5476.433, 5446.524, 5408.527, 
    5369.317,
  5484.307, 5509.756, 5533.785, 5552.797, 5562.677, 5563.494, 5557.622, 
    5544.128, 5528.934, 5508.729, 5481.069, 5447.091, 5411.016, 5368.424, 
    5325.768,
  5482.907, 5507.765, 5529.03, 5545.131, 5552.885, 5552.012, 5543.394, 
    5528.825, 5506.558, 5478.526, 5447.171, 5409.169, 5365.367, 5318.984, 
    5269.486,
  5485.332, 5506.317, 5524.27, 5537.3, 5540.107, 5535.521, 5522.25, 5503.393, 
    5478.952, 5448.089, 5408.895, 5362.846, 5314.011, 5261.356, 5208.376,
  5489.636, 5507.461, 5520.748, 5526.463, 5526.099, 5516.853, 5499.771, 
    5476.442, 5444.016, 5404.393, 5358.324, 5308.208, 5254.021, 5197.185, 
    5147.023,
  5493.355, 5505.06, 5512.525, 5515.638, 5507.521, 5492.2, 5469.26, 5436.997, 
    5399.04, 5353.358, 5302.866, 5246.935, 5187.887, 5135.156, 5089.808,
  5516.728, 5514.63, 5510.786, 5506.859, 5506.73, 5509.365, 5516.027, 
    5524.736, 5531.662, 5535.065, 5536.718, 5532.82, 5521.363, 5503.814, 
    5479.319,
  5501.769, 5502.256, 5501.561, 5500.29, 5500.875, 5503.044, 5508.832, 
    5512.346, 5518.674, 5523.497, 5519.812, 5513.448, 5500.408, 5482.305, 
    5454.708,
  5483.593, 5486.835, 5488.325, 5490.552, 5491.703, 5496.37, 5496.937, 
    5506.444, 5502.923, 5503.297, 5500.915, 5492.782, 5476.585, 5455.282, 
    5426.937,
  5462.044, 5467.64, 5471.482, 5474.141, 5478.435, 5479.511, 5486.888, 
    5482.126, 5489.636, 5485.6, 5477.608, 5468.266, 5450.809, 5427.594, 
    5395.218,
  5438.367, 5444.344, 5449.102, 5454.378, 5458.316, 5464.43, 5463.312, 
    5473.666, 5463.507, 5461.547, 5454.745, 5440.904, 5423.342, 5396.255, 
    5363.815,
  5413.074, 5418.073, 5422.199, 5427.502, 5431.699, 5437.168, 5441.677, 
    5438.483, 5441.091, 5435.591, 5423.875, 5409.889, 5390.029, 5362.601, 
    5330.555,
  5386.708, 5390.161, 5392.817, 5397.335, 5403.192, 5407.834, 5411.029, 
    5414.43, 5409.079, 5400.636, 5392.042, 5375.373, 5353.218, 5324.981, 
    5292.547,
  5360.461, 5361.455, 5361.995, 5365.579, 5369.326, 5375.732, 5378.87, 
    5377.812, 5375.227, 5369.46, 5356.398, 5339.209, 5316.607, 5288.298, 
    5255.189,
  5337.388, 5336.707, 5336.347, 5338.783, 5341.878, 5344.771, 5347.106, 
    5348.467, 5344.61, 5336.999, 5325.958, 5308.689, 5284.16, 5254.453, 
    5219.261,
  5318.851, 5316.443, 5317.246, 5319.876, 5322.253, 5326.595, 5330.427, 
    5330.652, 5327.734, 5319.509, 5303.74, 5280.884, 5252.492, 5219.538, 
    5181.205,
  5506.228, 5481.876, 5460.354, 5442.147, 5427.611, 5415.068, 5404.516, 
    5398.608, 5392.194, 5385.144, 5381.569, 5378.271, 5373.736, 5366.864, 
    5357.947,
  5475.431, 5451.258, 5432.811, 5416.272, 5403.247, 5392.603, 5388.96, 
    5380.286, 5378.044, 5376.358, 5370.875, 5366.601, 5359.642, 5351.515, 
    5338.71,
  5446.493, 5425.731, 5408.986, 5395.947, 5383.922, 5379.255, 5369.292, 
    5373.348, 5365.29, 5362.684, 5357.903, 5352.322, 5342.659, 5331.691, 
    5317.998,
  5422.314, 5404.605, 5389.826, 5377.773, 5368.886, 5360.562, 5360.909, 
    5351.41, 5353.64, 5349.092, 5342.967, 5335.487, 5324.626, 5312.018, 
    5294.959,
  5404.769, 5388.725, 5374.605, 5364.104, 5356.038, 5350.851, 5343.254, 
    5345.025, 5336.977, 5331.95, 5326.501, 5316.243, 5305.192, 5289.052, 
    5270.489,
  5390.192, 5374.978, 5360.948, 5350.852, 5341.298, 5335.592, 5331.326, 
    5324.313, 5321.311, 5316.853, 5307.896, 5297.466, 5284.909, 5265.835, 
    5241.847,
  5378.214, 5363.87, 5349.416, 5338.288, 5329.464, 5322.495, 5316.809, 
    5313.766, 5307.139, 5299.295, 5291.708, 5280.772, 5263.751, 5239.178, 
    5208.554,
  5367.392, 5352.76, 5337.939, 5326.818, 5316.208, 5310.316, 5304.879, 
    5298.847, 5293.4, 5288.009, 5278.556, 5262.833, 5239.534, 5208.394, 
    5171.18,
  5357.26, 5343.309, 5329.007, 5317.792, 5309.307, 5302.753, 5295.923, 
    5291.053, 5285.675, 5276.326, 5261.953, 5239.457, 5208.548, 5170.565, 
    5127.758,
  5347.652, 5332.768, 5318.987, 5309.836, 5300.195, 5293.378, 5289.223, 
    5283.241, 5275.062, 5260.494, 5238.719, 5208.314, 5170.683, 5127.874, 
    5080.961,
  5571.661, 5544.717, 5517.583, 5492.14, 5468.352, 5443.679, 5415.108, 
    5393.268, 5371.391, 5345.272, 5327.481, 5313.37, 5302.556, 5292.617, 
    5285.143,
  5556.394, 5530.631, 5506.82, 5483.531, 5461.44, 5433.423, 5415.058, 
    5379.79, 5357.544, 5341.391, 5322.853, 5307.661, 5294.952, 5284.118, 
    5272.812,
  5542.342, 5520.661, 5499.309, 5479.766, 5454.965, 5436.905, 5400.946, 
    5390.13, 5359.434, 5335.439, 5316.225, 5300.654, 5284.562, 5271.41, 
    5258.003,
  5529.6, 5510.826, 5492.448, 5472.65, 5451.222, 5424.236, 5405.238, 5368.73, 
    5349.182, 5330.88, 5308.166, 5290.722, 5273.369, 5257.558, 5240.117,
  5519.269, 5503.621, 5488.11, 5469.027, 5448.113, 5423.497, 5395.107, 
    5374.371, 5348.268, 5318.819, 5300.394, 5277.757, 5260.479, 5239.125, 
    5220.886,
  5509.387, 5495.906, 5481.119, 5463.831, 5441.063, 5416.723, 5391.229, 
    5360.486, 5334.23, 5311.634, 5287.942, 5264.395, 5243.89, 5219.357, 
    5195.599,
  5500.562, 5490.216, 5476.462, 5458.498, 5436.512, 5411.178, 5382.959, 
    5356.761, 5328.56, 5299.756, 5274.374, 5249.148, 5223.283, 5195.491, 
    5165.466,
  5492.714, 5482.332, 5467.51, 5449.779, 5425.139, 5399.823, 5371.376, 
    5340.734, 5311.898, 5285.948, 5258.161, 5229.617, 5200.086, 5166.912, 
    5130.91,
  5485.719, 5476.076, 5460.363, 5439.781, 5415.314, 5387.168, 5355.697, 
    5327.328, 5298.347, 5267.871, 5237.908, 5206.413, 5171.407, 5133.151, 
    5091.284,
  5477.358, 5463.275, 5445.063, 5424.228, 5396.244, 5366.437, 5335.67, 
    5304.551, 5274.726, 5246.251, 5213.946, 5178.003, 5139.126, 5095.32, 
    5052.383,
  5590.833, 5583.125, 5574.046, 5567.603, 5563.003, 5553.458, 5541.217, 
    5528.753, 5509.945, 5480.666, 5453.624, 5424.586, 5395.03, 5361.152, 
    5329.357,
  5580.264, 5573.269, 5565.105, 5559.544, 5553.311, 5544.248, 5535.724, 
    5512.144, 5493.062, 5473.849, 5446.658, 5416.686, 5384.272, 5350.776, 
    5313.164,
  5567.623, 5561.004, 5553.596, 5548.956, 5540.798, 5534.45, 5517.54, 
    5517.747, 5489.265, 5460.119, 5433.589, 5406.187, 5371.027, 5334.004, 
    5293.229,
  5551.177, 5544.938, 5538.757, 5533.375, 5526.433, 5516.491, 5508.332, 
    5483.337, 5472.125, 5452.59, 5420.61, 5390.686, 5355.361, 5315.535, 
    5270.487,
  5532.454, 5526.457, 5520.987, 5515.914, 5509.36, 5500.564, 5487.715, 
    5477.506, 5455.293, 5427.001, 5403.96, 5369.942, 5334.878, 5291.297, 
    5245.173,
  5510.779, 5505.904, 5500.141, 5496.571, 5489.853, 5482.145, 5469.83, 
    5449.898, 5431.646, 5410.436, 5381.755, 5347.851, 5309.854, 5264.993, 
    5216.166,
  5489.335, 5485.786, 5480.441, 5476.459, 5470.899, 5462.21, 5449.309, 
    5433.882, 5411.349, 5385.363, 5357.781, 5323.322, 5281.897, 5234.995, 
    5183.79,
  5468.341, 5464.374, 5459.426, 5456.389, 5449.935, 5441.552, 5427.25, 
    5408.247, 5387.51, 5364.652, 5333.775, 5296.231, 5253.478, 5205.23, 
    5151.854,
  5447.01, 5444.536, 5439.959, 5434.853, 5427.977, 5417.865, 5402.96, 
    5386.878, 5365.229, 5338.321, 5305.886, 5267.65, 5223.297, 5172.355, 
    5120.011,
  5423.532, 5418.789, 5414.273, 5410.575, 5403.257, 5392.247, 5377.078, 
    5358.001, 5336.499, 5310.925, 5277.375, 5237.419, 5191.823, 5141.02, 
    5090.627,
  5517.455, 5512.293, 5507.888, 5499.82, 5493.542, 5484.724, 5474.166, 
    5465.418, 5453.586, 5435.125, 5418.304, 5400.216, 5379.392, 5355.873, 
    5331.572,
  5490.237, 5484.247, 5480.406, 5472.72, 5465.461, 5457.898, 5453.34, 
    5434.425, 5422.632, 5413.38, 5395.191, 5377.716, 5357.318, 5337.345, 
    5311.766,
  5460.555, 5454.334, 5449.334, 5442.982, 5435.785, 5431.896, 5416.41, 
    5421.586, 5397.627, 5384.499, 5370.058, 5355.805, 5335.327, 5314.975, 
    5291.454,
  5427.981, 5423.041, 5417.741, 5411.942, 5406.055, 5398.043, 5397.687, 
    5376.663, 5377.098, 5363.735, 5347.475, 5333.115, 5315.482, 5296.023, 
    5271.762,
  5393.287, 5389.322, 5383.944, 5380.018, 5375.552, 5370.381, 5361.571, 
    5364.594, 5348.244, 5337.09, 5326.803, 5310.854, 5295.526, 5274.919, 
    5252.673,
  5358.154, 5355.711, 5350.534, 5349.464, 5344.899, 5342.616, 5338.054, 
    5328.216, 5324.474, 5317.309, 5303.496, 5290.498, 5275.187, 5255.448, 
    5232.088,
  5323.497, 5323.06, 5319.668, 5318.929, 5316.608, 5314.169, 5310.254, 
    5308.905, 5300.608, 5290.718, 5281.871, 5268.704, 5252.843, 5233.222, 
    5210.179,
  5293.46, 5292.925, 5290.154, 5291.16, 5289.049, 5288.721, 5284.669, 
    5278.965, 5274.074, 5268.748, 5258.109, 5245.323, 5230.585, 5211.39, 
    5188.33,
  5265.366, 5265.181, 5263.412, 5262.471, 5260.606, 5259.009, 5255.963, 
    5253.802, 5248.316, 5240.645, 5232.544, 5221.369, 5206.294, 5187.736, 
    5165.579,
  5237.98, 5235.561, 5233.453, 5233.529, 5232.262, 5229.929, 5226.298, 
    5221.001, 5217.037, 5212.893, 5205.708, 5195.29, 5181.966, 5164.838, 
    5143.142,
  5408.126, 5408.875, 5410.273, 5408.608, 5406.838, 5400.918, 5392.885, 
    5386.962, 5374.955, 5356.693, 5340.987, 5324.803, 5306.666, 5288.769, 
    5273.188,
  5370.484, 5372.963, 5375.022, 5372.682, 5367.946, 5363.025, 5361.42, 
    5344.729, 5332.937, 5326.778, 5309.178, 5294.542, 5277.442, 5263.974, 
    5247.425,
  5330.997, 5333.812, 5335.135, 5333.648, 5328.909, 5326.226, 5311, 5323.906, 
    5296.122, 5286.759, 5275.225, 5264.283, 5248.763, 5236.066, 5224.129,
  5282.564, 5286.091, 5287.609, 5286.187, 5282.765, 5276.971, 5281.146, 
    5259.137, 5266.034, 5253.287, 5241.798, 5232.979, 5223.521, 5212.758, 
    5202.156,
  5236.986, 5238.161, 5238.276, 5239.025, 5239.3, 5237.31, 5230.081, 
    5238.702, 5222.747, 5219.332, 5214.219, 5205.715, 5199.586, 5189.664, 
    5182.522,
  5192.671, 5193.929, 5193.497, 5196.416, 5196.08, 5197.837, 5196.736, 
    5188.783, 5191.24, 5191.689, 5184.019, 5181.464, 5176.301, 5170.18, 
    5163.747,
  5152.96, 5154.154, 5153.398, 5155.458, 5157.707, 5159.175, 5160.202, 
    5165.233, 5162.378, 5159.566, 5160.612, 5158.53, 5154.268, 5150.296, 
    5145.138,
  5113.528, 5113.463, 5112.968, 5117.572, 5120.297, 5125.844, 5128.629, 
    5129.738, 5133.095, 5137.643, 5137.176, 5136.542, 5135.463, 5132.673, 
    5128.39,
  5075.795, 5075.178, 5075.048, 5078.628, 5083.506, 5090.59, 5097.45, 
    5105.767, 5109.574, 5111.565, 5114.872, 5117.034, 5116.038, 5114.486, 
    5110.648,
  5044.486, 5039.186, 5036.812, 5040.14, 5045.235, 5053.418, 5062.209, 
    5070.539, 5079.453, 5088.085, 5093.308, 5096.604, 5097.422, 5096.285, 
    5091.741,
  5224.399, 5238.136, 5251.224, 5261.798, 5272.659, 5281.124, 5291.166, 
    5304.122, 5311.897, 5315.335, 5319.88, 5321.423, 5317.078, 5309.807, 
    5299.475,
  5195.491, 5209.279, 5224.256, 5236.329, 5245.211, 5256.112, 5267.915, 
    5273.175, 5280.495, 5291.19, 5290.184, 5290.27, 5285.165, 5279.554, 
    5265.775,
  5165.917, 5179.578, 5193.711, 5205.36, 5215.849, 5228.144, 5229.991, 
    5253.185, 5248.242, 5253.254, 5256.479, 5256.322, 5250.775, 5243.199, 
    5233.243,
  5133.329, 5144.476, 5157.349, 5167.43, 5179.565, 5183.91, 5206.138, 
    5197.581, 5219.556, 5220.914, 5218.33, 5217.166, 5215.977, 5208.027, 
    5197.831,
  5100.796, 5106.548, 5115.079, 5126.008, 5137.381, 5149.094, 5151.604, 
    5174.444, 5169.658, 5176.833, 5179.561, 5177.804, 5178.826, 5170.477, 
    5165.485,
  5074.271, 5075.224, 5078.057, 5083.935, 5089.462, 5097.659, 5107.61, 
    5108.199, 5126.564, 5135.164, 5133.407, 5138.501, 5138.689, 5135.513, 
    5131.774,
  5046.169, 5041.042, 5039.358, 5042.039, 5048.772, 5055.349, 5063.235, 
    5077.637, 5084.048, 5088.05, 5096.759, 5100.545, 5101.893, 5102.42, 
    5100.969,
  5030.703, 5017.257, 5007.18, 5003.684, 5002.348, 5008.357, 5015.567, 
    5022.493, 5035.208, 5049.216, 5056.217, 5062.895, 5068.624, 5071.272, 
    5071.726,
  5029.379, 5010.183, 4993.032, 4981.579, 4975.263, 4973.563, 4976.848, 
    4987.562, 4997.231, 5006.659, 5018.511, 5029.355, 5036.333, 5041.784, 
    5045.333,
  5043.798, 5018.139, 4996.816, 4980.689, 4966.506, 4960.277, 4959.285, 
    4962.875, 4973.139, 4986.667, 4997.746, 5006.9, 5014.442, 5020.351, 
    5023.787,
  5119.12, 5126.327, 5134.681, 5143.821, 5153.664, 5161.391, 5169.375, 
    5178.623, 5185.541, 5191.001, 5198.596, 5206.385, 5211.924, 5217.967, 
    5223.692,
  5098.463, 5103.446, 5109.565, 5117.56, 5124.863, 5134.707, 5144.686, 
    5149.104, 5156.092, 5166.463, 5170, 5177.023, 5181.898, 5189.018, 5191.477,
  5076.995, 5079.866, 5083.424, 5091.358, 5096.728, 5110.297, 5110.951, 
    5128.878, 5128.404, 5135.929, 5142.054, 5149.215, 5153.757, 5159.022, 
    5165.183,
  5061.95, 5059.639, 5060.785, 5063.229, 5070.327, 5072.378, 5090.42, 
    5085.813, 5103.171, 5108.155, 5113.741, 5119.12, 5125.925, 5131.089, 
    5135.903,
  5055.49, 5047.494, 5043.609, 5042.66, 5045.342, 5051.238, 5051.301, 
    5067.65, 5068.474, 5073.754, 5084.831, 5088.563, 5097.112, 5101.213, 
    5109.058,
  5059.386, 5045.682, 5035.269, 5030.439, 5026.743, 5026.868, 5032.051, 
    5029.033, 5037.91, 5044.683, 5046.934, 5053.568, 5059.604, 5064.936, 
    5071.678,
  5069.571, 5052.456, 5037.264, 5025.959, 5019.002, 5013.855, 5010.863, 
    5012.998, 5011.502, 5009.609, 5014.739, 5017.525, 5020.837, 5025.533, 
    5030.926,
  5084.678, 5065.847, 5047.205, 5032.25, 5017.768, 5008.112, 4999.755, 
    4991.602, 4987.38, 4985.345, 4981.489, 4979.731, 4980.571, 4982.047, 
    4985.548,
  5096.709, 5078.778, 5059.582, 5042.191, 5026.225, 5011.544, 4998.356, 
    4988.594, 4977.62, 4967.314, 4960.647, 4954.088, 4948.486, 4945.655, 
    4945.131,
  5108.284, 5088.592, 5068.551, 5050.395, 5030.653, 5013.758, 4997.893, 
    4982.684, 4971.068, 4960.952, 4951.256, 4942.322, 4935.669, 4930.895, 
    4927.916,
  5065.998, 5066.786, 5068.811, 5073.296, 5078.947, 5086.042, 5095.158, 
    5106.7, 5117.778, 5129.006, 5142.254, 5156.019, 5166.945, 5178.183, 
    5188.891,
  5061.762, 5058.326, 5056.12, 5056.619, 5057.647, 5062.751, 5069.673, 
    5075.002, 5084.533, 5097.09, 5105.771, 5118.095, 5128.285, 5141.72, 
    5149.204,
  5060.593, 5052.851, 5046.859, 5044.335, 5041.678, 5046.714, 5044.34, 
    5056.254, 5056.164, 5064.667, 5073.358, 5084.283, 5093.251, 5102.459, 
    5113.931,
  5059.878, 5049.403, 5041.178, 5033.486, 5029.562, 5024.063, 5031.119, 
    5025.041, 5035.443, 5039.096, 5044.823, 5052.24, 5061.401, 5070.213, 
    5077.91,
  5055.407, 5043.559, 5034.201, 5025.438, 5019.504, 5014.031, 5007.596, 
    5011.331, 5006.51, 5009.33, 5016.982, 5020.568, 5029.544, 5035.004, 
    5045.235,
  5047.962, 5033.875, 5022.502, 5013.96, 5005.423, 4999.714, 4996.212, 
    4989.081, 4989.437, 4989.292, 4987.806, 4991.069, 4996.771, 5002.384, 
    5010.31,
  5040.831, 5024.857, 5010.37, 4998.977, 4990.438, 4983.068, 4977.43, 
    4975.716, 4971.414, 4968.249, 4969.976, 4970.454, 4971.639, 4974.563, 
    4979.825,
  5037.598, 5017.046, 4998.132, 4984.273, 4971.016, 4962.545, 4955.604, 
    4950.363, 4948.333, 4949.086, 4948.359, 4950.041, 4952.81, 4955.621, 
    4958.796,
  5038.517, 5015.174, 4991.908, 4972.841, 4957.182, 4944.716, 4934.341, 
    4928.611, 4923.218, 4921.199, 4923.516, 4927.194, 4931.24, 4935.966, 
    4940.206,
  5044.979, 5015.372, 4988.504, 4966.032, 4944.923, 4929.413, 4917.037, 
    4906.894, 4901.08, 4898.219, 4897.354, 4899.66, 4905.066, 4912.647, 
    4919.666,
  5024.129, 5016.272, 5010.939, 5009.276, 5010.748, 5016.003, 5028.472, 
    5046.977, 5066.55, 5087.953, 5108.851, 5130.638, 5150.609, 5169.159, 
    5186.035,
  5018.775, 5010.791, 5004.744, 5001.459, 4999.067, 5002.021, 5007.302, 
    5015.518, 5031.119, 5052.199, 5069.813, 5090.177, 5106.735, 5127.98, 
    5140.41,
  5012.231, 5003.189, 4996.797, 4993.518, 4991.31, 4994.037, 4991.654, 
    5002.131, 5005.003, 5016.827, 5032.25, 5049.732, 5066.16, 5081.085, 
    5097.489,
  5004.913, 4993.789, 4986.847, 4981.917, 4980.738, 4977.927, 4986.418, 
    4979.167, 4990.802, 4996.235, 5005.651, 5016.962, 5031.301, 5045.975, 
    5058.376,
  4998.011, 4984.703, 4974.602, 4967.743, 4963.674, 4964.564, 4961.488, 
    4972.743, 4971.445, 4975.778, 4984.65, 4991.71, 5003.117, 5012.131, 
    5025.964,
  4994.341, 4978.031, 4964.154, 4953.603, 4945.077, 4940.485, 4942.009, 
    4938.984, 4947.835, 4958.073, 4962.931, 4972.479, 4981.31, 4989.879, 
    4999.971,
  4990.78, 4973.829, 4956.684, 4941.937, 4929.519, 4919.906, 4914.003, 
    4916.267, 4918.684, 4923.97, 4935.617, 4947.292, 4956.772, 4967.188, 
    4977.11,
  4987.298, 4969.198, 4948.807, 4931.083, 4913.069, 4899.688, 4890.208, 
    4884.482, 4885.561, 4894.296, 4904.436, 4916.087, 4928.951, 4941.362, 
    4953.759,
  4982.15, 4964.264, 4941.351, 4920.687, 4899.715, 4882.027, 4869.143, 
    4864.008, 4862.064, 4864.732, 4873.34, 4885.603, 4898.408, 4912.062, 
    4926.512,
  4977.893, 4957.876, 4932.165, 4909.862, 4886.161, 4866.236, 4851.729, 
    4842.457, 4841.646, 4846.226, 4853.199, 4861.521, 4871.943, 4884.434, 
    4899.026,
  4980.397, 4982.752, 4983.446, 4982.842, 4982.374, 4980.878, 4979.621, 
    4980.392, 4982.1, 4988.305, 5002.136, 5021.707, 5045.371, 5072.52, 
    5103.509,
  4966.796, 4969.836, 4970.506, 4969.137, 4966.979, 4966.118, 4966.107, 
    4962.639, 4963.207, 4969.713, 4977.696, 4994.643, 5013.891, 5042.021, 
    5068.792,
  4954.397, 4958.774, 4958.869, 4956.835, 4952.777, 4952.643, 4947.471, 
    4953.216, 4948.928, 4950.909, 4956.926, 4969.734, 4986.723, 5007.343, 
    5035.388,
  4946.007, 4948.678, 4946.421, 4941.619, 4937.186, 4931.836, 4936.101, 
    4928.362, 4936.05, 4937.264, 4941.418, 4948.803, 4963.186, 4983.049, 
    5006.151,
  4941.487, 4939.589, 4933.488, 4924.706, 4917.607, 4913.716, 4909.561, 
    4917.449, 4915.641, 4919.769, 4926.883, 4931.694, 4943.365, 4956.87, 
    4980.917,
  4941.238, 4932.983, 4923.359, 4909.889, 4898.526, 4892.338, 4890.718, 
    4887.748, 4894.195, 4902.922, 4908.404, 4916.671, 4926.021, 4938.312, 
    4956.897,
  4932.187, 4925.015, 4912.72, 4896.705, 4883.283, 4873.201, 4868.553, 
    4870.063, 4871.361, 4875.867, 4887.915, 4899.54, 4909.662, 4920.714, 
    4935.954,
  4930.773, 4917.581, 4901.332, 4883.653, 4865.196, 4853.559, 4844.992, 
    4841.11, 4844.03, 4852.917, 4863.785, 4878.634, 4893.975, 4907.396, 
    4920.868,
  4921.962, 4910.083, 4890.765, 4868.91, 4850.68, 4836.531, 4826.635, 
    4822.043, 4820.888, 4826.156, 4838.263, 4855.859, 4875.101, 4892.618, 
    4907.306,
  4911.017, 4896.647, 4874.71, 4854.864, 4834.837, 4818.61, 4806.333, 
    4799.104, 4799.588, 4806.217, 4817.456, 4833.976, 4856.431, 4878.381, 
    4896.333,
  4904.511, 4910.949, 4921.29, 4932.018, 4943.628, 4954.419, 4967.398, 
    4981.441, 4994.711, 5006.061, 5020.342, 5036.419, 5052.448, 5068.809, 
    5087.949,
  4883.843, 4892.065, 4903.016, 4915.092, 4926.615, 4939.526, 4953.254, 
    4964.682, 4977.867, 4993.109, 5004.854, 5019.066, 5032.609, 5050.233, 
    5064.156,
  4867.868, 4878.125, 4890.363, 4902.887, 4914.215, 4929.449, 4937.627, 
    4955.53, 4964.419, 4975.845, 4988.524, 5002.033, 5014.706, 5026.988, 
    5041.448,
  4863.202, 4874.433, 4887.021, 4898.099, 4910.616, 4916.373, 4933.011, 
    4933.328, 4949.613, 4959.87, 4971.336, 4982.407, 4995.694, 5008.487, 
    5020.583,
  4866.657, 4877.997, 4890.284, 4900.081, 4906.194, 4913.063, 4913.136, 
    4925.587, 4930.434, 4937.159, 4951.951, 4961.518, 4975.651, 4985.353, 
    4998.816,
  4880.504, 4892.444, 4900.126, 4905.713, 4904.756, 4901.388, 4902.225, 
    4898.824, 4905.143, 4916.284, 4924.382, 4937.066, 4950.653, 4963.241, 
    4976.166,
  4896.979, 4905.703, 4907.025, 4905.42, 4900.314, 4892.071, 4884.698, 
    4885.458, 4886.412, 4888.28, 4898.052, 4908.915, 4921.612, 4935.622, 
    4948.899,
  4906.92, 4906.905, 4900.812, 4894.42, 4882.476, 4870.154, 4861.287, 
    4856.424, 4857.297, 4865.143, 4871.135, 4879.997, 4892.807, 4907.222, 
    4922.131,
  4904.735, 4903.367, 4892.259, 4878.948, 4858.62, 4841.563, 4831.452, 
    4833.079, 4835.054, 4839.013, 4844.973, 4853.96, 4864.293, 4878.481, 
    4893.956,
  4897.462, 4888.017, 4873.159, 4853.865, 4832.206, 4817.455, 4808.111, 
    4805.358, 4808.203, 4815.508, 4821.676, 4829.702, 4840.31, 4854.694, 
    4870.648,
  4874.289, 4895.923, 4919.682, 4942.997, 4966.357, 4984.958, 5000.778, 
    5014.079, 5024.401, 5030.637, 5036.781, 5043.54, 5048.107, 5051.335, 
    5054.664,
  4854.52, 4873.731, 4895.395, 4918.846, 4940.454, 4961.029, 4979.506, 
    4990.689, 5001.056, 5013.269, 5020.009, 5028.953, 5034.799, 5041.618, 
    5044.562,
  4850.296, 4865.073, 4881.107, 4901.511, 4920.109, 4943.065, 4951.989, 
    4974.158, 4982.195, 4993.115, 5002.888, 5013.009, 5021.517, 5028.922, 
    5035.483,
  4863.864, 4870.108, 4879.534, 4890.971, 4906.029, 4917.292, 4939.862, 
    4942.469, 4961.719, 4974.253, 4986.419, 4996.063, 5007.404, 5017.034, 
    5026.382,
  4884.568, 4884.091, 4886.003, 4890.783, 4897.331, 4909.863, 4915.548, 
    4935.052, 4943.892, 4953.042, 4968.639, 4978.449, 4991.764, 5002.202, 
    5015.64,
  4900.384, 4898.246, 4895.984, 4896.741, 4896.868, 4900.273, 4909.668, 
    4913.578, 4924.917, 4940.98, 4950.319, 4963.908, 4976.3, 4989.571, 5003.83,
  4909.497, 4905.47, 4901.655, 4898.531, 4897.511, 4897.169, 4898.292, 
    4906.393, 4914.71, 4922.193, 4935.302, 4948.701, 4961.625, 4976.407, 
    4991.751,
  4897.491, 4891.467, 4886.399, 4883.066, 4878.514, 4877.608, 4879.754, 
    4883.574, 4892.352, 4907.406, 4920.812, 4934.213, 4948.952, 4964.435, 
    4980.241,
  4883.344, 4877.138, 4868.092, 4859.899, 4852.488, 4848.592, 4848.771, 
    4856.902, 4869.05, 4883.791, 4901.189, 4919.21, 4935.341, 4951.846, 
    4968.281,
  4871.889, 4862.064, 4851.967, 4842.752, 4833.058, 4826.252, 4823.57, 
    4825.134, 4835.813, 4856.416, 4880.12, 4901.978, 4921.417, 4938.983, 
    4955.301,
  4880.137, 4885.191, 4898.547, 4921.685, 4953.523, 4986.65, 5019.658, 
    5053.098, 5082.953, 5107.693, 5131.026, 5153.288, 5170.657, 5185.031, 
    5194.908,
  4883.574, 4882.078, 4887.257, 4903.662, 4927.61, 4960.776, 4996.169, 
    5026.35, 5056.328, 5088.221, 5112.25, 5134.625, 5152.387, 5168.627, 
    5176.943,
  4892.368, 4887.552, 4886.56, 4894.633, 4909.615, 4941.823, 4967.749, 
    5009.217, 5036.984, 5064.447, 5090.99, 5114.375, 5133.569, 5148.226, 
    5160.836,
  4899.952, 4891.761, 4890.89, 4891.681, 4902, 4913.858, 4953.004, 4971.647, 
    5011.617, 5043.073, 5071.425, 5093.773, 5115.377, 5131.291, 5143.072,
  4899.112, 4892.182, 4889.05, 4889.468, 4896.011, 4910.839, 4923.072, 
    4962.575, 4992.295, 5018.073, 5050.646, 5073.208, 5096.421, 5111.479, 
    5126.14,
  4887.312, 4880.222, 4880.715, 4885.966, 4890.812, 4899.589, 4918.224, 
    4932.436, 4964.6, 5001.922, 5027.973, 5055.077, 5076.821, 5094.774, 
    5108.142,
  4877.951, 4866.574, 4866.845, 4873.35, 4884.117, 4893.714, 4905.279, 
    4926.98, 4952.974, 4976.383, 5008.312, 5035.493, 5057.204, 5076.228, 
    5089.989,
  4874.233, 4860.826, 4854.77, 4860.145, 4870.652, 4884.194, 4896.738, 
    4908.69, 4929.109, 4960.745, 4990.332, 5016.363, 5040.136, 5059.252, 
    5073.834,
  4877.256, 4862.632, 4853.063, 4850.198, 4856.123, 4869.731, 4883.986, 
    4903.531, 4923.606, 4944.937, 4971.929, 4999.774, 5023.369, 5042.887, 
    5058.696,
  4880.977, 4862.992, 4850.587, 4845.422, 4843.975, 4852.795, 4866.663, 
    4883.549, 4903.554, 4929.959, 4957.912, 4985.126, 5009.313, 5029.626, 
    5046.263,
  4888.061, 4883.078, 4894.118, 4906.678, 4920.168, 4932.75, 4945.669, 
    4963.853, 4987.19, 5014.395, 5046.465, 5082.549, 5118.226, 5154.585, 
    5188.473,
  4895.812, 4890.301, 4894.559, 4908.191, 4921.203, 4935.53, 4952.296, 
    4968.957, 4991.32, 5022.529, 5054.27, 5089.408, 5123.854, 5160.155, 
    5191.614,
  4902.174, 4896.803, 4897.08, 4908.808, 4922.18, 4941.375, 4955.072, 
    4979.015, 5003.82, 5029.614, 5061.327, 5094.018, 5129.738, 5161.868, 
    5194.208,
  4903.588, 4901.442, 4900.761, 4907.694, 4923.731, 4936.335, 4963.188, 
    4977.158, 5004.275, 5033.672, 5065.771, 5097.665, 5132.235, 5165.823, 
    5195.653,
  4898.86, 4894.347, 4901.297, 4907.437, 4920.832, 4940.719, 4957.083, 
    4984.937, 5012.656, 5035.758, 5067.879, 5099.696, 5134.504, 5163.98, 
    5193.603,
  4896.977, 4886.451, 4892.247, 4903.918, 4917.963, 4934.862, 4959.326, 
    4979.585, 5003.497, 5038.17, 5066.817, 5101.13, 5133.978, 5166.257, 
    5192.564,
  4892.847, 4883.62, 4883.253, 4896.375, 4913.643, 4932.913, 4951.918, 
    4979.825, 5009.144, 5034.97, 5066.692, 5099.876, 5131.887, 5162.681, 
    5189.142,
  4893.554, 4880.292, 4877.584, 4888.564, 4905.356, 4925.575, 4947.867, 
    4967.951, 4994.353, 5028.856, 5062.365, 5095.341, 5128.723, 5159.399, 
    5185.863,
  4894.21, 4881.104, 4875.655, 4881.432, 4897.839, 4918.652, 4940.369, 
    4964.613, 4992.306, 5020.834, 5053.933, 5088.957, 5122.211, 5152.859, 
    5179.49,
  4901.508, 4884.496, 4875.251, 4877.931, 4890.705, 4910.428, 4933.655, 
    4953.537, 4977.442, 5009.034, 5044.677, 5081.063, 5115.163, 5146.729, 
    5173.714,
  4923.603, 4917.463, 4909.653, 4900.937, 4891.984, 4883.74, 4877.111, 
    4877.938, 4886.26, 4895.984, 4910.355, 4931.065, 4956.036, 4983.99, 
    5015.356,
  4926.397, 4921.628, 4912.511, 4901.866, 4890.254, 4879.087, 4872.461, 
    4872.333, 4879.182, 4896.875, 4916.635, 4941.479, 4968.61, 5000.859, 
    5032.114,
  4931.536, 4926.45, 4919.622, 4908.82, 4895.249, 4886.729, 4875.382, 
    4880.913, 4894.558, 4909.787, 4931.727, 4958.528, 4988.353, 5018.542, 
    5052.77,
  4935.269, 4933.688, 4929.85, 4918.799, 4911.735, 4896.303, 4899.244, 
    4896.443, 4908.633, 4929.314, 4955.541, 4981.945, 5013.558, 5046.23, 
    5080.625,
  4940.602, 4940.935, 4941.438, 4936.84, 4932.092, 4927.589, 4924.259, 
    4927.884, 4949.074, 4959.658, 4986.876, 5012.226, 5045.185, 5073.641, 
    5107.488,
  4946.198, 4950.02, 4952.884, 4953.641, 4953.253, 4952.36, 4958.327, 
    4964.252, 4972.95, 4997.552, 5020.057, 5047.166, 5075.833, 5106.02, 
    5133.055,
  4954.391, 4958.776, 4965.305, 4970.986, 4975.466, 4982.122, 4986.444, 
    4999.195, 5016.796, 5032.622, 5053.079, 5078.597, 5104.341, 5131.433, 
    5155.499,
  4962.824, 4968.481, 4976.162, 4985.431, 4991.83, 5001.691, 5013.608, 
    5025.247, 5037.891, 5059.003, 5080.898, 5104.687, 5129.906, 5154.062, 
    5175.239,
  4973.542, 4978.132, 4987.302, 4998.35, 5008.415, 5019.708, 5031.202, 
    5048.232, 5066.117, 5084.084, 5103.614, 5127.526, 5150.458, 5172.064, 
    5190.21,
  4985.647, 4987.097, 4994.513, 5007.088, 5017.94, 5032.385, 5046.864, 
    5062.182, 5078.84, 5099.912, 5122.4, 5145.658, 5167.72, 5188.297, 5204.586,
  4922.211, 4903.181, 4884.238, 4871.526, 4867.901, 4874.566, 4885.814, 
    4894.698, 4905.692, 4919.621, 4938.085, 4958.261, 4977.532, 4996.636, 
    5014.867,
  4919.37, 4893.636, 4868.749, 4851.191, 4846.628, 4856.365, 4876.026, 
    4888.543, 4899.998, 4918.277, 4937.095, 4955.53, 4972.152, 4989.997, 
    5005.716,
  4924.99, 4894.036, 4866.147, 4845.595, 4839.003, 4852.26, 4868.346, 
    4886.546, 4904.933, 4920.767, 4938.826, 4954.487, 4970.228, 4983.835, 
    5000.255,
  4939.134, 4907.154, 4878.93, 4855.833, 4850.451, 4852.279, 4874.414, 
    4887.219, 4905.036, 4923.884, 4942.634, 4956.073, 4970.576, 4984.233, 
    5001.086,
  4961.394, 4930.369, 4902.317, 4882.191, 4869.844, 4876.483, 4880.581, 
    4898.626, 4919.968, 4932.221, 4949.437, 4960.73, 4975.421, 4989.023, 
    5009.42,
  4991.92, 4962.422, 4934.49, 4914.834, 4901.94, 4897.902, 4909.338, 
    4917.669, 4927.542, 4946.273, 4959.549, 4974.277, 4990.276, 5008.591, 
    5026.711,
  5025.896, 5002.097, 4976.816, 4956.301, 4943.251, 4938.085, 4935.7, 
    4947.056, 4961.383, 4972.865, 4987.055, 5002.747, 5018.301, 5034.319, 
    5051.33,
  5058.432, 5042.542, 5023.613, 5008.024, 4993.87, 4988.596, 4989.495, 
    4992.181, 4998.746, 5012.639, 5025.01, 5037.973, 5051.1, 5064.731, 
    5077.508,
  5085.945, 5075.192, 5061.739, 5050.477, 5041.354, 5036.15, 5034.132, 
    5039.186, 5045.65, 5052.387, 5060.545, 5070.484, 5079.543, 5088.312, 
    5096.844,
  5109.011, 5101.945, 5094.163, 5086.016, 5078.923, 5075.566, 5074.421, 
    5074.515, 5077.127, 5083.124, 5088.965, 5094.573, 5099.691, 5104.584, 
    5108.665,
  4896.062, 4888.802, 4898.074, 4913.99, 4930.31, 4942.751, 4951.557, 
    4957.786, 4963.261, 4968.803, 4978.539, 4994.399, 5023.328, 5063.2, 
    5103.405,
  4916.868, 4903.36, 4903.459, 4914.43, 4929.399, 4941.377, 4950.833, 
    4955.738, 4957.034, 4962.104, 4970.137, 4982.615, 5006.031, 5046.769, 
    5086.364,
  4946.878, 4930.339, 4924.928, 4929.59, 4937.478, 4948.49, 4950.48, 
    4951.955, 4954.632, 4959.063, 4966.081, 4974.953, 4994.309, 5027.802, 
    5070.559,
  4978.835, 4960.106, 4950.799, 4946.607, 4950.53, 4947.674, 4951.29, 
    4950.42, 4954.051, 4960.319, 4967.106, 4972.402, 4987.723, 5018.53, 
    5058.889,
  5013.327, 4992, 4976.547, 4967.175, 4960.404, 4960.434, 4957.063, 4956.97, 
    4963.971, 4966.339, 4972.01, 4974.591, 4987.354, 5009.381, 5048.003,
  5050.185, 5027.917, 5007.641, 4994.547, 4982.295, 4972.914, 4971.021, 
    4971.179, 4971.211, 4976.318, 4979.276, 4982.087, 4991.928, 5011.813, 
    5042.125,
  5085.873, 5064.467, 5043.324, 5026.092, 5011.532, 5000.508, 4987.706, 
    4982.892, 4984.088, 4986.739, 4989.232, 4993.689, 5001.036, 5016.633, 
    5041.104,
  5117.467, 5098.617, 5078.031, 5061.883, 5045.684, 5032.285, 5020.166, 
    5009.901, 5001.616, 5000.73, 5002.918, 5007.671, 5015.501, 5028.472, 
    5047.365,
  5144.005, 5127.118, 5108.753, 5091.266, 5075.73, 5062.292, 5050.188, 
    5041.178, 5033.099, 5027.664, 5025.403, 5028.361, 5034.111, 5044.014, 
    5057.677,
  5166.811, 5150.376, 5135.017, 5119.276, 5102.335, 5088.536, 5076.758, 
    5067.367, 5059.401, 5054.358, 5051.221, 5051.508, 5054.887, 5062.078, 
    5071.973,
  4999.549, 4996.577, 4995.256, 4994.186, 4996.722, 5002.297, 5011.153, 
    5021.668, 5032.737, 5041.798, 5052.2, 5063.813, 5077.564, 5095.591, 
    5122.378,
  5014.455, 5007.77, 5006.241, 5004.413, 5006.122, 5009.509, 5018.381, 
    5027.069, 5036.678, 5048.784, 5060.535, 5074.784, 5089.984, 5112.499, 
    5139.061,
  5030.347, 5020.396, 5015.834, 5014.484, 5014.44, 5019.034, 5022.677, 
    5032.213, 5042.178, 5052.906, 5066.414, 5082.626, 5101.387, 5123.594, 
    5151.397,
  5055.673, 5038.375, 5026.24, 5020.188, 5019.267, 5019.403, 5026.509, 
    5031.034, 5040.028, 5052.881, 5067.287, 5084.926, 5106.702, 5132.218, 
    5160.714,
  5086.513, 5066.958, 5048.549, 5036.64, 5029.002, 5028.15, 5028.413, 
    5034.593, 5043.936, 5050.653, 5064.497, 5080.902, 5104.021, 5129.762, 
    5159.209,
  5115.772, 5095.848, 5074.79, 5059.426, 5046.39, 5040.304, 5038.536, 
    5039.913, 5041.416, 5051.274, 5058.158, 5072.192, 5093.819, 5123.356, 
    5154.12,
  5146.051, 5127.345, 5106.029, 5087.873, 5070.465, 5059.078, 5050.847, 
    5050.089, 5050.771, 5051.28, 5052.708, 5060.855, 5079.171, 5108.307, 
    5141.514,
  5172.796, 5154.453, 5134.199, 5116.771, 5097.424, 5080.835, 5067.167, 
    5057.943, 5052.643, 5051.787, 5050.008, 5051.458, 5066.152, 5093.69, 
    5128.191,
  5199.969, 5182.115, 5162.065, 5143.817, 5126.065, 5109.069, 5090.334, 
    5076.315, 5064.768, 5056.726, 5051.403, 5048.979, 5057.305, 5081.045, 
    5114.379,
  5225.374, 5204.339, 5183.971, 5165.216, 5145.801, 5129.869, 5113.841, 
    5096.729, 5080.194, 5067.453, 5057.742, 5052.896, 5056.222, 5074.798, 
    5105.613,
  5056.982, 5054.894, 5054.738, 5053.935, 5053.139, 5047.966, 5038.137, 
    5028.377, 5015.195, 4997.222, 4989.709, 4995.328, 5009.975, 5033.348, 
    5063.376,
  5069.632, 5064.238, 5063.719, 5061.454, 5061.051, 5053.077, 5048.083, 
    5028.768, 5009.311, 4992.959, 4982.855, 4988.734, 5005.139, 5031.507, 
    5062.513,
  5085.488, 5074.236, 5069.856, 5069.119, 5064.972, 5064.384, 5049.626, 
    5039.582, 5021.252, 4998.954, 4987.55, 4992.747, 5010.581, 5034.699, 
    5068.992,
  5109.509, 5091.43, 5079.542, 5072.045, 5071.888, 5063.823, 5062.079, 
    5044.386, 5025.04, 5012.361, 5003.882, 5009.152, 5026.232, 5052.677, 
    5087.774,
  5138.555, 5116.604, 5098.462, 5084.473, 5076.631, 5073.976, 5066.323, 
    5056.009, 5048.864, 5031.942, 5028.33, 5032.595, 5051.419, 5074.394, 
    5111.339,
  5164.241, 5142.763, 5121.489, 5103.804, 5089.351, 5078.965, 5076.666, 
    5068.227, 5057.356, 5053.982, 5053.095, 5060.326, 5078.71, 5106.538, 
    5138.9,
  5190.129, 5167.786, 5145.876, 5127.129, 5109.993, 5096.143, 5085.349, 
    5082.421, 5080.05, 5076.149, 5078.158, 5088.928, 5107.48, 5135.112, 
    5166.003,
  5210.85, 5191.609, 5169.226, 5148.632, 5129.129, 5114.153, 5102.77, 
    5094.544, 5090.954, 5095.27, 5102.154, 5115.772, 5136.47, 5162.562, 
    5189.994,
  5226.874, 5211.314, 5191.691, 5170.945, 5151.071, 5134.299, 5120.981, 
    5113.619, 5110.18, 5112.528, 5121.33, 5137.482, 5157.328, 5181.408, 
    5206.136,
  5236.729, 5225.25, 5208.844, 5189.157, 5167.882, 5150.527, 5137.893, 
    5128.533, 5123.637, 5124.953, 5133.471, 5149.138, 5169.375, 5191.818, 
    5215.317,
  5049.583, 5039.839, 5031.986, 5022.063, 5012.87, 5001.711, 4989.397, 
    4982.276, 4978.281, 4977.634, 4984.078, 4997.27, 5017.593, 5043.602, 
    5072.545,
  5047.871, 5036.729, 5028.675, 5018.814, 5008.952, 4992.546, 4986.921, 
    4970.6, 4965.548, 4967.926, 4978.176, 4994.569, 5016.677, 5046.19, 5073.53,
  5052.403, 5039.022, 5028.971, 5018.396, 5004.974, 4994.888, 4973.514, 
    4966.948, 4956.718, 4960.493, 4972.35, 4993.073, 5017.994, 5046.125, 
    5075.662,
  5060.045, 5045.542, 5032.798, 5019.412, 5005.371, 4985.77, 4973.862, 
    4958.939, 4952.298, 4956.217, 4972.552, 4994.409, 5022.08, 5052.967, 
    5082.738,
  5069.351, 5052.86, 5039.042, 5022.374, 5005.281, 4986.983, 4970.269, 
    4959.191, 4957.106, 4960.51, 4978.334, 5001.178, 5030.418, 5059.53, 
    5091.383,
  5080.956, 5063.904, 5045.799, 5028.718, 5009.169, 4991.446, 4977.797, 
    4968.504, 4964.434, 4973.553, 4990.515, 5014.071, 5042.562, 5074.117, 
    5102.63,
  5094.984, 5076.951, 5058.147, 5040.366, 5021.496, 5004.906, 4990.1, 
    4982.624, 4983.93, 4992.344, 5008.856, 5032.091, 5059.583, 5089.299, 
    5116.567,
  5111.271, 5093.664, 5075.762, 5057.1, 5038.703, 5023.385, 5012.065, 
    5004.824, 5004.854, 5015.652, 5032.875, 5055.733, 5082.602, 5109.31, 
    5133.731,
  5128.816, 5113.67, 5096.942, 5079.885, 5064.813, 5051.222, 5040.053, 
    5035.751, 5038.474, 5047.436, 5062.784, 5083.988, 5107.602, 5131.027, 
    5153.792,
  5148.208, 5134.423, 5120.151, 5105.674, 5091.862, 5082.073, 5075.51, 
    5071.981, 5074.193, 5083.321, 5097.691, 5116.199, 5135.955, 5156.016, 
    5176.792,
  5020.44, 5015.797, 5015.517, 5017.051, 5019.692, 5021.459, 5022.641, 
    5023.945, 5025.403, 5024.188, 5021.329, 5016.608, 5010.672, 5006.822, 
    5009.406,
  4997.392, 4992.236, 4992.062, 4995.917, 5001.352, 5005.501, 5011.68, 
    5013.122, 5014.563, 5017.035, 5014.553, 5010.617, 5005.613, 5006.157, 
    5011.151,
  4985.415, 4978.076, 4977.548, 4980.299, 4987.033, 4995.845, 4997.48, 
    5007.337, 5009.279, 5011.212, 5009.305, 5007.684, 5008.042, 5011.724, 
    5019.909,
  4979.259, 4971.548, 4970.419, 4972.293, 4978.978, 4984.201, 4994.228, 
    4997.154, 5002.082, 5006.191, 5009.573, 5012.688, 5019.702, 5026.627, 
    5037.805,
  4980.991, 4972.349, 4968.576, 4970.889, 4974.596, 4982.323, 4987.371, 
    4996.283, 5005.483, 5008.851, 5018.459, 5025.697, 5036.171, 5043.459, 
    5056.104,
  4987.994, 4978.557, 4972.806, 4974.21, 4976.74, 4983.045, 4992.062, 
    5000.588, 5008.732, 5022.549, 5033.464, 5044.303, 5054.319, 5063.757, 
    5073.782,
  5002.58, 4993.044, 4986.218, 4985.825, 4988.941, 4995.646, 5002.356, 
    5015.511, 5029.879, 5042.286, 5054.12, 5065.031, 5074.132, 5082.714, 
    5090.935,
  5025.882, 5015.406, 5007.798, 5006.685, 5008.552, 5016.812, 5027.422, 
    5038.737, 5050.786, 5065.006, 5076.359, 5085.871, 5094.006, 5101.073, 
    5108.118,
  5060.846, 5050.641, 5043.028, 5040.97, 5043.286, 5049.212, 5057.141, 
    5069.512, 5080.93, 5090.634, 5099.243, 5107.663, 5114.375, 5120.875, 
    5127.24,
  5100.164, 5089.464, 5082.19, 5078.452, 5078.474, 5083.437, 5090.801, 
    5098.505, 5106.952, 5115.834, 5123.638, 5130.527, 5136.498, 5142.307, 
    5147.607,
  4992.59, 5005.084, 5021.617, 5039.306, 5057.44, 5071.424, 5080.973, 
    5087.993, 5090.59, 5087.291, 5081.114, 5073.832, 5067.278, 5063.187, 
    5060.302,
  4971.395, 4982.998, 5000.405, 5021.354, 5040.846, 5058.668, 5072.468, 
    5078.511, 5079.946, 5078.689, 5070.841, 5063.54, 5056.085, 5051.228, 
    5044.502,
  4957.079, 4964.841, 4982.079, 5003.872, 5027.108, 5049.549, 5058.519, 
    5070.789, 5071.403, 5069.079, 5062.194, 5054.784, 5048.551, 5042.291, 
    5035.647,
  4952.689, 4957.973, 4973.242, 4992.608, 5016.605, 5033.85, 5053.942, 
    5055.372, 5062.135, 5058.892, 5055.634, 5051.837, 5048.698, 5042.401, 
    5036.209,
  4959.579, 4962.642, 4974.169, 4992.443, 5011.607, 5032.964, 5042.414, 
    5053.21, 5055.366, 5056.659, 5059.439, 5057.338, 5055.424, 5050.76, 
    5048.54,
  4977.043, 4979.247, 4986.169, 5001.25, 5016.201, 5029.923, 5043.769, 
    5049.757, 5056.918, 5063.57, 5066.136, 5066.714, 5065.168, 5063.303, 
    5061.045,
  4999.885, 5001.519, 5005.66, 5016.437, 5029.587, 5042.758, 5051.262, 
    5062.685, 5070.281, 5074.8, 5077.024, 5077.411, 5076.048, 5074.972, 
    5073.867,
  5031.78, 5032.29, 5034.383, 5042.435, 5050.172, 5061.452, 5070.522, 
    5077.066, 5081.759, 5086.557, 5087.884, 5088.232, 5087.211, 5085.828, 
    5084.562,
  5066.081, 5066.104, 5066.655, 5071.204, 5077.023, 5083.737, 5088.996, 
    5095.894, 5100.077, 5102.501, 5103.105, 5102.513, 5100.605, 5098.748, 
    5096.932,
  5100.73, 5098.539, 5098.268, 5100.058, 5102.837, 5107.942, 5112.515, 
    5115.574, 5117.644, 5119.064, 5118.546, 5117.071, 5114.66, 5111.984, 
    5109.354,
  4955.167, 4960.253, 4970.896, 4985.971, 5006.194, 5027.478, 5046.991, 
    5062.315, 5074.889, 5080.797, 5080.739, 5071.562, 5057.969, 5042.428, 
    5029.245,
  4949.076, 4954.425, 4966.125, 4982.89, 5003.609, 5025.229, 5044.648, 
    5059.185, 5070, 5076.426, 5074.282, 5064.938, 5052.196, 5039.263, 5025.288,
  4951.061, 4957.166, 4969.797, 4987.246, 5008.59, 5032.089, 5045.663, 
    5059.809, 5069.414, 5072.494, 5068.968, 5060.326, 5051.239, 5037.967, 
    5025.028,
  4960.643, 4966.526, 4981.466, 4997.839, 5020.856, 5034.204, 5052.437, 
    5058.16, 5066.798, 5066.582, 5064.214, 5059.839, 5053.166, 5044.123, 
    5033.432,
  4975.797, 4983.541, 4996.782, 5013.986, 5029.206, 5046.538, 5052.015, 
    5060.631, 5062.362, 5064.21, 5063.875, 5061.873, 5059.29, 5053.038, 
    5047.327,
  4996.845, 5003.387, 5012.926, 5027.948, 5039.575, 5047.143, 5053.686, 
    5056.814, 5059.09, 5063.838, 5065.562, 5065.538, 5064.129, 5062.484, 
    5059.453,
  5019.069, 5023.997, 5030.144, 5038.908, 5047.089, 5053.361, 5054.943, 
    5060.305, 5064.562, 5068.579, 5069.304, 5070.301, 5070.022, 5070.351, 
    5069.633,
  5042.219, 5043.089, 5044.726, 5050.208, 5053.043, 5057.271, 5061.564, 
    5065.395, 5068.356, 5071.855, 5073.334, 5074.55, 5074.554, 5075.549, 
    5076.525,
  5068.275, 5066.297, 5064.722, 5064.767, 5066.296, 5068.531, 5070.25, 
    5074.356, 5077.508, 5079.734, 5080.58, 5080.979, 5081.183, 5081.599, 
    5082.424,
  5094.41, 5088.48, 5084.038, 5081.845, 5079.743, 5079.751, 5081.316, 
    5082.806, 5084.32, 5086.285, 5087.798, 5088.555, 5088.421, 5088.632, 
    5089.146,
  5002.965, 4990.354, 4981.157, 4976.066, 4975.069, 4979.156, 4987.27, 
    5001.142, 5012.854, 5022.452, 5032.27, 5043.293, 5050.738, 5055.113, 
    5053.924,
  5004.357, 4990.907, 4980.304, 4975.286, 4975.941, 4982.004, 4997.098, 
    5008.7, 5017.165, 5028.413, 5038.344, 5046.646, 5051.406, 5053.225, 
    5050.022,
  5013.713, 5000.393, 4989.577, 4985.5, 4986.517, 4998.474, 5005.331, 
    5017.565, 5028.58, 5037.639, 5045.337, 5051.44, 5055.849, 5056.296, 
    5053.549,
  5027.64, 5015.298, 5007.521, 5001.761, 5006.846, 5009.119, 5022.679, 
    5028.283, 5037.548, 5045.729, 5053.807, 5059.043, 5063.708, 5063.062, 
    5059.22,
  5041.913, 5032.334, 5026.688, 5022.693, 5022.708, 5029.638, 5033.29, 
    5040.948, 5051.675, 5055.454, 5063.349, 5067.875, 5071.978, 5070.103, 
    5066.448,
  5051.778, 5044.827, 5039.332, 5037.125, 5037.68, 5039.013, 5047.396, 
    5052.849, 5057.459, 5065.748, 5072.17, 5077.392, 5079.882, 5078.54, 
    5073.369,
  5057.691, 5054.066, 5050.526, 5048.137, 5048.938, 5052.887, 5055.133, 
    5061.844, 5069.32, 5075.788, 5081.046, 5085.765, 5087.192, 5085.603, 
    5081.122,
  5061.25, 5058.107, 5054.991, 5055.301, 5056.19, 5060.014, 5065.842, 
    5071.103, 5076.378, 5083.532, 5089.155, 5093.065, 5094.636, 5093.584, 
    5090.206,
  5063.923, 5062.46, 5061.795, 5062.396, 5064.911, 5068.932, 5073.31, 
    5080.07, 5087.046, 5092.298, 5096.539, 5099.961, 5101.469, 5101.347, 
    5099.653,
  5062.651, 5060.265, 5062.045, 5065.734, 5069.932, 5075.867, 5082.885, 
    5089.08, 5094.706, 5100.373, 5105.097, 5108.678, 5110.978, 5112.088, 
    5111.638,
  5121.573, 5106.523, 5091.364, 5078.039, 5067.324, 5054.617, 5039.704, 
    5028.876, 5020.189, 5016.082, 5019.673, 5025.721, 5029.735, 5031.958, 
    5032.376,
  5113.419, 5100.753, 5089.072, 5080.852, 5074.169, 5062.471, 5055.392, 
    5043.863, 5034.344, 5030.792, 5029.373, 5030.394, 5030.771, 5030.68, 
    5029.617,
  5109.947, 5100.905, 5092.987, 5089.05, 5081.521, 5078.802, 5066.119, 
    5061.013, 5054.458, 5048.739, 5044.586, 5042.404, 5038.404, 5033.948, 
    5028.428,
  5109.875, 5102.833, 5098.969, 5094.375, 5092.947, 5085.603, 5083.701, 
    5075.27, 5066.911, 5062.587, 5057.459, 5050.981, 5043.868, 5034.732, 
    5025.579,
  5111.338, 5106.348, 5105.467, 5103.394, 5101.975, 5099.069, 5095.086, 
    5087.583, 5086.749, 5075.947, 5071.403, 5061.223, 5052.34, 5038.464, 
    5026.312,
  5114.22, 5111.536, 5110.86, 5111.149, 5110.893, 5108.435, 5106.818, 
    5102.432, 5095.29, 5090.368, 5082.976, 5073.513, 5063.141, 5050.481, 
    5037.604,
  5117.345, 5117.938, 5118.43, 5119.498, 5120.286, 5120.704, 5117.347, 
    5114.407, 5111.488, 5105.239, 5097.515, 5089.257, 5079.275, 5068.895, 
    5057.909,
  5122.359, 5123.77, 5124.931, 5127.749, 5128.747, 5129.434, 5128.905, 
    5126.443, 5122.029, 5118.22, 5112.69, 5105.873, 5097.97, 5089.7, 5081.27,
  5127.206, 5130.159, 5133.395, 5136.181, 5138.759, 5140.188, 5139.308, 
    5138.829, 5137.633, 5134.302, 5129.774, 5125.069, 5119.227, 5112.84, 
    5106.245,
  5132.674, 5135.803, 5140.133, 5143.983, 5146.796, 5149.065, 5151.209, 
    5151.56, 5150.712, 5149.506, 5147.579, 5144.621, 5140.867, 5136.466, 
    5131.823,
  5161.758, 5163.032, 5164.397, 5163.073, 5160.948, 5156.094, 5149.22, 
    5140.353, 5129.874, 5115.979, 5102.975, 5090.866, 5080.844, 5074.526, 
    5073.911,
  5149.686, 5150.412, 5152.024, 5151.489, 5150.048, 5146.122, 5141.991, 
    5131.201, 5119.084, 5107.246, 5092.338, 5078.155, 5064.994, 5059.106, 
    5059.27,
  5143.765, 5145.071, 5146.583, 5147.826, 5146.667, 5145.51, 5134.158, 
    5128.459, 5115.449, 5100.483, 5083.322, 5066.008, 5050.002, 5043.834, 
    5049.582,
  5144.526, 5146.294, 5148.15, 5148.593, 5146.903, 5141.354, 5136.108, 
    5123.052, 5111.125, 5096.625, 5078.145, 5057.877, 5040.996, 5035.047, 
    5043.34,
  5148.939, 5150.591, 5152.502, 5152.096, 5149.585, 5143.343, 5135.172, 
    5126.712, 5115.344, 5096.865, 5080.278, 5059.43, 5044.95, 5039.012, 
    5048.126,
  5154.922, 5156.55, 5156.886, 5156.092, 5151.856, 5146.691, 5139.891, 
    5129.677, 5117.148, 5104.048, 5087.912, 5072.031, 5060.563, 5056.663, 
    5062.304,
  5161.205, 5163.154, 5162.514, 5161.605, 5158.434, 5153.74, 5146.205, 
    5138.888, 5128.549, 5115.836, 5102.484, 5090.795, 5082.592, 5080.29, 
    5084.475,
  5168.011, 5169.332, 5168.691, 5168.154, 5164.879, 5161.372, 5155.994, 
    5148.255, 5139.034, 5130.084, 5120.789, 5112.593, 5107.774, 5107.326, 
    5111.446,
  5175.058, 5177.076, 5177.38, 5176.724, 5175.034, 5172.001, 5166.749, 
    5161.614, 5155.088, 5147.837, 5140.939, 5135.734, 5132.981, 5133.604, 
    5137.472,
  5182.898, 5183.713, 5185.109, 5185.699, 5184.776, 5183.021, 5179.595, 
    5174.451, 5169.232, 5164.962, 5161.308, 5158.868, 5158.082, 5160.115, 
    5165.031,
  5121.28, 5128.687, 5140.771, 5153.421, 5166.603, 5176.375, 5182.747, 
    5187.881, 5189.047, 5185.931, 5180.553, 5173.698, 5164.929, 5155.878, 
    5148.325,
  5123.11, 5128.114, 5135.242, 5144.225, 5151.555, 5157.734, 5164.546, 
    5164.877, 5163.562, 5161.378, 5153.304, 5145.576, 5135.055, 5129.417, 
    5122.15,
  5123.935, 5127.161, 5131.559, 5138.073, 5141.392, 5149.051, 5143.336, 
    5150.032, 5142.759, 5137.941, 5129.195, 5120.562, 5110.496, 5103.292, 
    5102.471,
  5126.884, 5127.981, 5130.905, 5132.637, 5135.337, 5134.174, 5139.373, 
    5130.048, 5129.671, 5121.746, 5112.422, 5101.561, 5095.066, 5093.847, 
    5098.446,
  5134.163, 5132.836, 5133.662, 5133.561, 5133.749, 5133.06, 5128.196, 
    5128.283, 5119.255, 5109.287, 5103.18, 5096.521, 5097.525, 5099.64, 
    5105.548,
  5140.957, 5138.716, 5137.017, 5136.101, 5133.794, 5131.906, 5128.563, 
    5120.873, 5115.457, 5111.313, 5107.677, 5107, 5109.042, 5112.345, 5116.579,
  5147.761, 5145.638, 5143.153, 5141.378, 5139.235, 5135.548, 5129.865, 
    5125.833, 5121.094, 5118.429, 5119.005, 5121.696, 5125.411, 5130.348, 
    5136.462,
  5154.894, 5152.441, 5149.098, 5146.39, 5142.872, 5140.199, 5136.217, 
    5132.181, 5131.251, 5133.863, 5138.013, 5143.739, 5150.593, 5157.601, 
    5165.191,
  5161.674, 5158.97, 5155.854, 5152.372, 5149.924, 5147.106, 5145.335, 
    5146.209, 5149.542, 5155.122, 5162.599, 5170.64, 5178.512, 5186.061, 
    5193.217,
  5168.857, 5164.362, 5160.404, 5156.89, 5154.646, 5155.137, 5157.817, 
    5163.086, 5170.944, 5180.214, 5189.521, 5198.191, 5205.703, 5211.443, 
    5214.864,
  5098.555, 5105.259, 5119.336, 5133.985, 5152.921, 5167.702, 5182.573, 
    5199.529, 5212.476, 5223.112, 5233.701, 5243.813, 5250.306, 5255.726, 
    5257.58,
  5106.96, 5110.175, 5120.171, 5133.119, 5145.974, 5160.708, 5178.495, 
    5188.565, 5202.008, 5214.984, 5221.599, 5228.82, 5231.562, 5234.692, 
    5231.377,
  5113.787, 5116.162, 5122.877, 5133.28, 5144.092, 5158.282, 5164.007, 
    5184.205, 5189.892, 5198.157, 5204.603, 5208.913, 5208.748, 5205.832, 
    5200.737,
  5118.217, 5118.246, 5124.33, 5129.444, 5139.972, 5146.537, 5162.265, 
    5163.265, 5178.148, 5184.25, 5186.082, 5185.073, 5181.812, 5177.011, 
    5168.769,
  5122.119, 5120.298, 5124.051, 5128.454, 5134.974, 5143.186, 5148.007, 
    5159.549, 5162.031, 5160.201, 5165.673, 5161.026, 5157.514, 5149.583, 
    5143.567,
  5128.963, 5124.001, 5122.129, 5124.131, 5127.59, 5132.62, 5140.21, 
    5141.477, 5146.273, 5150.796, 5147.981, 5144.712, 5141.281, 5136.028, 
    5131.422,
  5135.808, 5133.25, 5128.872, 5127.749, 5128.999, 5131.692, 5133.863, 
    5137.989, 5139.426, 5139.699, 5142.643, 5143.74, 5141.897, 5137.238, 
    5130.776,
  5145.709, 5138.263, 5133.587, 5131.292, 5131.457, 5134.806, 5139.671, 
    5143.83, 5148.592, 5153.607, 5153.931, 5151.961, 5148.832, 5143.828, 
    5136.952,
  5151.497, 5148.541, 5146.763, 5146.286, 5148.941, 5154.068, 5160.802, 
    5166.769, 5167.861, 5164.348, 5160.146, 5155.379, 5150.677, 5147.344, 
    5143.194,
  5151.39, 5152.242, 5155.017, 5160.131, 5167.292, 5175.171, 5181.21, 
    5182.143, 5178.732, 5171.893, 5161.334, 5150.322, 5142.947, 5141.101, 
    5142.624,
  5163.227, 5163.681, 5167.154, 5173.262, 5180.809, 5186.954, 5192.622, 
    5198.818, 5205.626, 5215.742, 5228.882, 5243.335, 5258.786, 5274.993, 
    5292.476,
  5164.986, 5166.438, 5169.963, 5177.634, 5187.004, 5193.779, 5201.75, 
    5205.893, 5212.937, 5223.358, 5232.878, 5245.351, 5258.236, 5272.721, 
    5285.882,
  5164.946, 5167.485, 5172.138, 5180.142, 5187.588, 5197.769, 5202.633, 
    5213.163, 5217.151, 5223.039, 5231.576, 5241.426, 5252.739, 5263.504, 
    5275.63,
  5162.313, 5166.256, 5172.71, 5178.923, 5188.46, 5195.346, 5205.209, 
    5208.288, 5216.97, 5223.944, 5229.568, 5236.735, 5245.167, 5254.381, 
    5261.846,
  5158.536, 5160.812, 5170.306, 5178.277, 5186.619, 5194.117, 5199.918, 
    5207.819, 5211.654, 5212.967, 5218.625, 5221.891, 5228.671, 5233.885, 
    5242.17,
  5158.057, 5157.441, 5165.757, 5175.032, 5184.221, 5191.12, 5196.292, 
    5197.544, 5200.441, 5203.604, 5204.919, 5206.436, 5210.464, 5214.007, 
    5219.136,
  5162.809, 5157.838, 5164.128, 5174.273, 5182.487, 5188.234, 5190.174, 
    5190.53, 5187.737, 5182.15, 5179.67, 5178.886, 5181.14, 5185.227, 5191.382,
  5168.272, 5162.25, 5169.355, 5176.277, 5184.662, 5188.961, 5190.051, 
    5184.79, 5177.558, 5169.929, 5162.564, 5157.735, 5158.608, 5162.306, 
    5167.961,
  5174.474, 5178.04, 5183.854, 5192.533, 5199.237, 5201.88, 5197.746, 
    5189.201, 5175.936, 5160.528, 5147.644, 5141.273, 5139.771, 5144.171, 
    5150.369,
  5190.683, 5196.871, 5204.034, 5210.367, 5212.825, 5211.44, 5203.855, 
    5190.152, 5171.299, 5150.648, 5131.533, 5119.916, 5118.203, 5123.701, 
    5132.322,
  5280.925, 5268.982, 5259.799, 5253.287, 5248.632, 5243.238, 5237.778, 
    5234.409, 5231.646, 5231.621, 5235.208, 5241.167, 5250.329, 5261.221, 
    5276.143,
  5271.608, 5260.789, 5253.829, 5249.393, 5247.806, 5245.321, 5244.613, 
    5242.062, 5240.88, 5240.013, 5239.34, 5241.652, 5245.752, 5255.075, 
    5266.279,
  5260.241, 5251.288, 5244.333, 5242.75, 5243.91, 5246.794, 5246.462, 
    5247.465, 5246.885, 5246.199, 5245.855, 5245.577, 5247.205, 5250.767, 
    5260.484,
  5246.836, 5239.375, 5233.165, 5231.811, 5236.07, 5241.318, 5246.963, 
    5246.895, 5247.885, 5248.408, 5248.647, 5249.143, 5250.985, 5253.462, 
    5259.227,
  5233.062, 5226.293, 5221.283, 5222.186, 5227.786, 5237.706, 5241.217, 
    5247.973, 5247.533, 5247.749, 5247.008, 5246.588, 5248.282, 5251.233, 
    5257.272,
  5218.768, 5213.044, 5209.008, 5212.272, 5219.219, 5230.753, 5238.175, 
    5240.167, 5242.439, 5242.861, 5240.814, 5239.862, 5240.117, 5243.292, 
    5248.675,
  5205.698, 5201.354, 5200.544, 5208.503, 5217.851, 5228.599, 5234.514, 
    5238.812, 5237.681, 5234.041, 5229.582, 5225.748, 5223.633, 5225.524, 
    5231.789,
  5195.578, 5193.968, 5198.33, 5207.663, 5216.598, 5226.543, 5231.909, 
    5233.105, 5230.606, 5226.983, 5220.451, 5213.839, 5207.676, 5205.286, 
    5208.993,
  5190.369, 5193.062, 5202.078, 5212.464, 5222.098, 5230.167, 5232.546, 
    5231.705, 5228.278, 5223.114, 5216.11, 5206.053, 5194.956, 5186.41, 
    5185.779,
  5190.554, 5199.219, 5209.647, 5218.729, 5226.019, 5229.077, 5229.273, 
    5226.783, 5225.048, 5221.531, 5212.714, 5199.047, 5183.156, 5170.339, 
    5165.331,
  5284.223, 5292.753, 5300.054, 5303.064, 5303.104, 5302.048, 5301.346, 
    5301.06, 5296.824, 5293.356, 5293.651, 5298.333, 5304.034, 5309.219, 
    5313.639,
  5261.095, 5272.433, 5282.558, 5288.803, 5290.755, 5290.648, 5293.145, 
    5293.363, 5292.953, 5291.775, 5287.514, 5288.23, 5290.042, 5295.711, 
    5297.871,
  5237.865, 5252.467, 5264.717, 5274.755, 5278.841, 5282.836, 5281.76, 
    5288.643, 5288.876, 5289.151, 5288.013, 5285.702, 5283.598, 5281.879, 
    5282.423,
  5215.643, 5232.836, 5246.892, 5258.258, 5265.118, 5268.3, 5275.72, 
    5275.028, 5282.009, 5284.745, 5285.428, 5284.035, 5282.144, 5278.838, 
    5274.104,
  5195.825, 5213.978, 5230.551, 5243.521, 5252.38, 5258.463, 5262.128, 
    5271.781, 5275.314, 5278.531, 5281.747, 5279.083, 5274.425, 5268.629, 
    5264.305,
  5180.408, 5198.949, 5215.478, 5229.116, 5237.943, 5245.049, 5252.667, 
    5257.864, 5267.044, 5274.025, 5275.093, 5271.896, 5266.517, 5259.272, 
    5251.99,
  5168.172, 5187.63, 5204.623, 5217.853, 5227.877, 5235.694, 5243.176, 
    5252.825, 5261.653, 5267.437, 5269.54, 5266.594, 5260.763, 5251.101, 
    5239.498,
  5160.568, 5179.689, 5195.022, 5207.675, 5217.434, 5226.907, 5235.875, 
    5244.491, 5255.07, 5262.845, 5265.136, 5265.038, 5258.501, 5245.395, 
    5228.009,
  5155.269, 5174.049, 5189.504, 5202.298, 5212.533, 5221.875, 5231.618, 
    5242.625, 5252.79, 5260.051, 5265.62, 5264.907, 5255.876, 5239.815, 
    5217.98,
  5154.264, 5170.814, 5184.468, 5196.968, 5207.076, 5217.374, 5228.004, 
    5238.647, 5249.475, 5259.628, 5265.595, 5264.119, 5254.375, 5236.646, 
    5211.36,
  5224.07, 5231.092, 5242.814, 5256.864, 5271.896, 5283.762, 5292.431, 
    5300.063, 5304.688, 5306.195, 5306.774, 5304.82, 5301.457, 5299.094, 
    5299.934,
  5210.066, 5216.489, 5226.953, 5241.089, 5255.167, 5268.026, 5280.374, 
    5286.644, 5292.809, 5297.914, 5299.792, 5299.589, 5297.238, 5294.498, 
    5292.139,
  5195.246, 5202.621, 5213.088, 5227.097, 5241.858, 5256.613, 5264.759, 
    5278.927, 5283.701, 5288.276, 5292.035, 5294.312, 5293.24, 5290.286, 
    5286.298,
  5178.535, 5185.963, 5198.222, 5211.612, 5227.281, 5240.134, 5257.332, 
    5262.017, 5274.195, 5280.195, 5284.772, 5286.987, 5287.46, 5284.223, 
    5278.517,
  5163.324, 5170.114, 5182.332, 5197.751, 5213.047, 5229.935, 5240.609, 
    5258.587, 5264.683, 5270.285, 5276.654, 5279.676, 5279.91, 5275.178, 
    5268.277,
  5149.918, 5156.099, 5166.429, 5181.608, 5197.768, 5214.102, 5231.358, 
    5242.002, 5254.321, 5264.165, 5268.975, 5272.699, 5272.382, 5266.889, 
    5257.405,
  5139.286, 5146.372, 5155.593, 5168.993, 5186.031, 5202.706, 5218.104, 
    5234.927, 5246.393, 5254.716, 5262.524, 5266.621, 5265.843, 5258.944, 
    5245.394,
  5130.531, 5139.909, 5148.155, 5158.916, 5173.311, 5191.454, 5208.126, 
    5222.181, 5234.788, 5247.282, 5255.969, 5261.24, 5260.859, 5251.779, 
    5233.146,
  5124.778, 5134.888, 5144.596, 5154.921, 5167.907, 5183.689, 5199.897, 
    5215.754, 5228.479, 5240.383, 5250.845, 5258.265, 5257.64, 5245.722, 
    5222.207,
  5124.791, 5132.935, 5141.433, 5150.682, 5163.209, 5178.55, 5194.164, 
    5207.315, 5220.977, 5235.763, 5248.266, 5256.954, 5256.334, 5241.926, 
    5217.946,
  5261.351, 5232.215, 5206.916, 5188.038, 5179.811, 5181.411, 5191.453, 
    5205.039, 5221.08, 5238.297, 5255.713, 5269.536, 5278.342, 5281.751, 
    5282.405,
  5246.909, 5217.633, 5194.149, 5178.246, 5171.256, 5175.606, 5187.634, 
    5200.309, 5216.023, 5234.176, 5249.654, 5262.03, 5270.742, 5275.071, 
    5275.467,
  5231.266, 5203.673, 5183.116, 5170.54, 5166.811, 5173.343, 5181.823, 
    5199.99, 5213.651, 5229.091, 5243.532, 5255.345, 5262.695, 5266.479, 
    5267.267,
  5214.208, 5189.209, 5171.363, 5161.718, 5162.35, 5167.701, 5182.848, 
    5192.551, 5210.036, 5225.624, 5238.208, 5248.125, 5254.829, 5257.788, 
    5256.412,
  5198.398, 5176.996, 5162.311, 5155.836, 5158.6, 5167.818, 5177.844, 
    5195.77, 5209.936, 5220.577, 5233.669, 5241.584, 5247.028, 5247.771, 
    5245.375,
  5183.382, 5166.25, 5153.801, 5150.014, 5154.738, 5164.55, 5178.224, 
    5190.478, 5203.733, 5219.113, 5228.345, 5235.743, 5239.67, 5238.7, 
    5233.538,
  5171.595, 5160.349, 5150.062, 5148.397, 5153.695, 5164.464, 5175.388, 
    5191.625, 5205.233, 5215.676, 5224.496, 5231.185, 5232.822, 5230.356, 
    5220.952,
  5163.983, 5156.633, 5149.121, 5148.251, 5152.036, 5163.105, 5174.136, 
    5186.791, 5198.877, 5212.193, 5220.821, 5227.183, 5227.472, 5223.297, 
    5209.093,
  5160.325, 5155.65, 5153.222, 5149.618, 5153.049, 5161.478, 5172.292, 
    5185.883, 5198.643, 5209.926, 5218.291, 5224.083, 5224.151, 5216.205, 
    5200.155,
  5158.605, 5155.879, 5154.904, 5151.257, 5151.28, 5158.663, 5170.002, 
    5181.402, 5193.562, 5206.273, 5216.674, 5221.39, 5221.484, 5211.698, 5200,
  5329.404, 5314.024, 5296.086, 5273.505, 5248.91, 5223.325, 5200.719, 
    5185.137, 5176.155, 5176.073, 5186.512, 5208.991, 5235.299, 5255.67, 
    5271.803,
  5300.101, 5286.966, 5270.922, 5250.234, 5227.81, 5203.36, 5189.404, 
    5176.119, 5169.811, 5174.31, 5185.816, 5207.967, 5232.438, 5252.435, 
    5265.949,
  5269.369, 5259.351, 5245.31, 5229.196, 5207.465, 5194.706, 5173.106, 
    5172.772, 5167.493, 5174.267, 5186.167, 5206.829, 5229.043, 5246.141, 
    5259.214,
  5238.444, 5231.156, 5220.052, 5205.776, 5189.077, 5172.52, 5169.064, 
    5158.683, 5164.131, 5172.739, 5187, 5205.816, 5225.403, 5241.23, 5250.453,
  5214.453, 5208.575, 5200.008, 5186.958, 5173.537, 5163.874, 5155.411, 
    5160.784, 5164.599, 5172.897, 5188.01, 5204.807, 5221.643, 5233.562, 
    5241.341,
  5196.021, 5190.72, 5181.91, 5170.334, 5158.451, 5151.626, 5151.195, 
    5154.569, 5162.088, 5175.348, 5188.358, 5204.094, 5217.531, 5227.202, 
    5232.084,
  5184.492, 5177.397, 5168.784, 5157.341, 5149.664, 5146.615, 5148.63, 
    5156.866, 5167.105, 5177.347, 5190.294, 5203.322, 5214.541, 5221.106, 
    5221.707,
  5174.906, 5167.372, 5157.059, 5146.966, 5141.881, 5144.031, 5149.049, 
    5156.86, 5167.121, 5179.807, 5192.005, 5203.094, 5211.741, 5216.185, 
    5213.028,
  5166.773, 5159.101, 5150.527, 5143.182, 5141.696, 5145.615, 5151.235, 
    5161.724, 5172.839, 5183.521, 5193.762, 5203.676, 5210.312, 5211.314, 
    5206.531,
  5162.898, 5156.768, 5149.689, 5142.787, 5141.639, 5145.812, 5153.62, 
    5163.317, 5174.053, 5185.223, 5195.166, 5203.628, 5208.695, 5208.328, 
    5208.727,
  5299.877, 5282.601, 5268.4, 5254.344, 5242.774, 5231.41, 5221.241, 
    5214.553, 5209.832, 5205.539, 5205.786, 5209.023, 5218.341, 5233.542, 
    5250.92,
  5264.499, 5245.264, 5229.787, 5215.469, 5204.59, 5194.181, 5191.034, 
    5184.559, 5182.557, 5182.969, 5184.471, 5189.601, 5200.416, 5218.928, 
    5237.736,
  5229.304, 5211.25, 5195.804, 5184.011, 5175.467, 5174.316, 5164.348, 
    5168.713, 5164.54, 5165.502, 5168.014, 5174.371, 5186.153, 5204.763, 
    5226.524,
  5207.233, 5189.781, 5175.617, 5166.413, 5160.687, 5155.489, 5158.016, 
    5150.884, 5152.856, 5153.242, 5156.317, 5162.911, 5175.727, 5195.744, 
    5218.286,
  5194.023, 5178.649, 5166.063, 5156.387, 5150.901, 5148.385, 5144.308, 
    5146.864, 5143.811, 5143.204, 5148.94, 5155.831, 5170.297, 5188.708, 
    5212.271,
  5189.025, 5173.279, 5158.73, 5149.152, 5141.367, 5138.575, 5137.467, 
    5135.186, 5137.337, 5141.081, 5145.595, 5154.875, 5168.848, 5188.616, 
    5211.387,
  5188.367, 5172.499, 5157.221, 5145.969, 5138.028, 5131.881, 5128.335, 
    5129.56, 5133.187, 5138.303, 5147.238, 5158.806, 5173.668, 5192.401, 
    5213.748,
  5191.822, 5174.665, 5157.434, 5144.448, 5134.22, 5128.11, 5125.341, 
    5127.055, 5133.513, 5143.695, 5155.254, 5167.99, 5182.867, 5200.271, 
    5218.439,
  5199.071, 5182.357, 5164.514, 5150.212, 5141.174, 5134.738, 5131.53, 
    5135.375, 5142.979, 5153.261, 5165.726, 5178.491, 5192.592, 5207.811, 
    5222.838,
  5209.89, 5192.328, 5174.096, 5158.61, 5147.256, 5142.109, 5141.481, 
    5144.967, 5152.865, 5164.373, 5175.881, 5188.737, 5201.44, 5214.707, 
    5227.057,
  5290.714, 5265.595, 5242.954, 5219.83, 5199.88, 5182.759, 5168.401, 
    5160.407, 5155.033, 5149.311, 5146.408, 5145.779, 5149.804, 5159.324, 
    5174.772,
  5275.08, 5249.563, 5225.666, 5201.51, 5181.108, 5161.359, 5153.55, 
    5143.517, 5140.459, 5137.169, 5133.726, 5132.515, 5134.923, 5144.339, 
    5159.456,
  5267.179, 5242.339, 5216.998, 5193.536, 5170.531, 5156.806, 5142.132, 
    5140.553, 5136.224, 5132.599, 5127.861, 5126.593, 5128.106, 5135.194, 
    5150.536,
  5266.771, 5240.742, 5214.497, 5189.839, 5168.593, 5148.989, 5143.413, 
    5136.184, 5133.135, 5129.421, 5124.834, 5123.604, 5126.951, 5136.151, 
    5151.787,
  5271.043, 5245.254, 5219.82, 5194.994, 5173.577, 5156.274, 5142.77, 
    5138.367, 5134.571, 5129.502, 5125.338, 5125.439, 5130.619, 5140.484, 
    5157.799,
  5279.924, 5252.936, 5225.91, 5202.821, 5179.653, 5160.863, 5149.317, 
    5140.147, 5134.415, 5130.995, 5128.94, 5131.034, 5138.141, 5150.696, 
    5166.672,
  5291.735, 5266.067, 5238.228, 5215.41, 5194.715, 5175.312, 5157.396, 
    5147.48, 5139.859, 5135.017, 5134.297, 5139.071, 5147.437, 5160.696, 
    5177.071,
  5307.157, 5280.443, 5251.384, 5227.854, 5206.26, 5188.791, 5172.019, 
    5158.105, 5147.775, 5143.738, 5143.795, 5149.416, 5159.507, 5174.068, 
    5192.177,
  5324.995, 5299.105, 5270.285, 5245.259, 5224.179, 5206.66, 5189.6, 
    5176.853, 5165.697, 5159.062, 5158.409, 5164.431, 5175.52, 5191.149, 
    5210.254,
  5345.164, 5316, 5286.816, 5260.562, 5236.012, 5219.5, 5206.709, 5194.662, 
    5183.879, 5178.068, 5177.891, 5183.971, 5195.471, 5211.193, 5229.139,
  5301.953, 5271.786, 5242.655, 5212.382, 5183.648, 5157.846, 5132.897, 5117, 
    5103.785, 5090.821, 5082.248, 5076.817, 5075.032, 5079.283, 5090.469,
  5316.898, 5284.203, 5252.131, 5220.143, 5190.825, 5159.662, 5141.202, 
    5117.434, 5102.518, 5093.87, 5086.806, 5082.393, 5079.798, 5084.012, 
    5093.497,
  5335.024, 5301.002, 5266.694, 5234.693, 5200.332, 5176.776, 5143.415, 
    5129.763, 5112.869, 5099.873, 5091.737, 5088.473, 5087.063, 5090.515, 
    5100.78,
  5354.527, 5318.663, 5283.107, 5246.886, 5216.404, 5181.57, 5161.892, 
    5134.555, 5116.485, 5107.182, 5099.996, 5095.536, 5096.374, 5101.11, 
    5114.659,
  5375.239, 5339.075, 5303.296, 5265.738, 5232.904, 5201.932, 5173.193, 
    5152.478, 5138.874, 5119.824, 5114.56, 5108.676, 5112.21, 5117.062, 
    5132.385,
  5394.145, 5358.34, 5321.09, 5284.784, 5249.38, 5217.709, 5193.84, 5169.551, 
    5150.662, 5140.382, 5133.372, 5130.032, 5133.05, 5140.638, 5154.11,
  5410.727, 5378.216, 5341.966, 5305.912, 5271.626, 5239.608, 5211.939, 
    5194.126, 5178.551, 5165.798, 5157.668, 5156.271, 5158.832, 5166.965, 
    5179.1,
  5423.658, 5392.641, 5358.22, 5324.109, 5290.111, 5258.76, 5232.817, 5214.1, 
    5199.362, 5190.485, 5185.535, 5184.147, 5187.535, 5195.03, 5205.98,
  5434.565, 5405.707, 5374.673, 5342.495, 5310.74, 5280.013, 5252.26, 
    5235.581, 5224.846, 5216.115, 5211.488, 5211.582, 5214.98, 5221.677, 
    5230.385,
  5441.305, 5411.133, 5381.808, 5353.583, 5323.104, 5296.387, 5271.246, 
    5251.798, 5241.72, 5237.285, 5235.295, 5236.599, 5239.604, 5245.241, 
    5251.759,
  5277.076, 5247.836, 5216.808, 5180.212, 5144.789, 5112.677, 5080.955, 
    5059.109, 5043.912, 5030.458, 5022.54, 5017.792, 5015.929, 5017.196, 
    5024.673,
  5276.079, 5247.922, 5218.382, 5183.034, 5149.541, 5114.352, 5091.035, 
    5063.965, 5044.635, 5032.934, 5023.572, 5018.229, 5016.433, 5020.639, 
    5028.449,
  5275.671, 5249.473, 5222.779, 5190.652, 5156.547, 5133.54, 5097.035, 
    5079.865, 5060.758, 5045.458, 5034, 5028.615, 5027.687, 5032.177, 5041.015,
  5275.52, 5250.786, 5228.766, 5196.826, 5170.781, 5139.266, 5122.386, 
    5095.796, 5077.693, 5065.484, 5057.501, 5051.143, 5052.786, 5057.307, 
    5069.265,
  5275.383, 5253.47, 5236.048, 5207.536, 5184.474, 5159.991, 5139.938, 
    5119.529, 5112.008, 5093.537, 5089.276, 5082.492, 5086.608, 5088.921, 
    5100.715,
  5275.772, 5256.287, 5241.163, 5218.69, 5197.282, 5176.486, 5162.243, 
    5146.601, 5132.092, 5125.363, 5120.328, 5117.081, 5119.25, 5123.602, 
    5132.049,
  5276.582, 5260.585, 5248.171, 5231.368, 5213.914, 5198.298, 5182.669, 
    5172.565, 5164.861, 5157.797, 5152.53, 5151.91, 5153.02, 5157.118, 
    5163.034,
  5279.379, 5265.903, 5255.19, 5243.278, 5227.477, 5215.698, 5205.5, 
    5197.657, 5188.978, 5186.045, 5183.965, 5183.314, 5184.528, 5188.075, 
    5192.452,
  5284.127, 5272.947, 5263.821, 5256.408, 5244.726, 5235.72, 5225.835, 
    5221.931, 5217.916, 5214.922, 5212.625, 5213.238, 5213.977, 5216.398, 
    5218.822,
  5290.878, 5280.296, 5272.539, 5267.445, 5257.151, 5251.967, 5247.009, 
    5243.732, 5240.024, 5239.374, 5239.049, 5239.804, 5240.725, 5243.089, 
    5245.011,
  5181.213, 5165.707, 5147.877, 5124.596, 5098.744, 5070.687, 5040.175, 
    5020.875, 5006.39, 4997.396, 4996.369, 5001.143, 5008.67, 5019.099, 
    5032.034,
  5185.78, 5172.559, 5155.232, 5135.476, 5112.388, 5083.059, 5062.489, 
    5036.297, 5016.018, 5005.978, 5000.773, 5002.261, 5006.658, 5016.105, 
    5026.66,
  5194.965, 5182.864, 5167.637, 5152.509, 5127.826, 5113.97, 5078.095, 
    5063.412, 5044.352, 5026.621, 5013.227, 5008.041, 5008.537, 5014.177, 
    5023.266,
  5207.421, 5196.143, 5184.649, 5167.127, 5153.189, 5125.216, 5113.686, 
    5086.418, 5066.127, 5051.029, 5037.935, 5023.922, 5019.124, 5018.937, 
    5026.245,
  5221.472, 5211.93, 5203.301, 5188.83, 5174.386, 5156.493, 5133.798, 
    5111.339, 5099.83, 5073.503, 5061.846, 5045.642, 5037.104, 5030.146, 
    5033.904,
  5236.907, 5229.935, 5221.106, 5210.859, 5196.684, 5179.15, 5163.37, 
    5141.115, 5117.638, 5101.219, 5083.645, 5067.942, 5056.393, 5047.772, 
    5046.276,
  5253.056, 5248.203, 5240.855, 5232.852, 5222.241, 5208.303, 5188.37, 
    5170.11, 5150.764, 5128.842, 5108.544, 5091.911, 5077.341, 5067.111, 
    5062.055,
  5270.267, 5266.625, 5260.157, 5254.4, 5244.261, 5233.113, 5218.73, 
    5199.972, 5177.371, 5156.708, 5135.798, 5116.93, 5100.632, 5088.787, 
    5081.41,
  5287.468, 5284.554, 5279.844, 5275.311, 5268.991, 5258.991, 5244.539, 
    5229.816, 5211.833, 5190.079, 5166.862, 5146.459, 5128.106, 5114.115, 
    5104.545,
  5304.691, 5301.423, 5298.469, 5294.277, 5287.302, 5280.476, 5270.786, 
    5256.317, 5238.766, 5220.237, 5199.234, 5178.144, 5158.897, 5143.478, 
    5132.234,
  5205.749, 5193.532, 5179.445, 5161.033, 5140.401, 5117.3, 5088.255, 
    5063.886, 5040.306, 5018.733, 5007.248, 5004.081, 5009.648, 5025.249, 
    5057.521,
  5217.974, 5206.022, 5190.184, 5170.512, 5149.305, 5120.64, 5097.61, 
    5063.713, 5037.722, 5017.867, 5004.323, 5000.265, 5001.923, 5015.911, 
    5040.54,
  5231.077, 5220.166, 5204.024, 5186.277, 5158.966, 5139.417, 5101.046, 
    5078.111, 5049.405, 5023.958, 5005.856, 4999.877, 5000.361, 5008.289, 
    5028.614,
  5244.874, 5233.803, 5219.079, 5197.899, 5176.897, 5143.587, 5121.902, 
    5084.442, 5055.05, 5032.221, 5013.006, 5002.527, 5002.755, 5008.612, 
    5024.378,
  5256.275, 5246.324, 5233.193, 5213.017, 5190.679, 5163.384, 5130.922, 
    5102.028, 5078.166, 5043.819, 5024.608, 5008.356, 5007.37, 5008.464, 
    5022.1,
  5265.747, 5256.458, 5242.658, 5225.095, 5201.525, 5174.479, 5146.704, 
    5114.284, 5085.792, 5062.79, 5037.904, 5019.478, 5013.745, 5014.045, 
    5022.994,
  5272.661, 5264.86, 5252.042, 5235.416, 5213.76, 5187.149, 5156.807, 
    5130.768, 5107.076, 5081.318, 5056.713, 5034.785, 5022.412, 5020.045, 
    5024.157,
  5278.31, 5270.23, 5257.871, 5242.07, 5219.439, 5193.73, 5166.081, 5139.041, 
    5115.379, 5095.945, 5075.074, 5053.231, 5035.928, 5028.536, 5029.606,
  5282.304, 5274.96, 5262.767, 5247.205, 5225.574, 5199.399, 5171.586, 
    5148.961, 5128.98, 5110.901, 5090.987, 5071.273, 5053.454, 5039.604, 
    5034.933,
  5285.681, 5276.804, 5265.063, 5248.35, 5224.809, 5200.521, 5175.444, 
    5152.102, 5132.92, 5118.441, 5104.35, 5087.191, 5070.495, 5056.384, 
    5045.317,
  5207.026, 5206.018, 5201.89, 5192.436, 5179.86, 5162.428, 5140.527, 
    5120.168, 5099.689, 5079.863, 5064.806, 5053.165, 5047.684, 5046.605, 
    5054.798,
  5208.872, 5204.125, 5194.618, 5181.52, 5164.428, 5141.893, 5124.52, 
    5098.109, 5079.306, 5064.755, 5048.892, 5038.46, 5029.694, 5028.39, 
    5032.027,
  5206.172, 5197.858, 5183.958, 5168.969, 5147.061, 5131.199, 5098.546, 
    5084.953, 5064.311, 5052.116, 5037.788, 5025.804, 5015.592, 5010.864, 
    5012.654,
  5200.735, 5188.344, 5171.638, 5152.023, 5130.794, 5104.49, 5089.841, 
    5061.719, 5053.663, 5043.66, 5030.373, 5014.593, 5003.843, 4996.5, 
    4997.617,
  5193.568, 5177.947, 5159.711, 5137.519, 5115.517, 5094.081, 5069.093, 
    5060.223, 5048.595, 5038.655, 5024.634, 5006.002, 4994.068, 4984.552, 
    4985.484,
  5186.042, 5168.397, 5147.694, 5125.624, 5102.113, 5081.444, 5066.041, 
    5051.365, 5044.79, 5037.286, 5020.575, 5001.609, 4987.69, 4978.187, 
    4976.536,
  5180.286, 5162.122, 5141.185, 5119.433, 5098.429, 5078.398, 5061.954, 
    5054.792, 5048.038, 5036.928, 5020.875, 5001.164, 4985.146, 4975.674, 
    4972.411,
  5178.208, 5159.989, 5138.831, 5117.124, 5095.263, 5076.89, 5064.441, 
    5054.505, 5047.639, 5039.653, 5024.39, 5004.942, 4987.75, 4978.075, 
    4974.875,
  5180.236, 5163.01, 5142.448, 5121.256, 5100.419, 5081.877, 5067.286, 
    5060.582, 5053.672, 5044.274, 5030.518, 5012.561, 4994.616, 4984.027, 
    4981.346,
  5186.395, 5169.28, 5150.088, 5128.602, 5105.966, 5087.63, 5073.727, 
    5063.249, 5056.46, 5048.839, 5037.792, 5022.589, 5005.34, 4993.229, 
    4989.929,
  5169.21, 5166.477, 5162.876, 5158.297, 5154.098, 5149.624, 5145.339, 
    5143.601, 5140.547, 5136.88, 5134.933, 5133.12, 5131.82, 5130.841, 
    5130.922,
  5163.226, 5155.919, 5146.833, 5137.865, 5128.483, 5120.356, 5116.166, 
    5109.62, 5106.374, 5104.894, 5100.696, 5100.267, 5098.006, 5099.718, 
    5098.1,
  5153.208, 5141.942, 5127.473, 5114.59, 5099.705, 5092.96, 5077.326, 
    5078.304, 5069.716, 5068.727, 5066.91, 5067.997, 5067.292, 5067.971, 
    5068.485,
  5146.741, 5132.203, 5114.682, 5097.497, 5081.697, 5067.042, 5064.434, 
    5050.907, 5050.829, 5048.049, 5047.398, 5047.189, 5046.393, 5046, 5044.082,
  5146.613, 5130.707, 5112.276, 5092.198, 5075.696, 5063.109, 5049.763, 
    5048.396, 5040.877, 5037.964, 5037.576, 5034.446, 5031.319, 5026.28, 
    5024.013,
  5150.572, 5134.167, 5113.948, 5093.773, 5073.646, 5059.208, 5049.481, 
    5038.672, 5034.621, 5033.084, 5028.68, 5023.716, 5017.179, 5009.608, 
    5003.917,
  5157.772, 5142.156, 5121.975, 5100.334, 5080.409, 5061.788, 5047.174, 
    5039.623, 5032.055, 5025.216, 5020.398, 5013.389, 5003.746, 4993.718, 
    4985.015,
  5165.862, 5149.727, 5129.851, 5108.352, 5085.082, 5064.942, 5048.493, 
    5034.93, 5025.204, 5018.637, 5011.107, 5002.361, 4991.068, 4979.066, 
    4968.548,
  5173.159, 5157.971, 5138.818, 5117.293, 5094.298, 5071.332, 5050.824, 
    5035.55, 5022.291, 5011.073, 5001.394, 4991.141, 4978.632, 4966.145, 
    4955.288,
  5178.775, 5162.21, 5144.094, 5124.111, 5100.062, 5076.431, 5054.097, 
    5033.377, 5016.879, 5004.214, 4992.855, 4981.422, 4968.57, 4955.883, 
    4945.305,
  5176.677, 5174.774, 5172.436, 5168.506, 5163.885, 5157.759, 5151.833, 
    5149.626, 5145.755, 5141.632, 5142.724, 5146.204, 5152.428, 5159.802, 
    5170.776,
  5172.997, 5167.647, 5161.17, 5152.725, 5143.58, 5133.863, 5126.527, 
    5114.926, 5110.811, 5110.276, 5106.891, 5109.692, 5113.004, 5123.432, 
    5130.566,
  5173.832, 5167.334, 5158.632, 5149.172, 5136.616, 5126.722, 5109.558, 
    5105.577, 5089.813, 5081.65, 5077.82, 5077.139, 5078.627, 5083.71, 
    5093.238,
  5178.16, 5169.941, 5159.597, 5147.321, 5133.318, 5116.855, 5105.07, 
    5081.735, 5075.144, 5063.921, 5053.031, 5048.282, 5047.798, 5051.338, 
    5057.488,
  5181.764, 5172.605, 5161.153, 5145.903, 5128.918, 5110.528, 5088.382, 
    5074.864, 5051.791, 5038.19, 5030.298, 5021.884, 5021.786, 5020.954, 
    5028.113,
  5184.753, 5173.664, 5158.27, 5140.905, 5118.679, 5096.391, 5072.636, 
    5045.334, 5026.529, 5012.053, 4998.292, 4993.469, 4994.555, 4997.297, 
    5003.654,
  5187.003, 5173.863, 5155.532, 5133.572, 5108.75, 5079.145, 5048.737, 
    5020.182, 4992.216, 4970.474, 4960.436, 4957.865, 4961.041, 4969.314, 
    4978.635,
  5188.986, 5171.362, 5149.054, 5123.221, 5091.254, 5056.298, 5017.594, 
    4978.71, 4948.213, 4927.114, 4915.074, 4914.167, 4923.495, 4937.762, 
    4953.167,
  5189.586, 5170.719, 5145.904, 5115.021, 5078.036, 5033.466, 4983.671, 
    4941.27, 4903.599, 4877.963, 4867.857, 4872.523, 4886.357, 4906.236, 
    4926.127,
  5191.289, 5168.387, 5139.475, 5103.917, 5058.377, 5007.437, 4951.351, 
    4900.434, 4858.631, 4833.828, 4824.925, 4834.258, 4854.272, 4879.576, 
    4903.47,
  5221.204, 5219.215, 5217.509, 5217.266, 5217.519, 5217.478, 5215.975, 
    5219.054, 5217.405, 5213.406, 5212.906, 5213.454, 5213.498, 5214.994, 
    5217.69,
  5223.806, 5222.071, 5218.052, 5215.012, 5208.769, 5204.589, 5200.268, 
    5188.722, 5184.46, 5182.908, 5175.195, 5172.708, 5170.335, 5172.727, 
    5171.844,
  5230.106, 5227.7, 5221.917, 5215.686, 5205.215, 5197.289, 5179.865, 
    5179.954, 5161.855, 5151.88, 5145.066, 5140.34, 5136.092, 5135.061, 
    5137.581,
  5234.863, 5228.495, 5218.709, 5205.906, 5192.304, 5174.228, 5164.267, 
    5135.045, 5128.021, 5113.705, 5100.204, 5092.999, 5089.581, 5089.603, 
    5092.484,
  5236.061, 5226.157, 5212.754, 5195.688, 5174.237, 5154.283, 5127.425, 
    5114.936, 5084.837, 5063.354, 5050.224, 5036.559, 5033.847, 5031.51, 
    5039.73,
  5233.63, 5219.366, 5200.083, 5176.783, 5151.245, 5124.156, 5095.506, 
    5060.471, 5034.526, 5012.609, 4989.654, 4975.961, 4969.625, 4969.086, 
    4978.125,
  5229.216, 5211.201, 5186.622, 5159.78, 5128.576, 5094.137, 5057.283, 
    5023.195, 4989.057, 4959.435, 4939.426, 4922.613, 4911.79, 4909.905, 
    4917.704,
  5222.595, 5198.779, 5170.962, 5137.908, 5101.475, 5061.122, 5018.405, 
    4979.638, 4949.655, 4924.425, 4897.914, 4875.183, 4860.157, 4854.859, 
    4862.441,
  5214.409, 5189.567, 5157.275, 5119.53, 5077.868, 5031.424, 4989.052, 
    4957.514, 4924.639, 4890.745, 4859.467, 4831.384, 4810.374, 4802.063, 
    4809.179,
  5208.348, 5176.404, 5140.372, 5099.14, 5052.715, 5007.918, 4968.866, 
    4935.001, 4900.52, 4866.274, 4831.014, 4797.889, 4772.998, 4762.443, 
    4770.412,
  5300.206, 5294.299, 5288.229, 5280.356, 5271.519, 5260.518, 5245.934, 
    5236.986, 5225.402, 5210.868, 5202.72, 5197.891, 5195.594, 5196.188, 
    5200.839,
  5292.26, 5287.211, 5280.448, 5271.963, 5260.386, 5245.601, 5235.147, 
    5211.934, 5198.604, 5188.946, 5175.079, 5167.486, 5162.359, 5163.585, 
    5164.939,
  5285.209, 5280.58, 5271.962, 5262.538, 5246.159, 5234.303, 5205.354, 
    5199.122, 5172.942, 5154.94, 5141.805, 5132.183, 5124.663, 5122.552, 
    5125.196,
  5277.69, 5271.563, 5261.306, 5245.971, 5228.766, 5203.207, 5189.173, 
    5150.684, 5135.679, 5116.489, 5100.04, 5088.367, 5081.325, 5078.136, 
    5079.178,
  5270.542, 5261.544, 5248.336, 5229.809, 5205.402, 5180.545, 5146.451, 
    5130.54, 5099.598, 5072.513, 5059.277, 5042.592, 5035.976, 5028.647, 
    5031.553,
  5261.182, 5248.733, 5230.625, 5206.179, 5178.078, 5146.467, 5115.667, 
    5078.941, 5054.813, 5035.268, 5014.575, 4999.439, 4990.37, 4983.073, 
    4982.512,
  5251.204, 5234.787, 5210.601, 5183.749, 5151.183, 5114.701, 5081.548, 
    5055.279, 5026.915, 4998.669, 4979.045, 4963.158, 4951.694, 4943.787, 
    4939.634,
  5238.157, 5215.891, 5189.542, 5156.525, 5120.022, 5086.511, 5055.26, 
    5021.786, 4992.23, 4968.372, 4948.381, 4933.242, 4921.959, 4911.344, 
    4903.004,
  5222.806, 5199.342, 5168.076, 5132.888, 5097.841, 5065.295, 5032.617, 
    5000.404, 4968.372, 4943.505, 4926.929, 4913.806, 4899.879, 4884.695, 
    4870.182,
  5207.846, 5178.85, 5146.496, 5110.908, 5078.821, 5046.993, 5011.089, 
    4973.111, 4945.22, 4928.851, 4915.74, 4900.852, 4882.352, 4860.514, 
    4837.609,
  5350.989, 5355.964, 5357.429, 5353.867, 5347.85, 5338.058, 5324.455, 
    5313.105, 5295.044, 5270.035, 5246.187, 5220.782, 5195.291, 5169.375, 
    5148.402,
  5334.287, 5339.408, 5339.382, 5335.522, 5327.742, 5316.244, 5305.569, 
    5281.059, 5260.561, 5241.791, 5212.076, 5184.712, 5155.312, 5133.287, 
    5107.344,
  5316.577, 5321.747, 5319.862, 5317.191, 5306.828, 5299.45, 5273.882, 
    5267.074, 5235.318, 5206.426, 5176.985, 5147.761, 5116.62, 5090.592, 
    5066.726,
  5298.355, 5302.204, 5300.965, 5295.464, 5286.603, 5268.831, 5258.263, 
    5219.608, 5198.537, 5169.454, 5138.578, 5108.759, 5078.373, 5053.095, 
    5030.447,
  5280.176, 5283.023, 5281.553, 5275.542, 5263.8, 5249.214, 5220.683, 
    5207.621, 5172.549, 5133.554, 5105.671, 5070.289, 5043.084, 5017.12, 
    5000.405,
  5262.756, 5264.642, 5261.814, 5254.25, 5239.96, 5220.655, 5197.654, 
    5160.604, 5130.32, 5100.634, 5066.45, 5036.21, 5012.394, 4991.463, 
    4976.073,
  5248.354, 5248.671, 5243.954, 5233.366, 5217.999, 5194.455, 5166.295, 
    5139.073, 5105.604, 5067.841, 5036.305, 5009.9, 4988.003, 4969.885, 
    4954.361,
  5237.078, 5233.788, 5225.835, 5212.915, 5192.651, 5167.91, 5138.543, 
    5103.14, 5068.263, 5036.491, 5009.358, 4987.465, 4969.305, 4951.737, 
    4934.76,
  5224.616, 5219.382, 5208.619, 5191.777, 5169.761, 5141.818, 5110.889, 
    5078.124, 5043.233, 5013.233, 4990.746, 4971.641, 4952.592, 4933.157, 
    4913.713,
  5211.508, 5202.288, 5189.028, 5170.757, 5145.329, 5116.066, 5082.984, 
    5046.002, 5016.06, 4994.72, 4975.93, 4957.159, 4937.322, 4916.093, 4893.84,
  5246.489, 5260, 5274.195, 5286.835, 5299.531, 5308.977, 5318.171, 5326.925, 
    5331.749, 5331.82, 5330.799, 5325.519, 5315.507, 5300.158, 5282.018,
  5231.547, 5246.124, 5259.509, 5272.93, 5282.873, 5293.929, 5302.421, 
    5306.375, 5309.792, 5312.928, 5306.354, 5299.314, 5285.434, 5270.875, 
    5247.541,
  5212.735, 5228.574, 5242.795, 5256.345, 5267.218, 5278.337, 5280.346, 
    5292.039, 5288.39, 5286.073, 5280.765, 5270.875, 5254.031, 5234.291, 
    5210.665,
  5192.14, 5208.606, 5224.226, 5236.993, 5248.851, 5255.284, 5267.704, 
    5259.097, 5267.073, 5261.091, 5251.78, 5238.096, 5220.872, 5198.043, 
    5171.31,
  5170.477, 5186.929, 5203.246, 5216.917, 5227.987, 5237.115, 5238.081, 
    5248.321, 5239.366, 5230.64, 5223.709, 5204.454, 5185.652, 5157.104, 
    5133.61,
  5151.44, 5165.694, 5181.694, 5195.85, 5206.259, 5213.582, 5218.937, 
    5212.975, 5212.957, 5205.405, 5188.738, 5169.148, 5146.139, 5118.743, 
    5093.23,
  5136.136, 5147.065, 5161.234, 5174.055, 5184.785, 5190.858, 5193.308, 
    5195.117, 5186.629, 5172.106, 5157.187, 5133.536, 5107.394, 5079.903, 
    5053.763,
  5127.656, 5134.857, 5144.783, 5156.273, 5164.895, 5170.608, 5171.483, 
    5165.853, 5157.663, 5144.672, 5121.335, 5095.949, 5069.665, 5042.563, 
    5015.924,
  5121.689, 5128.118, 5135.603, 5143.091, 5148.604, 5151.583, 5150.466, 
    5145.591, 5131.563, 5110.492, 5087.42, 5062.138, 5033.942, 5006.214, 
    4979.304,
  5121.573, 5126.467, 5130.935, 5135.298, 5138.192, 5137.553, 5131.309, 
    5119.018, 5102.116, 5081.108, 5054.777, 5028.071, 5001.28, 4975.146, 
    4947.213,
  5070.486, 5073.565, 5080.797, 5090.636, 5104.85, 5120.699, 5140.559, 
    5165.574, 5190.327, 5210.774, 5228.364, 5244.318, 5256.688, 5268.252, 
    5278.448,
  5058.879, 5062.389, 5069.442, 5079.27, 5089.709, 5104.338, 5121.936, 
    5140.128, 5162.59, 5186.892, 5204.241, 5220.552, 5233.281, 5245.477, 
    5252.1,
  5051.671, 5055.039, 5062.383, 5072.784, 5082.998, 5097.635, 5108.03, 
    5128.365, 5142.734, 5161.459, 5179.976, 5195.785, 5208.504, 5216.599, 
    5226.062,
  5045.761, 5048.508, 5058.209, 5068.327, 5080.363, 5089.626, 5106.532, 
    5113.026, 5131.224, 5144.93, 5159.578, 5172.092, 5183.183, 5191.58, 
    5195.32,
  5041.613, 5043.901, 5054.335, 5066.537, 5078.508, 5091.508, 5099.708, 
    5112.888, 5121.675, 5130.17, 5142.517, 5149.736, 5158.386, 5161.24, 
    5166.016,
  5041.955, 5040.413, 5051.783, 5064.968, 5078.435, 5088.821, 5100.739, 
    5105.482, 5114.028, 5122.208, 5127.371, 5131.333, 5135.049, 5134.618, 
    5134.488,
  5044.365, 5041.981, 5049.704, 5063.271, 5076.849, 5087.438, 5094.679, 
    5102.232, 5106.306, 5106.908, 5109.805, 5108.988, 5107.589, 5102.983, 
    5098.198,
  5050.209, 5046.398, 5050.72, 5061.187, 5072.051, 5080.263, 5086.388, 
    5088.522, 5090.031, 5091.205, 5088.154, 5083.77, 5077.779, 5069.724, 
    5059.73,
  5059.25, 5055.692, 5055.112, 5060.345, 5066.641, 5072.294, 5074.803, 
    5076.042, 5072.992, 5067.064, 5060.603, 5052.889, 5042.475, 5030.333, 
    5016.101,
  5070.359, 5065.338, 5062.986, 5063.005, 5063.142, 5063.623, 5061.916, 
    5057.397, 5051.546, 5044.131, 5034.063, 5021.854, 5007.96, 4991.885, 
    4973.485,
  5033.944, 5017.806, 5003.918, 4992.293, 4982.29, 4974.183, 4968.271, 
    4969.061, 4976.799, 4989.065, 5006.152, 5026.237, 5045.485, 5065.402, 
    5087.038,
  5024.259, 5008.662, 4995.59, 4983.206, 4972.511, 4961.97, 4957.198, 
    4950.917, 4954.191, 4967.054, 4983.552, 5005.396, 5026.664, 5050.236, 
    5069.506,
  5019.288, 5004.672, 4992.141, 4980.878, 4968.3, 4958.402, 4945.97, 
    4944.196, 4940.91, 4947.91, 4963.314, 4985.849, 5008.832, 5031.613, 
    5054.442,
  5017.223, 5003.494, 4991.809, 4978.809, 4967.391, 4955.332, 4947.098, 
    4936.276, 4932.558, 4935.461, 4946.8, 4967.365, 4991.693, 5015.999, 
    5037.529,
  5017.44, 5004.528, 4994.105, 4981.482, 4970.748, 4959.606, 4949.243, 
    4940.472, 4935.936, 4931.302, 4939.326, 4952.923, 4976.065, 4997.716, 
    5020.508,
  5019.136, 5005.625, 4994.458, 4983.072, 4972.749, 4964.198, 4956.873, 
    4947.348, 4940.661, 4938.021, 4939.122, 4946.349, 4961.941, 4980.761, 
    4999.847,
  5022.317, 5008.912, 4996.119, 4984.402, 4974.186, 4965.849, 4959.507, 
    4955.965, 4951.886, 4947.147, 4945.596, 4948.063, 4955.53, 4967.102, 
    4980.73,
  5028.324, 5012.341, 4996.805, 4983.253, 4970.625, 4961.466, 4956.495, 
    4952.8, 4950.504, 4950.325, 4949.74, 4950.171, 4951.547, 4955.576, 
    4961.351,
  5035.765, 5019.423, 5001.088, 4984.431, 4968.211, 4956.52, 4948.789, 
    4945.82, 4944.181, 4942.624, 4941.637, 4941.616, 4941.626, 4942.152, 
    4942.655,
  5044.276, 5025.252, 5005.7, 4986.743, 4967.852, 4953.366, 4943.768, 
    4937.36, 4933.734, 4931.682, 4929.492, 4926.797, 4923.136, 4919.119, 
    4914.616,
  5075.027, 5068.882, 5062.326, 5053.927, 5044.554, 5031.743, 5014.509, 
    5000.851, 4985.784, 4969.611, 4959.016, 4951.369, 4945.744, 4942.164, 
    4941.431,
  5062.641, 5056.536, 5049.079, 5039.353, 5027.36, 5009.977, 4997.31, 
    4974.658, 4959.877, 4948.246, 4935.321, 4927.317, 4919.914, 4917.646, 
    4913.404,
  5053.876, 5046.534, 5037.188, 5027.559, 5011.063, 4998.722, 4971.464, 
    4964.446, 4943.455, 4929.479, 4915.593, 4907.286, 4898.439, 4893.311, 
    4890.701,
  5045.617, 5037.841, 5028.183, 5014.498, 4997.562, 4975.525, 4964.341, 
    4938.906, 4928.728, 4917.004, 4902.817, 4891.38, 4881.697, 4875.509, 
    4870.874,
  5037.938, 5030.011, 5020.686, 5005.111, 4986.577, 4966.91, 4944.408, 
    4936.06, 4920.797, 4904.449, 4893.368, 4879.067, 4869.684, 4861.02, 
    4858.698,
  5029.316, 5022.878, 5012.805, 4997.693, 4977.343, 4955.191, 4937.924, 
    4918.303, 4906.849, 4898.262, 4883.683, 4870.32, 4859.738, 4852.511, 
    4849.948,
  5020.304, 5015.663, 5006.887, 4994.852, 4974.443, 4949.83, 4928.349, 
    4915.586, 4901.959, 4886.708, 4874.192, 4861.641, 4850.992, 4845.201, 
    4843.831,
  5012.272, 5009.162, 5003.2, 4990.672, 4967.947, 4944.434, 4923.143, 
    4904.009, 4888.2, 4876.204, 4862.273, 4850.253, 4841.06, 4835.163, 4834.95,
  5004.723, 5002.777, 4997.598, 4985.499, 4967.295, 4942.983, 4919.515, 
    4900.333, 4881.603, 4863.218, 4847.268, 4834.556, 4825.357, 4821.519, 
    4822.884,
  5003.381, 4999.12, 4994.162, 4983.373, 4963.901, 4942.129, 4918.021, 
    4893.616, 4871.179, 4850.89, 4831.959, 4816.227, 4805.233, 4800.321, 
    4802.162,
  5078.076, 5088.17, 5098.341, 5106.371, 5113.229, 5117.208, 5119.141, 
    5119.875, 5114.986, 5105.646, 5095.616, 5084.51, 5072.472, 5061.064, 
    5051.945,
  5058.603, 5066.913, 5074.988, 5082.759, 5087.475, 5091.922, 5094.613, 
    5090.214, 5084.989, 5079.707, 5066.433, 5055.145, 5041.863, 5033.732, 
    5022.043,
  5047.484, 5053.487, 5058.773, 5064.987, 5067.855, 5074.227, 5065.905, 
    5070.747, 5057.78, 5048.113, 5036.51, 5025.069, 5011.575, 5000.425, 
    4991.459,
  5040.892, 5045.021, 5048.432, 5051.197, 5052.796, 5049.796, 5053.727, 
    5036.703, 5033.745, 5021.921, 5006.118, 4991.342, 4977.32, 4965.04, 
    4953.34,
  5037.441, 5040.042, 5041.827, 5042.375, 5041.942, 5038.813, 5028.338, 
    5024.853, 5005.619, 4986.982, 4973.22, 4952.204, 4936.676, 4919.599, 
    4910.032,
  5037.642, 5036.922, 5035.381, 5033.308, 5027.395, 5021.144, 5011.345, 
    4991.472, 4973.907, 4954.183, 4929.738, 4907.71, 4889.083, 4872.378, 
    4862.059,
  5041.148, 5038.402, 5033.144, 5028.02, 5020.202, 5008.255, 4990.795, 
    4971.958, 4946.36, 4918.154, 4894.025, 4869.769, 4848.348, 4831.869, 
    4821.594,
  5049.535, 5043.188, 5035.259, 5026.338, 5012.307, 4995.973, 4975.28, 
    4949.693, 4923.504, 4897.301, 4868.286, 4840.542, 4816.343, 4798.064, 
    4788.062,
  5061.209, 5052.869, 5041.754, 5029.4, 5013.41, 4994.213, 4971.441, 4946.53, 
    4916.546, 4882.969, 4850.478, 4818.382, 4790.266, 4770.148, 4759.896,
  5075.93, 5064.222, 5051.691, 5037.286, 5018.63, 4998.426, 4973.644, 
    4943.603, 4911.607, 4876.9, 4840.899, 4805.164, 4774.208, 4751.412, 
    4739.828,
  5051.277, 5057.664, 5072.805, 5092.708, 5116.441, 5137.491, 5158.846, 
    5179.927, 5198.32, 5213.203, 5225.749, 5235.376, 5240.582, 5242.003, 
    5240.519,
  5052.652, 5058.632, 5067.631, 5085.196, 5104, 5124.311, 5144.148, 5160.524, 
    5176.511, 5193.561, 5202.585, 5210.558, 5212.122, 5213.859, 5206.857,
  5053.278, 5058.651, 5065.979, 5078.542, 5092.965, 5113.979, 5123.055, 
    5147.269, 5156.384, 5166.896, 5174.659, 5179.793, 5179.627, 5176.29, 
    5171.166,
  5052.842, 5056.048, 5062.509, 5069.528, 5082.419, 5090.925, 5111.885, 
    5111.826, 5131.306, 5141.206, 5145.966, 5148.205, 5147.359, 5143.761, 
    5134.639,
  5053.485, 5053.091, 5057.744, 5063.368, 5071.638, 5082.919, 5088.894, 
    5103.596, 5109.774, 5109.048, 5118.453, 5116.464, 5116.409, 5108.838, 
    5103.348,
  5056.188, 5051.971, 5050.701, 5053.877, 5058.564, 5064.701, 5074.101, 
    5075.453, 5082.251, 5091.481, 5091.598, 5090.96, 5088.904, 5081.874, 
    5073.396,
  5061.827, 5055.771, 5051.078, 5048.688, 5051.678, 5055.906, 5060.229, 
    5067.632, 5070.948, 5069.264, 5070.183, 5068.305, 5062.965, 5054.808, 
    5043.839,
  5066.896, 5060.329, 5054.549, 5052.292, 5049.52, 5049.688, 5051.016, 
    5050.642, 5051.289, 5053.364, 5050.801, 5045.575, 5038.308, 5028.071, 
    5015.418,
  5065.928, 5058.871, 5052.36, 5047.71, 5044.843, 5043.465, 5041.646, 
    5041.314, 5038.166, 5032.479, 5027.105, 5020.213, 5010.197, 4998.611, 
    4984.798,
  5061.404, 5051.074, 5042.262, 5036.619, 5031.259, 5027.274, 5023.356, 
    5017.818, 5012.812, 5007.985, 5000.621, 4990.888, 4979.342, 4966.988, 
    4953.005,
  5061.824, 5049.009, 5039.227, 5034.908, 5031.499, 5029.071, 5029.516, 
    5038.226, 5051.409, 5068.461, 5091.699, 5122.748, 5157.716, 5189.366, 
    5217.708,
  5061.49, 5050.657, 5042.122, 5040.246, 5040.291, 5039.406, 5043.341, 
    5050.098, 5063.867, 5086.187, 5112.036, 5145.046, 5175.969, 5206.084, 
    5231.269,
  5061.16, 5051.625, 5045.234, 5045.228, 5047.994, 5052.059, 5055.033, 
    5068.76, 5085.511, 5104.863, 5132.993, 5162.825, 5190.971, 5214.861, 
    5238.443,
  5059.913, 5050.759, 5048.36, 5047.028, 5054.971, 5057.713, 5070.633, 
    5077.617, 5097.132, 5119.778, 5148.419, 5174.762, 5199.656, 5222.926, 
    5241.426,
  5058.949, 5048.824, 5047.481, 5048.312, 5055.369, 5066.84, 5075.633, 
    5091.418, 5114.362, 5131.054, 5157.053, 5179.421, 5202.453, 5219.954, 
    5236.099,
  5058.879, 5048.755, 5043.351, 5045.862, 5052.892, 5063.225, 5079.824, 
    5094.368, 5108.862, 5134.636, 5154.852, 5177.182, 5196.79, 5213.531, 
    5226.51,
  5055.736, 5048.459, 5042.379, 5040.848, 5046.116, 5057.312, 5070.758, 
    5089.563, 5110.585, 5127.437, 5147.918, 5167.18, 5183.797, 5197.626, 
    5207.971,
  5051.571, 5045.696, 5039.841, 5037.758, 5038.652, 5045.298, 5058.754, 
    5072.897, 5089.864, 5111.707, 5131.654, 5148.923, 5165.527, 5178.257, 
    5187.82,
  5039.703, 5034.625, 5030.537, 5028.564, 5027.679, 5032.603, 5041.35, 
    5057.084, 5074.262, 5091.034, 5107.984, 5126.141, 5141.598, 5154.242, 
    5163.354,
  5025.468, 5019.47, 5014.313, 5013.107, 5013.568, 5016.1, 5022.251, 
    5033.424, 5047.9, 5066.029, 5084.123, 5101.133, 5116.369, 5129.458, 
    5138.821,
  5106.018, 5095.672, 5084.41, 5072.747, 5060.401, 5046.901, 5029.889, 
    5018.1, 5009.977, 5006.869, 5011.451, 5023.024, 5040.246, 5058.782, 
    5077.641,
  5094.265, 5083.924, 5072.589, 5061.95, 5050.234, 5034.628, 5020.307, 
    5005.615, 4999.447, 5002.936, 5012.787, 5030.624, 5050.342, 5071.931, 
    5092.319,
  5084.5, 5075.249, 5065.26, 5056.539, 5043.77, 5031.953, 5009.729, 5004.521, 
    5001.924, 5008.464, 5023.344, 5044.408, 5066.196, 5087.894, 5115.283,
  5075.817, 5067.337, 5058.888, 5049.907, 5041.177, 5024.665, 5013.808, 
    4999.987, 5004.157, 5018.755, 5041.078, 5063.256, 5087.746, 5116.567, 
    5146.366,
  5066.528, 5060.062, 5054.047, 5047.026, 5041.024, 5027.688, 5014.838, 
    5007.591, 5024.565, 5035.412, 5062.129, 5085.105, 5115.524, 5143.895, 
    5171.815,
  5055.465, 5051.112, 5047.387, 5042.813, 5038.074, 5030.572, 5020.811, 
    5021.43, 5029.161, 5057.717, 5082.709, 5110.551, 5141.758, 5170.594, 
    5193.587,
  5042.685, 5041.193, 5040.008, 5039.227, 5037.796, 5035.022, 5027.665, 
    5033.283, 5054.363, 5078.184, 5104.535, 5134.413, 5164.029, 5189.298, 
    5209.659,
  5027.379, 5026.616, 5028.573, 5032.006, 5032.515, 5034.402, 5036.042, 
    5042.549, 5063.796, 5092.934, 5122.393, 5151.916, 5181.074, 5204.067, 
    5221.939,
  5009.606, 5007.442, 5012.382, 5022.038, 5029.307, 5033.991, 5038.155, 
    5051.977, 5079.538, 5106.833, 5135.067, 5165.291, 5191.669, 5212.625, 
    5228.149,
  4987.762, 4981.145, 4987.166, 5000.068, 5013.198, 5025.295, 5036.531, 
    5051.763, 5079.116, 5110.347, 5141.061, 5171.36, 5196.999, 5217.342, 
    5230.257,
  5097.769, 5083.916, 5074.954, 5072.387, 5071.059, 5069.216, 5067.02, 
    5066.809, 5065.781, 5064.901, 5066.174, 5071.089, 5078.797, 5088.789, 
    5099.886,
  5089.184, 5071.64, 5061.695, 5059.188, 5058.962, 5059.113, 5057.879, 
    5054.269, 5050.983, 5049.481, 5050.635, 5057.207, 5067.763, 5081.398, 
    5093.263,
  5081.439, 5058.674, 5048.444, 5046.751, 5048.818, 5051.438, 5046.383, 
    5044.379, 5038.723, 5036.369, 5039.823, 5050.033, 5064.066, 5078.515, 
    5094.625,
  5071.823, 5045.927, 5033.678, 5031.387, 5037.704, 5038.915, 5042.295, 
    5032.773, 5031.359, 5029.964, 5039.237, 5051.421, 5069.04, 5089.259, 
    5106.641,
  5062.818, 5031.624, 5017.888, 5018.208, 5027.834, 5034.365, 5032.182, 
    5032.333, 5029.683, 5033.585, 5045.957, 5063.116, 5086.786, 5105.887, 
    5119.461,
  5054.935, 5018.525, 5001.881, 5005.126, 5017.262, 5027.512, 5029.334, 
    5029.936, 5032.27, 5044.041, 5060.484, 5084.754, 5107.316, 5122.87, 
    5129.806,
  5047.731, 5008.4, 4990.483, 4997.387, 5013.272, 5024.616, 5026.784, 
    5032.664, 5042.173, 5058.733, 5081.834, 5106.826, 5125.958, 5136.651, 
    5138.499,
  5043.014, 5001.252, 4982.637, 4992.699, 5009.257, 5022.148, 5027.354, 
    5036.629, 5052.632, 5076.816, 5103.69, 5128.198, 5143.7, 5150.511, 
    5147.788,
  5041.034, 4997.054, 4980.158, 4993.588, 5011.798, 5023.633, 5030.462, 
    5046.501, 5068.872, 5096.796, 5124.961, 5147.503, 5159.931, 5164.473, 
    5159.152,
  5041.976, 4995.66, 4979.42, 4993.293, 5011.966, 5025.446, 5036.307, 
    5056.855, 5083.553, 5115.083, 5143.716, 5164.923, 5176.766, 5179.122, 
    5173.519,
  5104.166, 5062.714, 5033.79, 5022.152, 5024.423, 5032.058, 5034.106, 
    5037.114, 5038.078, 5038.003, 5038.354, 5039.276, 5041.406, 5045.388, 
    5053.957,
  5109.419, 5068.773, 5040.826, 5029.643, 5032.335, 5035.19, 5038.019, 
    5036.225, 5036.002, 5036.912, 5037.609, 5039.234, 5041.973, 5046.323, 
    5052.001,
  5118.586, 5079.173, 5052.56, 5041.579, 5040.266, 5045.76, 5040.312, 
    5039.075, 5036.684, 5035.623, 5036.87, 5039.711, 5043.039, 5047.284, 
    5053.164,
  5129.186, 5092.563, 5068.099, 5053.617, 5053.654, 5048.892, 5048.637, 
    5039.897, 5034.791, 5033.569, 5035.344, 5037.807, 5042.683, 5047.341, 
    5053.811,
  5143.292, 5108.242, 5086.519, 5071.13, 5067.224, 5062.686, 5053.997, 
    5045.417, 5039.005, 5034.567, 5037.125, 5040.311, 5047.06, 5051.217, 
    5057.704,
  5160.547, 5123.891, 5104.237, 5090.337, 5082.762, 5074.498, 5066.369, 
    5056.02, 5049.658, 5048.342, 5049.837, 5052.6, 5056.171, 5059.375, 
    5062.046,
  5179.126, 5140.481, 5122.878, 5109.522, 5100.321, 5091.321, 5079.866, 
    5072.054, 5067.015, 5063.725, 5062.342, 5063.046, 5063.729, 5066.519, 
    5069.551,
  5200.032, 5158.16, 5137.854, 5126.781, 5115.528, 5106.773, 5097.093, 
    5088.323, 5079.674, 5074.987, 5072.031, 5071.526, 5072.499, 5075.976, 
    5081.536,
  5220.092, 5178.618, 5153.997, 5141.757, 5131.946, 5124.434, 5115.271, 
    5107.626, 5098.543, 5090.917, 5085.106, 5084.293, 5087.097, 5093.424, 
    5101.302,
  5238.085, 5196.833, 5167.914, 5153.802, 5144.08, 5138.917, 5133.722, 
    5126.513, 5116.116, 5109.011, 5104.494, 5104.872, 5108.47, 5115.217, 
    5122.271,
  5272.583, 5238.435, 5203.131, 5166.612, 5134.628, 5111.873, 5094.193, 
    5085.696, 5079.112, 5070.026, 5062.96, 5055.397, 5049.953, 5044.99, 
    5044.802,
  5288.412, 5255.5, 5220.438, 5183.454, 5149.308, 5117.156, 5104.603, 
    5089.401, 5080.996, 5075.129, 5067.371, 5060.609, 5054.062, 5047.809, 
    5044.109,
  5304.924, 5273.691, 5239.087, 5204.547, 5164.261, 5139.943, 5107.375, 
    5101.013, 5089.455, 5082.234, 5073.51, 5066.702, 5059.117, 5054.32, 
    5049.294,
  5319.131, 5288.749, 5257.388, 5221.117, 5186.357, 5147.051, 5127.31, 
    5106.385, 5095.624, 5089.023, 5081.572, 5073.711, 5066.836, 5060.673, 
    5055.733,
  5333.388, 5303.133, 5274.186, 5239.036, 5205.525, 5169.429, 5138.181, 
    5120.129, 5110.528, 5098.379, 5092.481, 5083.545, 5077.726, 5068.999, 
    5063.788,
  5345.072, 5315.392, 5286.234, 5254.353, 5220.84, 5186.26, 5154.684, 
    5130.847, 5116.608, 5109.56, 5102.938, 5095.606, 5089.244, 5081.473, 
    5074.358,
  5354.065, 5327.549, 5298.786, 5267.711, 5236.133, 5203.797, 5171.704, 
    5145.438, 5131.278, 5121.017, 5114.088, 5108.417, 5101.539, 5093.842, 
    5085.22,
  5359.806, 5335.983, 5307.314, 5277.503, 5245.515, 5214.59, 5185.375, 
    5158.532, 5139.6, 5130.388, 5124.072, 5118.506, 5112.317, 5104.272, 
    5093.704,
  5362.716, 5342.052, 5315.307, 5284.619, 5253.594, 5223.235, 5194.856, 
    5170.104, 5151.496, 5139.961, 5132.434, 5126.903, 5120.165, 5111.245, 
    5099.395,
  5364.069, 5341.626, 5314.793, 5285.719, 5253.037, 5222.488, 5197.158, 
    5174.158, 5155.256, 5144.089, 5137.145, 5131.206, 5124.228, 5114.642, 
    5101.046,
  5409.601, 5384.834, 5354.381, 5322.114, 5290.472, 5259.274, 5225.589, 
    5201.287, 5175.863, 5147.022, 5125.797, 5107.054, 5092.953, 5080.219, 
    5073.162,
  5410.117, 5384.368, 5354.493, 5322.779, 5290.304, 5253.674, 5227.46, 
    5186.274, 5161.4, 5141.836, 5119.873, 5103.19, 5089.423, 5078.615, 
    5069.913,
  5409.302, 5383.102, 5352.979, 5321.835, 5284.712, 5256.106, 5209.561, 
    5190.404, 5152.117, 5127.068, 5110.168, 5097.046, 5085.034, 5075.635, 
    5067.123,
  5406.614, 5378.407, 5348.561, 5313.021, 5275.65, 5231.878, 5200.657, 
    5151.52, 5129.131, 5106.47, 5093.186, 5085.045, 5080.109, 5073.034, 
    5066.05,
  5403.285, 5374.588, 5342.802, 5304.007, 5262.136, 5216.207, 5167.702, 
    5137.46, 5103.021, 5080.323, 5073.448, 5069.24, 5071.269, 5068.474, 
    5065.042,
  5398.494, 5367.713, 5331.005, 5288.913, 5240.099, 5187.809, 5140.154, 
    5094.252, 5064.681, 5051.121, 5044.037, 5049.579, 5057.298, 5061.866, 
    5062.343,
  5393.086, 5361.363, 5320.88, 5273.434, 5217.911, 5160.677, 5107.212, 
    5066.058, 5036.109, 5019.187, 5019.267, 5029.064, 5040.833, 5051.191, 
    5054.879,
  5387.631, 5351.443, 5305.632, 5252.219, 5188.816, 5126.894, 5071.511, 
    5025.487, 4998.223, 4989.812, 4994.52, 5008.644, 5025.87, 5039.241, 
    5045.665,
  5382.403, 5345.412, 5296.921, 5236.681, 5168.875, 5100.475, 5040.916, 
    4999.472, 4974.357, 4965.645, 4975.62, 4994.295, 5012.895, 5026.991, 
    5033.912,
  5377.979, 5334.979, 5279.88, 5214.803, 5139.501, 5070.24, 5015.231, 
    4973.682, 4951.655, 4950.904, 4965.1, 4985.045, 5003.19, 5016.219, 
    5021.487,
  5346.058, 5295.255, 5243.748, 5192.291, 5145.1, 5098.292, 5046.657, 
    5011.37, 4983.521, 4957.521, 4948.878, 4951.78, 4963.781, 4981.077, 
    5003.088,
  5348.996, 5296.648, 5240.183, 5185.396, 5134.771, 5076.273, 5035.226, 
    4975.2, 4942.365, 4926.328, 4916.952, 4920.889, 4932.8, 4956.763, 4979.138,
  5355.167, 5302.137, 5241.625, 5185.601, 5125.519, 5081.961, 5009.867, 
    4979.775, 4933.995, 4907.019, 4894.612, 4898.893, 4912.118, 4935.409, 
    4963.32,
  5362.916, 5307.974, 5246.944, 5184.256, 5129.608, 5066.78, 5026.263, 
    4961.57, 4922.312, 4900.114, 4887.33, 4888.407, 4903.951, 4928.875, 
    4956.749,
  5371.941, 5317.738, 5256.543, 5192.727, 5137.668, 5082.916, 5026.682, 
    4978.184, 4941.226, 4904.081, 4893.697, 4891.532, 4908.819, 4931.2, 
    4959.849,
  5380.666, 5327.923, 5266.265, 5204.911, 5148.315, 5097.819, 5047.339, 
    4992.838, 4948.334, 4922.756, 4908.716, 4908.676, 4924.783, 4947.438, 
    4969.517,
  5390.568, 5341.65, 5283.052, 5222.195, 5169.169, 5120.999, 5068.993, 
    5023.208, 4982.418, 4949.543, 4933.88, 4934.561, 4946.861, 4965.487, 
    4980.503,
  5400.542, 5353.853, 5298.46, 5240.278, 5186.218, 5141.639, 5096.072, 
    5049.276, 5008.773, 4980.917, 4965.384, 4963.398, 4972.117, 4983.93, 
    4991.948,
  5409.808, 5367.601, 5317.428, 5261.288, 5210.1, 5166.16, 5122.299, 
    5082.387, 5046.95, 5016.253, 4998.181, 4992.763, 4994.47, 4998.339, 
    5000.099,
  5417.346, 5376.428, 5329.922, 5278.584, 5225.724, 5183.916, 5145.449, 
    5106.036, 5072.292, 5045.5, 5026.466, 5016.207, 5010.872, 5006.836, 
    5001.066,
  5417.716, 5384.351, 5350.047, 5311.114, 5272.017, 5231.913, 5187.29, 
    5150.679, 5111.872, 5070.562, 5039.029, 5014, 4998.613, 4990.369, 4991.618,
  5418.924, 5387.547, 5355.4, 5320.27, 5284.99, 5242.818, 5211.121, 5163.681, 
    5125.612, 5092.36, 5059.732, 5032.624, 5010.532, 4998.622, 4992.176,
  5417.679, 5388.421, 5357.437, 5327.329, 5290.253, 5263.296, 5212.939, 
    5188.47, 5151.223, 5114.639, 5080.157, 5051.982, 5027.126, 5010.23, 
    4998.976,
  5410.849, 5382.968, 5355.231, 5324.975, 5295.816, 5259.349, 5235.005, 
    5193.292, 5160.112, 5130.322, 5098.536, 5069.63, 5043.794, 5023.87, 
    5009.873,
  5401.409, 5375.23, 5349.93, 5321.81, 5295.254, 5266.202, 5233.028, 
    5207.503, 5177.385, 5139.716, 5112.055, 5082.168, 5058.172, 5035.515, 
    5020.353,
  5387.423, 5362.811, 5337.823, 5313.543, 5287.423, 5261.235, 5235.97, 
    5202.977, 5172.181, 5146.558, 5118.46, 5090.856, 5065.684, 5043.657, 
    5026.565,
  5370.809, 5348.491, 5324.534, 5302.014, 5279.122, 5255.615, 5229.43, 
    5205.767, 5178.517, 5148.224, 5119.9, 5093.531, 5067.287, 5045.348, 
    5026.709,
  5351.991, 5329.387, 5306.145, 5286.097, 5263.605, 5243.265, 5220.91, 
    5195.368, 5168.858, 5144.948, 5117.984, 5090.619, 5064.149, 5041.536, 
    5022.294,
  5332.151, 5310.146, 5288.787, 5268.769, 5249.292, 5230.03, 5209.214, 
    5188.986, 5165.28, 5138.889, 5110.978, 5083.545, 5056.396, 5033.705, 
    5013.423,
  5312.89, 5288.197, 5267.493, 5249.511, 5230.867, 5213.622, 5195.863, 
    5174.612, 5152.378, 5129.412, 5102.422, 5073.313, 5046.21, 5023.033, 
    5002.068,
  5323.524, 5290.958, 5262.263, 5237.886, 5220.254, 5205.839, 5192.206, 
    5184.491, 5177.089, 5166.431, 5158.817, 5150.649, 5141.177, 5129.247, 
    5118.006,
  5320.211, 5285.875, 5255.628, 5229.254, 5208.902, 5190.29, 5182.103, 
    5166.773, 5159.652, 5155.484, 5147.96, 5141.051, 5132.36, 5123.278, 
    5110.887,
  5320.779, 5285.319, 5253.834, 5227.085, 5202.11, 5188.459, 5164.42, 
    5162.082, 5148.158, 5140.829, 5134.613, 5129.569, 5121.382, 5111.963, 
    5101.361,
  5323.241, 5287.051, 5254.747, 5224.79, 5200.636, 5174.911, 5163.566, 
    5140.381, 5135.184, 5128.972, 5121.347, 5116.094, 5109.626, 5101.901, 
    5089.591,
  5327.715, 5291.607, 5259.094, 5228.422, 5201.632, 5177.197, 5152.816, 
    5139.944, 5124.414, 5113.166, 5108.71, 5101.681, 5096.996, 5087.743, 
    5078.429,
  5332.116, 5295.949, 5262.545, 5232.282, 5202.486, 5175.854, 5152.646, 
    5129.269, 5113.223, 5103.817, 5095.027, 5089.109, 5083.782, 5075.454, 
    5064.353,
  5336.12, 5302.283, 5269.025, 5238.84, 5209.229, 5180.625, 5152.965, 
    5131.336, 5110.158, 5093.277, 5083.477, 5076.775, 5069.561, 5060.77, 
    5048.426,
  5340.212, 5306.781, 5273.436, 5243.896, 5212.502, 5184.396, 5156.388, 
    5129.479, 5105.41, 5088.012, 5073.47, 5063.989, 5056.108, 5045.61, 
    5032.147,
  5344.177, 5312.643, 5280.691, 5251.112, 5221.412, 5191.991, 5161.823, 
    5134.929, 5107.84, 5084.935, 5065.987, 5052.603, 5039.665, 5028.218, 
    5015.916,
  5346.515, 5314.386, 5283.706, 5255.117, 5224.403, 5195.775, 5166.814, 
    5136.718, 5108.684, 5083.951, 5061.383, 5042.277, 5028.285, 5016.791, 
    5008.154,
  5347.691, 5319.251, 5293.052, 5268.705, 5247.098, 5226.345, 5203.96, 
    5186.632, 5167.684, 5148.247, 5135.462, 5128.772, 5129.159, 5132.512, 
    5137.528,
  5347.757, 5317.707, 5291.268, 5266.395, 5246.115, 5222.797, 5207.618, 
    5181.719, 5161.685, 5144.878, 5128.748, 5118.591, 5116.179, 5120.143, 
    5124.623,
  5347.149, 5316.474, 5289.211, 5265.785, 5242.888, 5228.163, 5201.922, 
    5188.51, 5165.642, 5142.965, 5123.988, 5110.862, 5104.343, 5106.541, 
    5112.451,
  5345.059, 5312.917, 5285.214, 5260.359, 5239.669, 5218.342, 5206.495, 
    5182.271, 5161.38, 5143.113, 5121.7, 5105.98, 5097.107, 5096.127, 5099.531,
  5342.505, 5309.36, 5281.497, 5256.672, 5236.187, 5217.653, 5199.757, 
    5186.216, 5168.112, 5141.448, 5121.961, 5102.49, 5092.422, 5086.775, 
    5090.106,
  5338.309, 5303.484, 5274.166, 5250.539, 5229.118, 5210.939, 5197.295, 
    5179.756, 5162.081, 5143.777, 5122.153, 5102.678, 5089.834, 5082.331, 
    5081.446,
  5332.133, 5298.009, 5268.027, 5244.643, 5224.073, 5207.145, 5191.44, 
    5180.327, 5164.927, 5144.604, 5123.043, 5103.382, 5087.35, 5077.932, 
    5072.857,
  5324.346, 5289.042, 5258.165, 5235.767, 5215.167, 5199.554, 5185.697, 
    5172.012, 5157.26, 5142.729, 5123.712, 5104.037, 5086.703, 5073.96, 
    5065.193,
  5315.161, 5281.084, 5251.404, 5228.305, 5208.801, 5193.483, 5179.366, 
    5168.424, 5154.245, 5137.954, 5120.722, 5102.763, 5085.326, 5070.638, 
    5058.09,
  5305.031, 5269.49, 5240.029, 5219.088, 5199.779, 5184.379, 5170.988, 
    5156.867, 5142.585, 5129.042, 5113.889, 5098.339, 5081.702, 5067.141, 
    5054.572,
  5307.778, 5269.66, 5240.018, 5219.187, 5204.417, 5189.23, 5174.527, 
    5168.746, 5166.813, 5160.299, 5151.858, 5137.5, 5123.04, 5110.836, 
    5107.983,
  5313.324, 5271.022, 5240.906, 5217.633, 5203.723, 5185.231, 5175.259, 
    5163.299, 5161.655, 5156.939, 5149.02, 5136.623, 5122.533, 5110.136, 
    5103.592,
  5318.486, 5272.891, 5242.452, 5218.625, 5203.159, 5189.93, 5171.738, 
    5166.004, 5160.65, 5154.506, 5146.347, 5135.381, 5122.598, 5109.464, 
    5101.237,
  5322.819, 5273.691, 5242.178, 5216.773, 5202.822, 5185.301, 5175.372, 
    5161.456, 5156.117, 5150.204, 5142.57, 5132.734, 5122.003, 5110.302, 
    5100.479,
  5325.919, 5274.518, 5242.87, 5216.622, 5202.07, 5187.586, 5173.579, 
    5163.223, 5155.176, 5146.554, 5138.584, 5128.052, 5119.031, 5108.599, 
    5100.443,
  5326.182, 5273.042, 5240.022, 5214.229, 5198.313, 5183.608, 5172.879, 
    5159.478, 5150.22, 5140.973, 5132.11, 5121.874, 5113.138, 5104.158, 
    5097.115,
  5323.425, 5273.082, 5239.083, 5213.418, 5196.314, 5181.696, 5169.162, 
    5157.52, 5146.278, 5134.434, 5123.781, 5113.189, 5103.649, 5095.691, 
    5089.545,
  5319.577, 5269.941, 5234.702, 5209.64, 5190.709, 5175.696, 5163.26, 
    5150.024, 5137.006, 5124.736, 5112.294, 5101.264, 5091.546, 5084.189, 
    5078.63,
  5315.706, 5267.988, 5234.304, 5207.982, 5188.124, 5171.646, 5156.951, 
    5142.761, 5127.884, 5112.747, 5098.724, 5086.419, 5076.007, 5069.213, 
    5064.471,
  5310.582, 5262.147, 5228.536, 5203.438, 5181.867, 5163.378, 5147.936, 
    5131.049, 5114.593, 5097.962, 5082.4, 5068.733, 5057.936, 5051.244, 
    5047.574,
  5336.96, 5293.757, 5256.798, 5226.369, 5202, 5182.56, 5164.37, 5153.049, 
    5144.915, 5136.152, 5131.636, 5125.979, 5120.909, 5113.726, 5106.691,
  5337.541, 5292.789, 5255.078, 5223.566, 5199.4, 5175.517, 5163.983, 
    5144.909, 5136.878, 5130.493, 5124.041, 5118.714, 5113.915, 5110.231, 
    5104.955,
  5335.867, 5290.922, 5252.775, 5221.983, 5196.178, 5178.462, 5153.085, 
    5145.358, 5130.56, 5120.876, 5114.761, 5109.921, 5105.522, 5102.44, 
    5100.016,
  5330.586, 5286.118, 5248.472, 5216.288, 5190.824, 5164.44, 5151.473, 
    5126.193, 5117.354, 5109.372, 5101.946, 5097.441, 5094.626, 5092.89, 
    5092.376,
  5324.37, 5281.053, 5244.833, 5212.242, 5186.263, 5160.877, 5134.82, 
    5122.173, 5104.559, 5090.063, 5085.984, 5080.631, 5080.188, 5079.029, 
    5081.246,
  5315.897, 5273.896, 5237.734, 5205.826, 5176.129, 5147.668, 5124.218, 
    5096.732, 5080.326, 5071.224, 5062.685, 5059.885, 5060.369, 5062.597, 
    5065.991,
  5305.962, 5268.181, 5231.918, 5200.172, 5169.042, 5138.007, 5106.83, 
    5084.539, 5062.867, 5045.475, 5037.058, 5035.072, 5036.708, 5041.773, 
    5047.82,
  5296.243, 5260.55, 5223.987, 5191.671, 5156.285, 5122.608, 5089.923, 
    5058.49, 5032.781, 5017.063, 5006.793, 5005.146, 5008.857, 5017.75, 
    5026.95,
  5287.379, 5254.188, 5219.252, 5185.028, 5148.354, 5110.421, 5071.477, 
    5038.64, 5008.849, 4984.983, 4972.615, 4971.309, 4977.291, 4989.509, 
    5003.872,
  5280.087, 5246.576, 5211.701, 5175.89, 5134.608, 5093.316, 5052.301, 
    5012.033, 4977.144, 4949.859, 4935.338, 4933.289, 4942.138, 4957.705, 
    4977.603,
  5202.927, 5172.902, 5148.093, 5125.718, 5106.002, 5086.863, 5067.766, 
    5055.583, 5045.229, 5036.445, 5035.917, 5039.318, 5044.461, 5050.906, 
    5058.783,
  5199.43, 5167.589, 5141.252, 5115.884, 5093.721, 5069.117, 5055.844, 
    5033.97, 5023.114, 5018.856, 5015.918, 5019.65, 5026.76, 5037.024, 5045.65,
  5197.337, 5164.175, 5135.647, 5108.369, 5081.445, 5063.833, 5033.725, 
    5025.827, 5007.774, 4996.934, 4993.685, 4997.042, 5005.759, 5017.705, 
    5030.826,
  5193.908, 5158.239, 5127.659, 5096.083, 5069.175, 5040.213, 5026.844, 
    4996.127, 4985.3, 4976.105, 4969.247, 4970.949, 4981.278, 4998.142, 
    5014.779,
  5190.73, 5152.954, 5120.029, 5086.179, 5057.736, 5032.326, 5003.947, 
    4989.667, 4968.361, 4948.329, 4943, 4941.4, 4953.856, 4973.039, 4997.186,
  5186.472, 5144.941, 5108.46, 5074.484, 5043.72, 5016.14, 4993.014, 
    4963.271, 4941.514, 4926.708, 4913.266, 4911.727, 4923.114, 4947.816, 
    4977.402,
  5181.467, 5138.36, 5099.837, 5064.92, 5034.607, 5005.943, 4976.865, 
    4952.982, 4927.162, 4901.743, 4885.778, 4882.82, 4893.027, 4921.828, 
    4957.126,
  5176.062, 5129.571, 5088.729, 5052.987, 5021.127, 4992.244, 4963.111, 
    4931.183, 4901.75, 4878.359, 4858.022, 4852.584, 4864.289, 4896.674, 
    4939.853,
  5170.865, 5123.688, 5082.616, 5045.849, 5014.852, 4983.271, 4949.374, 
    4918.569, 4886.52, 4856.056, 4833.019, 4826.607, 4839.456, 4875.42, 
    4926.011,
  5166.289, 5114.786, 5072.674, 5036.839, 5004.239, 4971.406, 4937.068, 
    4900.193, 4866.146, 4836.368, 4813.378, 4805.776, 4819.846, 4861.353, 
    4915.841,
  5129.912, 5081.58, 5046.263, 5017.958, 4999.131, 4984.742, 4974.133, 
    4970.429, 4969.601, 4974.578, 4986.448, 5002.956, 5022.52, 5039.679, 
    5056.934,
  5110.282, 5061.994, 5029.177, 5001.833, 4983.5, 4967.636, 4962.08, 4953.15, 
    4954.979, 4960.926, 4971.53, 4987.814, 5007.175, 5030.132, 5048.314,
  5092.129, 5045.856, 5014.509, 4987.619, 4968.841, 4958.701, 4944.557, 
    4945.875, 4942.053, 4947.614, 4958.953, 4973.431, 4993.651, 5014.766, 
    5037.553,
  5073.209, 5029.597, 4997.818, 4970.533, 4953.336, 4938.37, 4937.766, 
    4926.616, 4932.506, 4935.452, 4946.51, 4960.923, 4979.824, 5003.964, 
    5028.368,
  5056.658, 5013.899, 4981.034, 4953.635, 4936.184, 4926.586, 4918.268, 
    4919.729, 4918.176, 4923.805, 4934.386, 4948.302, 4967.494, 4989.475, 
    5017.201,
  5040.956, 4996.917, 4960.125, 4932.739, 4913.864, 4904.856, 4903.183, 
    4900.316, 4904.219, 4911.896, 4920.644, 4936.156, 4954.668, 4978.533, 
    5006.235,
  5027.541, 4983.868, 4943.199, 4913.804, 4893.084, 4884.235, 4880.632, 
    4884.961, 4888.866, 4896.192, 4908.06, 4923.653, 4942.77, 4966.669, 
    4995.342,
  5019.359, 4972.502, 4927.243, 4894.616, 4869.401, 4858.693, 4857.272, 
    4861.332, 4869.268, 4881.471, 4894.25, 4911.294, 4932.097, 4957.25, 
    4988.12,
  5017.054, 4968.937, 4920.173, 4882.457, 4853.884, 4838.897, 4835.284, 
    4843.292, 4853.415, 4866.009, 4881.769, 4900.77, 4922.996, 4949.713, 
    4982.377,
  5021.017, 4968.335, 4916.034, 4876.138, 4842.033, 4824.097, 4819.845, 
    4826.508, 4839.59, 4855.567, 4873.048, 4893.366, 4917.388, 4946.759, 
    4982.876,
  5032.557, 4993.119, 4960.844, 4937.852, 4925.505, 4923.08, 4928.734, 
    4940.915, 4952.162, 4960.052, 4970.882, 4990.277, 5017.595, 5049.138, 
    5078.564,
  5006.956, 4962.175, 4928.576, 4903.645, 4895.022, 4897.754, 4911.79, 
    4923.292, 4936.193, 4948.713, 4961.648, 4983.733, 5013.061, 5048.712, 
    5076.984,
  4986.545, 4937.644, 4902.021, 4876.931, 4874.672, 4884.337, 4895.805, 
    4917.97, 4931.116, 4941.726, 4955.375, 4978.978, 5012.095, 5045.42, 
    5075.178,
  4968.704, 4917.179, 4879.131, 4853.846, 4853.856, 4863.371, 4891.594, 
    4905.548, 4923.703, 4936.208, 4951.92, 4977.703, 5013.774, 5049.056, 
    5077.544,
  4958.499, 4905.621, 4865.169, 4838.864, 4837.518, 4855.117, 4879.485, 
    4910.126, 4925.081, 4934.735, 4951.125, 4980.276, 5017.679, 5050.094, 
    5079.612,
  4957.289, 4903.104, 4861.69, 4834.849, 4831.314, 4846.805, 4884.112, 
    4905.67, 4921.381, 4936.261, 4954.336, 4986.543, 5023.235, 5056.105, 
    5084.138,
  4964.77, 4913.489, 4873.495, 4847.576, 4841.441, 4858.72, 4887.079, 
    4914.935, 4928.512, 4940.847, 4961.622, 4994.707, 5029.835, 5060.774, 
    5088.789,
  4981.802, 4931.583, 4893.498, 4870.69, 4863.322, 4878.312, 4901.406, 
    4916.295, 4929.793, 4948.062, 4971.498, 5004.281, 5037.623, 5068.531, 
    5095.921,
  5003.653, 4955.216, 4919.349, 4896.896, 4890.837, 4898.58, 4913.103, 
    4929.057, 4943.163, 4959.348, 4983.307, 5014.81, 5045.428, 5075.634, 
    5102.461,
  5032.119, 4981.296, 4944.955, 4924.303, 4914.127, 4917.997, 4928.17, 
    4938.098, 4951.797, 4971.124, 4996.173, 5025.626, 5054.931, 5084.299, 
    5110.851,
  5039.333, 4992.756, 4951.955, 4919.501, 4892.571, 4869.741, 4855.527, 
    4867.909, 4907.269, 4947.762, 4980.851, 5010.924, 5034.936, 5057.592, 
    5082.934,
  5032.187, 4987.288, 4949.385, 4920.095, 4896.537, 4870.911, 4861.036, 
    4871.649, 4910.608, 4951.53, 4982.82, 5009.11, 5029.899, 5053.544, 
    5078.488,
  5031.163, 4989.551, 4955.218, 4931.156, 4908.859, 4896.232, 4881.2, 
    4893.02, 4930.052, 4960.751, 4986.383, 5007.271, 5027.347, 5047.739, 
    5075.448,
  5033.281, 4994.456, 4964.431, 4941.436, 4928.507, 4910.196, 4912.937, 
    4918.703, 4944.434, 4969.019, 4990.903, 5006.427, 5026.32, 5049.201, 
    5078.46,
  5038.856, 5003.524, 4976.579, 4956.384, 4945.322, 4938.574, 4936.069, 
    4942.8, 4965.297, 4975.89, 4993.928, 5007.197, 5028.811, 5051.982, 
    5083.729,
  5046.033, 5013.057, 4988.063, 4970.455, 4959.613, 4952.801, 4954.47, 
    4960.437, 4966.897, 4983.839, 4996.048, 5012.848, 5035.414, 5062.99, 
    5093.405,
  5054.112, 5024.065, 5001.227, 4984.109, 4973.001, 4968.247, 4965.178, 
    4970.694, 4980.614, 4990.288, 5002.9, 5023.607, 5047.483, 5075.887, 
    5106.616,
  5063.396, 5033.52, 5010.836, 4995.279, 4982.274, 4975.296, 4974.391, 
    4977.073, 4983.744, 4998.71, 5016.912, 5040.023, 5065.296, 5093.841, 
    5124.308,
  5073.927, 5044.733, 5021.91, 5006.011, 4995.237, 4989.144, 4986.396, 
    4992.315, 5003.772, 5018.375, 5038.003, 5061.27, 5085.089, 5113.271, 
    5141.548,
  5087.569, 5055.76, 5032.059, 5017.645, 5007.005, 5002.94, 5004.639, 
    5010.846, 5022.666, 5041.056, 5061.808, 5083.584, 5106.86, 5132.647, 
    5159.285,
  5106.44, 5080.213, 5057.04, 5037.677, 5019.111, 5000.201, 4977.594, 
    4963.324, 4952.836, 4955.694, 4965.642, 4976.135, 4991.439, 5004.748, 
    5022.677,
  5097.475, 5073.111, 5053.274, 5039.106, 5027.562, 5012.54, 5004.883, 
    4994.104, 4988.175, 4994.422, 5002.874, 5015.41, 5024.82, 5038.811, 
    5053.903,
  5093.806, 5070.77, 5054.699, 5046.132, 5036.524, 5038.007, 5025.872, 
    5026.414, 5029.082, 5031.677, 5037.612, 5046.035, 5057.296, 5067.501, 
    5079.277,
  5093.34, 5070.455, 5057.888, 5048.834, 5050.074, 5042.417, 5052.695, 
    5050.274, 5051.321, 5057.945, 5066.061, 5071.827, 5079.986, 5088.75, 
    5100.056,
  5096.427, 5075.035, 5062.807, 5056.52, 5058.78, 5062.982, 5065.932, 
    5068.82, 5078.408, 5077.996, 5085.024, 5088.664, 5097.227, 5101.399, 
    5111.218,
  5104.219, 5083.402, 5067.931, 5062.283, 5063.402, 5066.468, 5074.822, 
    5078.92, 5081.151, 5089.202, 5092.917, 5097.374, 5103.081, 5109.664, 
    5117.534,
  5116.222, 5096.927, 5080.305, 5071.054, 5069.212, 5074.021, 5076.996, 
    5084.409, 5089.206, 5089.978, 5092.377, 5098.139, 5104.212, 5111.233, 
    5120.185,
  5131.876, 5112.773, 5095.38, 5083.684, 5075.068, 5073.479, 5076.077, 
    5078.164, 5078.157, 5081.011, 5085.217, 5092.594, 5102.297, 5113.048, 
    5125.362,
  5150.343, 5131.388, 5114.893, 5102.211, 5092.196, 5084.712, 5078.378, 
    5076.858, 5075.258, 5075.034, 5079.225, 5090.56, 5103.522, 5117.806, 
    5135.303,
  5170.923, 5148.567, 5133.421, 5121.802, 5109.64, 5100.389, 5092.881, 
    5084.875, 5079.759, 5080.259, 5086.822, 5098.815, 5114.509, 5134, 5155.432,
  5220.375, 5205.972, 5196.5, 5185.473, 5173.897, 5160.727, 5142.17, 5125.2, 
    5101.208, 5067.478, 5029.519, 4984.564, 4941.575, 4913.162, 4911.73,
  5228.468, 5210.33, 5198.65, 5185.315, 5173.568, 5157.153, 5147.191, 
    5124.822, 5106.449, 5083.542, 5050.164, 5012.755, 4971.25, 4941.52, 
    4929.261,
  5237.888, 5216.486, 5201.08, 5187.2, 5171.006, 5160.654, 5140.217, 
    5133.556, 5117.06, 5097.951, 5073.385, 5042.05, 5007.96, 4975.935, 
    4957.738,
  5247.719, 5223.098, 5203.192, 5185.772, 5169.777, 5152.413, 5143.492, 
    5125.408, 5118.286, 5108.778, 5091.973, 5068.897, 5043.998, 5018.46, 
    4999.535,
  5258.359, 5231.98, 5208.232, 5187.487, 5169.46, 5152.507, 5135.341, 
    5125.202, 5117.622, 5114.081, 5106.702, 5090.527, 5074.483, 5056.52, 
    5043.956,
  5268.209, 5240.977, 5214.131, 5189.853, 5167.645, 5148.169, 5131.678, 
    5114.222, 5108.732, 5113.891, 5113.695, 5107.258, 5097.383, 5087.491, 
    5079.459,
  5277.232, 5250.534, 5222.589, 5196.306, 5171.031, 5148.32, 5127.22, 
    5110.958, 5103.547, 5108.596, 5115.161, 5117.057, 5114.584, 5111.64, 
    5108.574,
  5285.84, 5257.492, 5229.872, 5202.675, 5174.738, 5150.146, 5127.878, 
    5106.171, 5094.525, 5100.687, 5111.705, 5120.322, 5124.726, 5127.808, 
    5130.292,
  5292.484, 5265.488, 5238.696, 5210.099, 5182.685, 5157.741, 5134.408, 
    5113.352, 5099.218, 5098.143, 5108.673, 5121.562, 5130.785, 5137.735, 
    5144.303,
  5299.965, 5271.871, 5243.742, 5216.113, 5188.566, 5164.863, 5144.587, 
    5124.182, 5109.857, 5107.241, 5115.1, 5126.406, 5135.78, 5144.765, 5153.93,
  5355.981, 5326.38, 5297.473, 5263.915, 5232.907, 5200.637, 5169.739, 
    5141.989, 5124.05, 5100.173, 5067.523, 5021.561, 4976.563, 4944.202, 
    4928.658,
  5351.06, 5321.69, 5292.868, 5259.036, 5228.493, 5191.595, 5172.68, 
    5137.495, 5124.239, 5107.69, 5077.199, 5038.033, 4994.041, 4965.452, 
    4948.879,
  5347.191, 5318.854, 5289.676, 5257.885, 5223.585, 5197.738, 5160.024, 
    5144.338, 5128.746, 5116.83, 5090.916, 5058.259, 5019.946, 4987.533, 
    4968.266,
  5342.936, 5314.542, 5285.886, 5253.06, 5220.972, 5186.705, 5166.863, 
    5139.151, 5133.017, 5124.634, 5106.779, 5080.872, 5049.688, 5020.094, 
    4995.177,
  5339.449, 5311.549, 5283.96, 5250.799, 5219.117, 5186.771, 5160.135, 
    5141.645, 5138.381, 5132.694, 5121.024, 5100.812, 5077.285, 5050.764, 
    5028.369,
  5335.788, 5308.359, 5279.568, 5248.461, 5214.736, 5182.046, 5161.892, 
    5140.82, 5138.752, 5139.254, 5132.06, 5118.944, 5099.515, 5078.279, 
    5056.693,
  5332.925, 5306.339, 5278.255, 5247.893, 5213.245, 5181.882, 5160.951, 
    5143.83, 5141.7, 5144.32, 5140.547, 5132.626, 5117.74, 5100.635, 5080.706,
  5330.973, 5303.351, 5276.035, 5245.604, 5209.553, 5180.213, 5162.81, 
    5144.197, 5141.072, 5147.075, 5146.356, 5141.555, 5130.492, 5117.83, 
    5101.494,
  5328.84, 5302.345, 5276.231, 5245.389, 5211.373, 5181.749, 5164.894, 
    5148.553, 5142.658, 5148.126, 5148.575, 5145.812, 5138.058, 5128.428, 
    5116.231,
  5327.512, 5299.734, 5274.324, 5244.892, 5210.313, 5181.941, 5168.139, 
    5152.041, 5143.677, 5147.205, 5149.052, 5146.71, 5141.245, 5134.668, 
    5125.716,
  5363.641, 5339.406, 5317.307, 5293.528, 5271.25, 5242.751, 5212.103, 
    5189.458, 5172.267, 5161.963, 5153.77, 5139.383, 5118.431, 5091.135, 
    5067.996,
  5356.197, 5330.413, 5307.174, 5282.782, 5259.038, 5223.611, 5199.417, 
    5174.083, 5160.559, 5157.359, 5150.334, 5139.425, 5119.973, 5099.142, 
    5073.688,
  5351.137, 5325.09, 5300.742, 5276.394, 5248.268, 5220.945, 5182.394, 
    5172.104, 5155.412, 5151.914, 5146.519, 5137.93, 5120.707, 5100.441, 
    5079.272,
  5347.38, 5320.208, 5295.381, 5267.909, 5240.723, 5200.834, 5183.671, 
    5157.288, 5149.217, 5146.429, 5143.004, 5135.332, 5119.805, 5102.641, 
    5083.263,
  5345.27, 5318.164, 5292.833, 5263.992, 5235.181, 5199.702, 5173.156, 
    5159.643, 5144.718, 5141.454, 5138.934, 5131.396, 5116.456, 5099.837, 
    5083.715,
  5343.809, 5316.353, 5289.373, 5260.158, 5229.612, 5193.378, 5173.421, 
    5152.759, 5139.773, 5138.712, 5134.661, 5127.045, 5111.92, 5097.597, 
    5082.847,
  5343.054, 5316.787, 5289.683, 5258.854, 5229.535, 5193.789, 5172.671, 
    5155.662, 5141.375, 5136.265, 5131.005, 5121.772, 5106.627, 5093.005, 
    5077.709,
  5343.332, 5316.447, 5288.616, 5257.005, 5227.205, 5193.193, 5174.304, 
    5155.065, 5140.31, 5135.878, 5128.638, 5117.875, 5102.787, 5088.603, 
    5071.946,
  5343.697, 5318.057, 5290.663, 5257.772, 5229.804, 5196.5, 5177.265, 
    5160.671, 5145.506, 5137.643, 5127.701, 5115.898, 5099.641, 5082.197, 
    5061.629,
  5344.814, 5317.875, 5290.17, 5257.424, 5229.798, 5198.261, 5180.821, 
    5164.518, 5148.809, 5140.771, 5129.409, 5116.726, 5098.496, 5077.496, 
    5053.343,
  5373.774, 5347.798, 5319.373, 5286.067, 5256.653, 5227.247, 5198.209, 
    5178.599, 5159.162, 5140.243, 5127.388, 5120.497, 5117.604, 5116.428, 
    5115.388,
  5374.928, 5347.784, 5317.612, 5282.135, 5250.947, 5216.196, 5194.536, 
    5167.038, 5147.209, 5133.685, 5120.252, 5113.44, 5108.698, 5106.944, 
    5102.167,
  5375.737, 5348.472, 5317.043, 5281.729, 5246.582, 5220.038, 5183.438, 
    5170.616, 5146.559, 5128.886, 5114.224, 5107.233, 5099.391, 5094.106, 
    5086.706,
  5375.724, 5347.312, 5316.019, 5278.25, 5244.349, 5208.186, 5188.14, 
    5158.401, 5138.584, 5125.053, 5108.918, 5098.274, 5087.177, 5078.224, 
    5068.836,
  5375.142, 5346.871, 5316.385, 5278.007, 5243.201, 5210.59, 5180.275, 
    5163.466, 5141.007, 5118.296, 5102.374, 5085.583, 5071.463, 5058.58, 
    5049.583,
  5373.578, 5345.242, 5314.3, 5276.672, 5240.181, 5207.933, 5181.826, 
    5155.483, 5131.501, 5114.066, 5092.643, 5072.959, 5054.947, 5040.93, 
    5030.864,
  5371.219, 5344.098, 5314.065, 5276.778, 5241.474, 5209.941, 5181.309, 
    5160.199, 5134.989, 5110.107, 5085.802, 5064.124, 5043.215, 5029.715, 
    5019.203,
  5368.357, 5341.585, 5311.465, 5275.253, 5239.859, 5210.145, 5182.907, 
    5158.085, 5131.49, 5109.697, 5084.36, 5060.333, 5039.044, 5025.993, 
    5018.252,
  5364.515, 5339.929, 5311.114, 5275.964, 5242.768, 5213.641, 5185.98, 
    5163.625, 5138.004, 5113.66, 5087.306, 5063.268, 5041.963, 5029.82, 
    5022.542,
  5360.647, 5336.086, 5307.406, 5274.316, 5242.432, 5215.363, 5189.559, 
    5165.789, 5140.989, 5119.714, 5095.717, 5072.855, 5052.992, 5042.352, 
    5036.199,
  5404.487, 5382.597, 5357.474, 5327.497, 5293.623, 5259.089, 5225.065, 
    5200.962, 5179.593, 5155.401, 5136.762, 5121.581, 5110.751, 5102.846, 
    5101.42,
  5396.3, 5374.178, 5348.963, 5317.473, 5283.208, 5245.351, 5221.877, 
    5191.798, 5168.791, 5150.2, 5129.988, 5112.227, 5097.538, 5089.253, 
    5084.752,
  5388.841, 5367.954, 5341.716, 5311.237, 5274.404, 5249.124, 5209.548, 
    5196.627, 5172.724, 5147.845, 5124.246, 5104.447, 5085.345, 5073.434, 
    5068.063,
  5382.249, 5361.107, 5335.596, 5302.391, 5268.731, 5233.801, 5216.061, 
    5188.604, 5167.262, 5148.714, 5122.749, 5099.007, 5076.844, 5060.003, 
    5051.571,
  5377.543, 5356.475, 5331.942, 5298.346, 5266.381, 5236.491, 5210.101, 
    5194.284, 5177.341, 5149.238, 5126.043, 5097.212, 5072.861, 5049.664, 
    5038.506,
  5373.902, 5353.319, 5328.111, 5296.289, 5263.11, 5233.416, 5212.835, 
    5193.09, 5174.975, 5155.348, 5130.302, 5100.822, 5072.609, 5046.173, 
    5029.754,
  5371.232, 5352.409, 5327.779, 5297.729, 5267.131, 5238.29, 5213.77, 
    5200.189, 5184.716, 5162.491, 5136.357, 5106.65, 5074.503, 5044.758, 
    5023.597,
  5369.253, 5351.676, 5327.761, 5299.971, 5269.535, 5241.55, 5218.397, 
    5200.848, 5185.237, 5168.247, 5143.863, 5113.791, 5080.045, 5046.208, 
    5020.267,
  5367.597, 5351.61, 5329.907, 5304.834, 5277.907, 5250.179, 5224.505, 
    5207.81, 5193.474, 5174.235, 5150.279, 5121.626, 5087.385, 5050.532, 
    5020.109,
  5365.765, 5350.112, 5331.085, 5308.881, 5282.602, 5256.345, 5231.657, 
    5210.409, 5194.649, 5177.869, 5156.391, 5130.035, 5096.881, 5058.643, 
    5023.718,
  5445.806, 5422.126, 5396.785, 5368.527, 5342.764, 5322.634, 5307.936, 
    5297.342, 5281.997, 5258.688, 5236.381, 5212.519, 5193.63, 5177.657, 
    5166.429,
  5448.025, 5424.377, 5398.851, 5371.346, 5345.724, 5322.916, 5312.894, 
    5294.888, 5278.69, 5260.435, 5237.131, 5212.401, 5191.189, 5175.07, 
    5159.895,
  5449.66, 5426.621, 5401.414, 5375.802, 5348.592, 5331.743, 5309.744, 
    5302.104, 5283.02, 5259.24, 5235.951, 5211.654, 5188.338, 5170.162, 
    5151.695,
  5449.199, 5426.385, 5401.989, 5376.291, 5351.566, 5327.711, 5315.232, 
    5293.324, 5276.27, 5257.808, 5232.538, 5208.224, 5184.971, 5165.207, 
    5143.096,
  5446.818, 5424.795, 5401.688, 5376.822, 5353.412, 5331.739, 5310.874, 
    5297.705, 5278.978, 5251.956, 5229.903, 5202.194, 5180.199, 5156.828, 
    5133.613,
  5441.596, 5419.664, 5396.597, 5373.828, 5350.773, 5329.286, 5311.026, 
    5288.648, 5268.562, 5246.929, 5223.091, 5195.914, 5173.376, 5148.771, 
    5122.965,
  5433.661, 5413.506, 5390.501, 5368.54, 5347.74, 5327.892, 5307.917, 
    5290.139, 5268.727, 5242.343, 5216.373, 5189.174, 5164.661, 5139.194, 
    5110.096,
  5424.613, 5403.864, 5380.314, 5360.18, 5339.982, 5322.056, 5303.795, 
    5282.618, 5260.204, 5236.052, 5209.438, 5181.192, 5156.219, 5129.187, 
    5098.646,
  5414.797, 5394.138, 5371.183, 5350.829, 5332.786, 5315.598, 5297.3, 
    5278.443, 5256.159, 5229.698, 5202.026, 5172.73, 5146.716, 5118.497, 
    5086.958,
  5405.125, 5381.934, 5358.899, 5340.669, 5322.542, 5305.29, 5287.549, 
    5266.014, 5243.952, 5219.754, 5193.139, 5163.577, 5137.5, 5108.717, 
    5076.762,
  5533.108, 5509.543, 5486.41, 5460.799, 5437.783, 5414.406, 5391.234, 
    5373.114, 5355.959, 5336.781, 5322.623, 5308.337, 5295.289, 5282.988, 
    5274.46,
  5522.261, 5499.324, 5477.164, 5452.445, 5429.372, 5403.064, 5387.121, 
    5361.613, 5346.23, 5334.903, 5320.477, 5307.251, 5294.648, 5283.951, 
    5274.146,
  5509.405, 5488.252, 5466.049, 5444.119, 5418.833, 5401.515, 5371.242, 
    5363.454, 5342.932, 5327.524, 5314.505, 5302.768, 5289.45, 5278.585, 
    5268.074,
  5493.628, 5473.836, 5453.085, 5430.974, 5408.884, 5383.174, 5369.599, 
    5341.723, 5330.43, 5319.109, 5304.158, 5292.087, 5279.74, 5268.559, 
    5257.519,
  5477.814, 5459.622, 5440.133, 5419.351, 5397.669, 5376.041, 5351.896, 
    5340.722, 5321.051, 5302.432, 5290.235, 5274.426, 5263.209, 5250.227, 
    5241.17,
  5461.466, 5445.003, 5425.562, 5405.895, 5382.151, 5359.866, 5339.812, 
    5316.731, 5298.946, 5283.477, 5265.422, 5249.542, 5236.771, 5224.911, 
    5216.151,
  5446.859, 5432.112, 5412.886, 5392.383, 5369.539, 5345.843, 5322.195, 
    5301.774, 5277.974, 5253.22, 5233.22, 5215.023, 5200.284, 5189.81, 
    5182.293,
  5434.366, 5418.637, 5398.574, 5377.44, 5351.504, 5326.723, 5300.021, 
    5270.578, 5241.793, 5216.505, 5191.919, 5171.762, 5157.211, 5148.158, 
    5143.29,
  5422.805, 5408.07, 5387.586, 5363.648, 5336.306, 5306.343, 5272.362, 
    5240.127, 5207.214, 5175.172, 5149.828, 5130.041, 5116.715, 5109.203, 
    5106.344,
  5414.371, 5397.32, 5374.095, 5347.649, 5314.347, 5278.137, 5239.797, 
    5200.8, 5166.568, 5136.615, 5113.193, 5096.193, 5085.745, 5080.071, 
    5077.89,
  5454.753, 5435.97, 5421.438, 5406.688, 5394.879, 5380.817, 5363.196, 
    5348.423, 5331.439, 5313.116, 5301.019, 5291.369, 5284.423, 5277.903, 
    5274.465,
  5439.324, 5424.114, 5411.787, 5398.317, 5386.243, 5367.133, 5353.85, 
    5327.283, 5309.495, 5296.864, 5283.466, 5275.727, 5269.936, 5268.251, 
    5265.534,
  5429.352, 5418.119, 5405.938, 5394.274, 5376.937, 5362.631, 5330.27, 
    5317.107, 5290.174, 5272.216, 5259.765, 5252.95, 5247.636, 5247.113, 
    5247.831,
  5424.149, 5413.033, 5401.609, 5386.071, 5367.006, 5340.221, 5320.819, 
    5279.657, 5260.921, 5244.884, 5231.288, 5222.767, 5219.125, 5218.381, 
    5221.434,
  5421.729, 5411.588, 5399.034, 5380.25, 5357.089, 5328.389, 5289.833, 
    5266.771, 5238.788, 5214.255, 5202.98, 5189.937, 5185.145, 5180.778, 
    5185.278,
  5421.825, 5409.795, 5393.889, 5371.527, 5342.842, 5307.901, 5269.423, 
    5230.479, 5205.506, 5190.171, 5172.588, 5160.03, 5151.563, 5145.821, 
    5146.098,
  5422.593, 5408.792, 5390.35, 5363.614, 5332.379, 5290.419, 5244.953, 
    5215.989, 5189.415, 5166.886, 5149.91, 5136.773, 5125.076, 5117.622, 
    5113.519,
  5423.165, 5406.104, 5384.516, 5353.501, 5317.297, 5271.315, 5225.841, 
    5194.729, 5169.066, 5151.928, 5133.266, 5118.586, 5105.568, 5095.798, 
    5088.451,
  5423.218, 5404.848, 5380.368, 5345.808, 5307.839, 5257.748, 5213.751, 
    5189.208, 5162.941, 5140.727, 5119.825, 5103.762, 5088.529, 5077.128, 
    5067.26,
  5423.43, 5400.74, 5373.079, 5337.148, 5295.213, 5245.057, 5206.809, 
    5179.602, 5152.195, 5129.847, 5107.229, 5089.192, 5073.385, 5061.73, 
    5051.344,
  5441.712, 5415.572, 5388.348, 5358.289, 5327.541, 5293.655, 5258.684, 
    5232.291, 5205.948, 5180.793, 5166.658, 5160.173, 5160.018, 5165.544, 
    5175.458,
  5448.057, 5420.855, 5391.331, 5358.988, 5326.385, 5284.986, 5256.168, 
    5217.609, 5189.177, 5169.947, 5154.354, 5146.551, 5145.057, 5150.836, 
    5159.911,
  5454.002, 5426.624, 5395.181, 5363.186, 5325.505, 5293.948, 5244.462, 
    5223.845, 5191.525, 5164.482, 5145.601, 5136.642, 5132.177, 5136.122, 
    5144.572,
  5458.045, 5429.734, 5398.099, 5362.974, 5327.537, 5283.724, 5253.05, 
    5211.156, 5181.674, 5161.05, 5140.622, 5129.066, 5123.619, 5124.969, 
    5131.398,
  5461.407, 5433.079, 5401.673, 5365.692, 5330.126, 5290.1, 5247.433, 
    5220.577, 5190.588, 5157.005, 5137.746, 5121.708, 5115.736, 5114.162, 
    5119.652,
  5463.206, 5434.68, 5402.027, 5367.653, 5330.095, 5290.265, 5252.574, 
    5215.194, 5181.631, 5157.625, 5134.191, 5116.824, 5107.732, 5105.021, 
    5109.518,
  5463.597, 5436.685, 5404.099, 5369.852, 5333.774, 5294.595, 5254.058, 
    5223.08, 5189.955, 5158.496, 5132.525, 5113.175, 5099.749, 5095.336, 
    5097.712,
  5463.034, 5435.891, 5402.924, 5370.038, 5333.066, 5295.621, 5257.078, 
    5221.725, 5187.062, 5159.203, 5132.769, 5110.879, 5094.424, 5086.689, 
    5085.88,
  5461.241, 5435.769, 5403.813, 5370.674, 5335.479, 5297.903, 5258.89, 
    5226.609, 5193.512, 5161.897, 5133.486, 5109.627, 5090.336, 5079.222, 
    5075.079,
  5458.592, 5431.468, 5400.115, 5368.886, 5333.016, 5296.278, 5259.033, 
    5224.341, 5191.627, 5162.297, 5134.508, 5109.107, 5087.686, 5073.785, 
    5066.352,
  5497.081, 5467.053, 5437.551, 5406.764, 5376.479, 5345.138, 5309.008, 
    5279.282, 5247.766, 5213.065, 5186.432, 5166.417, 5154.583, 5151.333, 
    5157.686,
  5497.796, 5467.668, 5438.365, 5407.887, 5378.425, 5343.099, 5316.968, 
    5274.439, 5243.067, 5215.883, 5188.024, 5166.062, 5151.423, 5145.405, 
    5148.134,
  5496.625, 5466.989, 5437.459, 5408.748, 5376.423, 5351.776, 5307.612, 
    5288.136, 5249.881, 5216.308, 5187.472, 5164.955, 5147.426, 5138.934, 
    5138.203,
  5492.412, 5462.574, 5433.603, 5403.677, 5374.612, 5339.49, 5314.502, 
    5268.302, 5239.113, 5212.274, 5184.365, 5161.322, 5143.495, 5132.361, 
    5129.661,
  5486.446, 5457.139, 5428.576, 5399.283, 5369.669, 5338.358, 5301.606, 
    5275.235, 5239.801, 5202.627, 5179.661, 5155.456, 5138.695, 5124.404, 
    5120.806,
  5477.549, 5448.318, 5419.421, 5390.999, 5359.686, 5327.916, 5294.747, 
    5254.676, 5219.397, 5193.71, 5169.655, 5149.693, 5132.147, 5118.04, 
    5111.576,
  5466.372, 5438.9, 5410.296, 5381.027, 5350.098, 5315.905, 5279.101, 
    5245.918, 5211.144, 5182.029, 5159.543, 5142.209, 5124.506, 5111.094, 
    5101.865,
  5453.654, 5426.95, 5397.414, 5368.276, 5334.353, 5299.119, 5261.549, 
    5222.437, 5190.34, 5168.578, 5149.486, 5133.522, 5117, 5103.02, 5092.468,
  5440.26, 5415.417, 5386.564, 5355.3, 5320.022, 5282.264, 5242.415, 
    5208.138, 5180.655, 5158.126, 5140.063, 5124.75, 5108.235, 5094.136, 
    5083.774,
  5427.41, 5401.351, 5370.745, 5339.012, 5300.46, 5262.434, 5223.68, 
    5189.326, 5165.016, 5147.321, 5131.502, 5115.864, 5099.556, 5085.789, 
    5076.408,
  5429.18, 5409.384, 5386.724, 5360.991, 5336.649, 5313.485, 5288.626, 
    5270.586, 5250.89, 5228.266, 5209.423, 5194.103, 5182.182, 5174.137, 
    5171.302,
  5414.376, 5392.031, 5367.962, 5342.023, 5316.785, 5290.467, 5271.303, 
    5242.339, 5220.357, 5204.37, 5184.36, 5170.957, 5161.72, 5159.973, 
    5158.116,
  5398.296, 5375.448, 5350.233, 5324.812, 5296.026, 5277.897, 5241.865, 
    5230.353, 5199.107, 5174.218, 5155.268, 5144.125, 5139.108, 5141.178, 
    5144.816,
  5382.224, 5358.917, 5333.448, 5305.119, 5278.043, 5246.715, 5229.227, 
    5187.526, 5163.744, 5142.488, 5123.99, 5116.889, 5117.894, 5124.219, 
    5131.76,
  5368.556, 5345.34, 5318.618, 5288.239, 5257.901, 5231.074, 5194.698, 
    5176.616, 5145.127, 5112.849, 5101.649, 5096.211, 5101.804, 5109.838, 
    5120.156,
  5357.649, 5331.93, 5302.359, 5270.754, 5239.509, 5207.636, 5177.713, 
    5140.877, 5114.354, 5099.275, 5087.619, 5086.269, 5091.957, 5100.281, 
    5109.839,
  5347.23, 5320.978, 5289.095, 5256.35, 5223.228, 5191.924, 5158.717, 
    5135.796, 5113.65, 5093.644, 5083.598, 5082.327, 5085.32, 5092.304, 
    5099.961,
  5338.495, 5309.921, 5275.826, 5241.69, 5208.782, 5177.803, 5149.188, 
    5122.393, 5102.396, 5091.382, 5083.542, 5080.465, 5081.009, 5084.821, 
    5090.191,
  5331.311, 5301.623, 5265.716, 5231.137, 5198.627, 5169.849, 5144.04, 
    5125.702, 5108.879, 5093.456, 5082.988, 5077.439, 5074.797, 5075.643, 
    5078.88,
  5325.729, 5291.963, 5254.729, 5220.615, 5190.469, 5164.463, 5143.231, 
    5122.375, 5106.187, 5093.107, 5082.414, 5073.637, 5068.167, 5066.293, 
    5067.562,
  5285.19, 5257.106, 5231.075, 5203.16, 5175.385, 5149.103, 5123.287, 
    5106.149, 5093.216, 5083.774, 5084.299, 5095.126, 5112.88, 5132.834, 
    5153.121,
  5276.226, 5246.082, 5218.157, 5187.328, 5158.242, 5126.354, 5107.915, 
    5083.051, 5068.018, 5061.388, 5060.538, 5070.104, 5089.032, 5113.19, 
    5135.896,
  5269.115, 5238.431, 5208.714, 5178.071, 5145.521, 5124.953, 5090.18, 
    5079.12, 5059.517, 5045.502, 5040.386, 5050.426, 5070.26, 5094.406, 
    5121.421,
  5262.188, 5231.241, 5201.78, 5170.04, 5140.964, 5111.569, 5095.356, 
    5066.393, 5049.583, 5038.552, 5030.438, 5038.028, 5056.596, 5081.925, 
    5108.914,
  5258.568, 5228.459, 5199.4, 5168.75, 5142.622, 5117.591, 5091.791, 
    5073.979, 5057.373, 5038.477, 5031.554, 5033.423, 5050.554, 5070.841, 
    5098.974,
  5256.864, 5227.304, 5198.422, 5171.169, 5144.148, 5121.22, 5099.584, 
    5076.031, 5057.04, 5046.969, 5038.248, 5038.246, 5049.806, 5067.969, 
    5091.755,
  5257.911, 5230.199, 5202.14, 5177.035, 5153.523, 5130.957, 5106.758, 
    5088.221, 5070.434, 5054.855, 5046.661, 5046.408, 5052.5, 5067.928, 
    5087.449,
  5260.658, 5234.05, 5207.174, 5184.181, 5159.829, 5138.768, 5116.231, 
    5094.173, 5074.599, 5062.953, 5054.634, 5053.81, 5057.692, 5070.011, 
    5085.365,
  5266.98, 5242.157, 5216.423, 5194.705, 5172.893, 5150.323, 5125.956, 
    5105.603, 5086.042, 5070.01, 5059.761, 5057.646, 5060.581, 5070.09, 
    5083.353,
  5275.584, 5250.19, 5226.585, 5206.307, 5182.141, 5159.562, 5135.694, 
    5111.994, 5090.733, 5074.762, 5063.49, 5059.474, 5060.923, 5069.206, 
    5080.953,
  5274.243, 5238.24, 5205.558, 5172.02, 5142.307, 5115.976, 5090.421, 
    5073.784, 5061.435, 5049.23, 5045.489, 5050.368, 5066.802, 5092.999, 
    5124.096,
  5281.656, 5243.937, 5208.722, 5172.553, 5140.966, 5107.736, 5090.052, 
    5063.647, 5048.918, 5039.694, 5032.141, 5030.311, 5035.286, 5059.608, 
    5089.963,
  5291.651, 5252.483, 5214.24, 5177.255, 5139.992, 5115.043, 5080.561, 
    5067.85, 5050.112, 5037.048, 5026.259, 5019.066, 5018.877, 5031.695, 
    5060.394,
  5301.099, 5260.443, 5220.504, 5179.565, 5142.851, 5106.719, 5088.187, 
    5061.111, 5047.399, 5037.991, 5026.445, 5016.069, 5013.427, 5022.886, 
    5045.493,
  5312.454, 5271.113, 5229.789, 5186.933, 5148.411, 5114.158, 5085.236, 
    5068.378, 5056.401, 5042.619, 5032.213, 5019.373, 5018.076, 5022.763, 
    5044.078,
  5323.406, 5281.722, 5237.806, 5194.754, 5152.663, 5116.601, 5091.537, 
    5070.591, 5058.185, 5052.583, 5043.816, 5035.169, 5031.823, 5038.237, 
    5053.915,
  5335.114, 5294.998, 5250.204, 5206.406, 5163.884, 5125.967, 5095.764, 
    5079.325, 5069.954, 5063.209, 5058.86, 5056.053, 5056.365, 5061.862, 
    5074.41,
  5346.599, 5307.866, 5262.132, 5217.687, 5173.262, 5134.636, 5103.949, 
    5083.187, 5073.375, 5071.98, 5072.572, 5073.953, 5078.286, 5086.201, 
    5097.143,
  5358.921, 5323.307, 5278.529, 5234.207, 5191.064, 5150.004, 5114.61, 
    5092.776, 5082.651, 5079.845, 5081.82, 5086.993, 5093.188, 5102.412, 
    5113.159,
  5370.902, 5337.445, 5295.263, 5251.389, 5206.161, 5165.631, 5130.158, 
    5101.634, 5087.852, 5085.453, 5089.018, 5095.767, 5104.129, 5113.878, 
    5124.828,
  5348.679, 5306.256, 5258.361, 5208.819, 5164.389, 5138.485, 5114.596, 
    5098.539, 5086.397, 5076.581, 5082.741, 5099.737, 5123.761, 5151.623, 
    5178.894,
  5345.92, 5305.146, 5258.047, 5209.241, 5167.885, 5140.078, 5126.151, 
    5102.157, 5086.452, 5078.524, 5078.709, 5091.911, 5113.072, 5142.844, 
    5166.959,
  5344.124, 5306.096, 5259.766, 5213.852, 5172.673, 5155.646, 5130.326, 
    5117.236, 5100.508, 5084.27, 5077.942, 5084.572, 5101.171, 5124.827, 
    5153.159,
  5341.628, 5306.154, 5262.091, 5215.687, 5180.559, 5157.211, 5148.994, 
    5128.893, 5108.337, 5092.746, 5079.885, 5078.374, 5088.961, 5110.506, 
    5135.746,
  5340.482, 5308.291, 5266.012, 5221.425, 5188.813, 5170.539, 5159.088, 
    5142.861, 5132.043, 5107.445, 5090.819, 5076.854, 5078.504, 5090.915, 
    5115.366,
  5339.717, 5310.434, 5268.808, 5227.318, 5193.631, 5176.353, 5173.101, 
    5160.354, 5143.625, 5127.089, 5110.064, 5089.629, 5076.598, 5077.559, 
    5095.051,
  5340.214, 5314.378, 5274.437, 5234.773, 5202.37, 5184.239, 5179.505, 
    5175.22, 5165.787, 5149.186, 5130.293, 5112.703, 5092.916, 5076.983, 
    5078.505,
  5341.532, 5318.469, 5280.505, 5242.262, 5208.263, 5188.142, 5186.434, 
    5185.137, 5177.547, 5167.441, 5152.516, 5134.562, 5116.373, 5098.501, 
    5084.612,
  5344.433, 5324.562, 5289.881, 5252.474, 5220.441, 5196.741, 5189.469, 
    5193.149, 5192.428, 5184.934, 5172.811, 5157.881, 5140.709, 5123.828, 
    5108.133,
  5348.314, 5330.727, 5299.835, 5263.708, 5229.632, 5205.011, 5194.328, 
    5195.787, 5198.203, 5196.341, 5189.396, 5177.529, 5163.822, 5149.352, 
    5135.635,
  5315.725, 5298.936, 5281.152, 5260.623, 5240.042, 5227.013, 5204.231, 
    5179.663, 5153.112, 5138.117, 5147.826, 5160.447, 5172.204, 5179.445, 
    5184.97,
  5302.558, 5286.023, 5270.01, 5250.305, 5235.198, 5227.084, 5212.787, 
    5182.84, 5156.334, 5141.485, 5148.202, 5161.316, 5174.026, 5184.562, 
    5190.752,
  5291.82, 5275.942, 5259.95, 5242.997, 5234.283, 5235.067, 5215.465, 
    5197.638, 5173.843, 5151.412, 5149.268, 5159.698, 5173.789, 5184.935, 
    5193.006,
  5283.586, 5265.094, 5248.23, 5236.128, 5236.966, 5234.198, 5228.092, 
    5207.915, 5184.083, 5165.449, 5150.756, 5157.438, 5170.166, 5185.368, 
    5195.592,
  5278.424, 5257.474, 5243.811, 5236.893, 5242.068, 5242.887, 5234.855, 
    5218.631, 5204.797, 5179.101, 5163.082, 5152.518, 5163.778, 5179.129, 
    5193.389,
  5278.708, 5256.743, 5242.549, 5239.384, 5244.596, 5248.094, 5244.546, 
    5231.093, 5212.101, 5194.696, 5175.874, 5157.01, 5154.6, 5171.34, 5188.324,
  5286.055, 5262.244, 5248.586, 5245.345, 5251.071, 5256.497, 5251.396, 
    5243.395, 5229.662, 5210.248, 5189.576, 5170.724, 5154.222, 5159.586, 
    5178.478,
  5300.766, 5273.486, 5255.66, 5251.909, 5255.065, 5261.641, 5260.849, 
    5252.441, 5237.964, 5222.568, 5204.3, 5185.364, 5167.836, 5156.462, 
    5166.951,
  5316.565, 5291.431, 5268.436, 5260.947, 5262.849, 5267.688, 5266.915, 
    5262.118, 5252.341, 5236.76, 5218.458, 5200.224, 5182.921, 5168.161, 
    5160.527,
  5331.409, 5310.228, 5284.712, 5268.99, 5267.037, 5270.329, 5272.144, 
    5267.415, 5258.735, 5246.475, 5231.126, 5214.292, 5197.223, 5182.7, 
    5170.245,
  5270.064, 5267.675, 5265.128, 5258.854, 5253.381, 5251.713, 5240.846, 
    5226.942, 5209.08, 5188.538, 5185.479, 5190.6, 5194.576, 5191.699, 
    5183.364,
  5256.793, 5256.167, 5256.442, 5254.365, 5255.193, 5251.025, 5243.029, 
    5224.011, 5205.502, 5190.277, 5185.805, 5190.138, 5192.281, 5188.785, 
    5178.927,
  5253.254, 5252.663, 5256.102, 5259.953, 5259.417, 5257.362, 5243.073, 
    5230.886, 5214.068, 5194.431, 5185.619, 5188.917, 5190.418, 5186.681, 
    5175.859,
  5260.184, 5259.55, 5264.568, 5267.074, 5267.267, 5258.08, 5251.332, 
    5233.727, 5215.384, 5199.902, 5185.869, 5185.763, 5189.41, 5185.963, 
    5176.72,
  5275.149, 5273.838, 5277.217, 5277.04, 5274.751, 5266.784, 5254.9, 
    5240.795, 5227.626, 5205.012, 5190.744, 5182.334, 5187.264, 5186.169, 
    5180.923,
  5289.078, 5287.169, 5286.555, 5284.845, 5280.09, 5271.676, 5262.099, 
    5246.758, 5230.195, 5213.764, 5196.082, 5182.148, 5185.699, 5188.254, 
    5185.645,
  5298.731, 5295.382, 5293.241, 5289.958, 5285.042, 5277.303, 5265.67, 
    5254.568, 5241.63, 5224.005, 5205.574, 5189.774, 5185.188, 5191.09, 
    5191.197,
  5305.384, 5297.905, 5293.75, 5289.516, 5284.477, 5278.258, 5269.026, 
    5257.838, 5245.674, 5232.729, 5216.889, 5200.639, 5190.549, 5192.436, 
    5196.6,
  5309.219, 5301.314, 5292.814, 5287.034, 5283.118, 5278.107, 5269.622, 
    5261.358, 5252.832, 5241.869, 5227.599, 5212.5, 5200.105, 5194.939, 
    5199.026,
  5309.423, 5303.17, 5295.175, 5285.39, 5279.958, 5276.499, 5270.491, 
    5262.646, 5253.885, 5246.086, 5236.304, 5223.812, 5210.983, 5202.108, 
    5200.666,
  5292.786, 5289.949, 5286.886, 5282.022, 5276.565, 5268.86, 5257.485, 
    5246.473, 5233.481, 5216.563, 5201.722, 5195.371, 5194.889, 5196.052, 
    5197.511,
  5300.417, 5295.289, 5290.951, 5284.609, 5277.604, 5266.998, 5258.464, 
    5242.595, 5228.651, 5214.152, 5199.282, 5194.016, 5195.172, 5196.744, 
    5196.291,
  5307.668, 5301.455, 5294.59, 5287.654, 5278.081, 5270.266, 5254.213, 
    5244.459, 5229.984, 5213.458, 5197.32, 5191.435, 5191.852, 5192.355, 
    5189.3,
  5309.027, 5302.145, 5294.956, 5285.942, 5275.964, 5264.338, 5255.741, 
    5239.605, 5227.246, 5214.071, 5197.379, 5188.354, 5186.611, 5185.743, 
    5180.787,
  5308.558, 5301.504, 5293.857, 5283.24, 5273.884, 5264.318, 5250.834, 
    5241.357, 5230.293, 5214.254, 5199.056, 5186.444, 5182.754, 5178.45, 
    5172.826,
  5305.943, 5298.516, 5290.137, 5279.504, 5270.205, 5261.787, 5251.7, 
    5238.557, 5227.437, 5216.034, 5201.079, 5187.119, 5179.921, 5172.722, 
    5164.136,
  5303.886, 5297.479, 5289.104, 5278.658, 5271.508, 5263.628, 5252.39, 
    5242.646, 5231.547, 5218.126, 5203.261, 5188.917, 5176.952, 5167.724, 
    5154.82,
  5302.237, 5296.907, 5289.825, 5281.124, 5274.191, 5267.417, 5256.964, 
    5244.303, 5231.409, 5220.023, 5206.194, 5191.593, 5176.451, 5164.102, 
    5148.578,
  5300.664, 5298.1, 5293.997, 5288.116, 5282.829, 5275.597, 5264.037, 
    5251.755, 5237.548, 5223.431, 5209.295, 5195.166, 5178.845, 5162.327, 
    5145.273,
  5299.888, 5297.9, 5297.629, 5294.847, 5290.104, 5283.349, 5272.108, 
    5257.19, 5241.406, 5226.143, 5212.401, 5199.39, 5183.288, 5164.459, 
    5146.054,
  5336.579, 5324.366, 5313.89, 5302.496, 5290.613, 5278.035, 5264.065, 
    5252.198, 5240.142, 5227.128, 5215.689, 5204.242, 5197.083, 5193.694, 
    5191.296,
  5334.757, 5321.566, 5310.424, 5298.353, 5286.537, 5271.751, 5261.343, 
    5244.561, 5232.336, 5222.88, 5212.047, 5200.989, 5194.294, 5191.417, 
    5191.07,
  5334.234, 5321.61, 5310.323, 5299.539, 5285.504, 5275.289, 5255.679, 
    5246.019, 5231.431, 5218.73, 5208.026, 5198.174, 5190.108, 5185.906, 
    5184.508,
  5335.187, 5322.669, 5312.094, 5300.111, 5287.978, 5271.824, 5260.086, 
    5239.246, 5226.306, 5215.281, 5204.068, 5194.416, 5185.43, 5179.682, 
    5175.955,
  5336.336, 5325.223, 5316.275, 5304.973, 5292.91, 5277.624, 5258.091, 
    5243.619, 5227.876, 5210.533, 5200.244, 5188.561, 5180.375, 5172.062, 
    5167.739,
  5337.64, 5327.82, 5319.547, 5309.351, 5295.71, 5279.622, 5261.857, 
    5240.469, 5222.987, 5208.395, 5194.782, 5182.205, 5173.4, 5164.388, 
    5159.522,
  5338.556, 5331.29, 5324.156, 5314.135, 5300.988, 5284.246, 5263.949, 
    5245.158, 5226.527, 5206.42, 5190.208, 5176.399, 5165.396, 5155.485, 
    5150.001,
  5340.562, 5334.075, 5326.455, 5316.729, 5302.24, 5285.766, 5266.312, 
    5244.749, 5224.378, 5205.409, 5186.879, 5169.851, 5156.272, 5145.106, 
    5139.018,
  5343.27, 5337.612, 5329.916, 5319.299, 5305.594, 5288.678, 5268.464, 
    5248.761, 5228.373, 5206.412, 5184.469, 5163.729, 5146, 5132.194, 5126.265,
  5348.697, 5340.637, 5331.583, 5320.688, 5305.061, 5287.743, 5269.023, 
    5248.486, 5228.318, 5206.753, 5183.243, 5158.891, 5137.473, 5121.797, 
    5117.767,
  5339.441, 5327.639, 5318.339, 5305.983, 5292.312, 5276.251, 5258.632, 
    5244.766, 5231.084, 5216.526, 5206.402, 5198.561, 5193.404, 5191.076, 
    5191.738,
  5337.585, 5326.02, 5315.432, 5301.428, 5286.368, 5267.413, 5254.93, 
    5234.998, 5222.218, 5211.752, 5200.791, 5192.459, 5186.502, 5184.458, 
    5184.682,
  5337.227, 5325.6, 5313.036, 5298.128, 5279.88, 5266.337, 5243.137, 
    5235.318, 5218.076, 5205.317, 5194.542, 5185.785, 5178.318, 5175.216, 
    5175.458,
  5336.949, 5322.871, 5308.265, 5290.291, 5272.124, 5251.295, 5240.221, 
    5217.741, 5208.597, 5198.021, 5186.868, 5176.982, 5169.078, 5165.311, 
    5165.525,
  5336.389, 5320.76, 5303.374, 5282.549, 5262.247, 5243.066, 5223.13, 
    5214.357, 5199.519, 5186.834, 5177.408, 5165.456, 5157.49, 5152.505, 
    5154.083,
  5335.432, 5316.266, 5293.666, 5270.203, 5245.998, 5225.152, 5208.989, 
    5193.06, 5183.223, 5175.302, 5163.881, 5152.61, 5143.12, 5139.406, 
    5141.607,
  5333.326, 5310.815, 5282.757, 5254.576, 5228.051, 5205.627, 5189.803, 
    5181.063, 5172.401, 5161.395, 5150.617, 5137.267, 5126.159, 5124.427, 
    5129.555,
  5330.636, 5301.429, 5267.018, 5235.195, 5205.295, 5185.044, 5172.309, 
    5163.339, 5157.009, 5149.588, 5136.952, 5120.993, 5109.977, 5112.015, 
    5121.312,
  5327.836, 5294.282, 5255.954, 5219.972, 5190.347, 5170.787, 5160.279, 
    5155.943, 5150.088, 5139.354, 5124.387, 5106.537, 5099.521, 5107.368, 
    5120.009,
  5328.132, 5288.136, 5246.796, 5209.573, 5178.818, 5160.738, 5153.25, 
    5148.404, 5142.862, 5133.227, 5117.411, 5104.531, 5105.314, 5115.325, 
    5128.44,
  5300.11, 5288.958, 5280.089, 5271.908, 5265.716, 5259.091, 5252.855, 
    5249.483, 5244.771, 5238.82, 5235.761, 5230.974, 5225.025, 5218.289, 
    5214.984,
  5282.122, 5269.368, 5258.116, 5248.252, 5240.283, 5233.639, 5232.143, 
    5224.508, 5224.038, 5224.657, 5222.499, 5222.292, 5220.279, 5217.389, 
    5216.264,
  5265.633, 5250.712, 5236.826, 5225.809, 5213.983, 5209.94, 5197.404, 
    5204.143, 5197.439, 5201.415, 5205.875, 5210.155, 5212.464, 5213.417, 
    5214.522,
  5253.701, 5235.521, 5219.018, 5202.163, 5188.639, 5174.086, 5173.407, 
    5159.52, 5169.495, 5173.953, 5184.117, 5192.809, 5202.002, 5207.371, 
    5212.694,
  5245.535, 5224.637, 5204.425, 5184.776, 5166.747, 5150.698, 5135.106, 
    5135.038, 5130.333, 5139.482, 5158.318, 5173, 5188.28, 5197.902, 5208.053,
  5242.107, 5218.424, 5194.256, 5171.896, 5148.704, 5130.686, 5116.31, 
    5103.205, 5103.18, 5113.054, 5128.765, 5152.476, 5172.507, 5188.88, 
    5201.668,
  5242.738, 5218.859, 5193.604, 5170.122, 5147.302, 5126.12, 5109.1, 5100.41, 
    5093.195, 5095.066, 5111.982, 5136.089, 5157.991, 5178.377, 5194.288,
  5249.054, 5225.205, 5199.436, 5175.792, 5150.156, 5129.089, 5112.128, 
    5100.6, 5094.506, 5095.814, 5105.13, 5125.471, 5147.841, 5169.226, 5187.99,
  5259.887, 5236.876, 5211.849, 5187.938, 5162.417, 5137.124, 5117.964, 
    5108.82, 5101.354, 5097.923, 5104.066, 5120.566, 5139.587, 5161.292, 
    5182.302,
  5275.113, 5250.408, 5226.277, 5200.328, 5169.975, 5142.843, 5122.835, 
    5111.121, 5107.453, 5104.344, 5108.429, 5120.447, 5136.622, 5157.937, 
    5180.747,
  5275.029, 5262.151, 5250.612, 5239.976, 5231.156, 5223.279, 5217.033, 
    5215.503, 5215.283, 5217.292, 5224.909, 5234.424, 5244.205, 5250.41, 
    5251.077,
  5271.85, 5256.431, 5242.21, 5228.72, 5217.149, 5206.265, 5201.593, 
    5194.795, 5196.1, 5201.173, 5208.753, 5221.943, 5233.914, 5244.593, 
    5246.437,
  5270, 5252.206, 5235.832, 5220.979, 5206.134, 5197.495, 5183.72, 5183.801, 
    5178.795, 5184.122, 5195.205, 5210.788, 5226.522, 5239.014, 5243.787,
  5263.608, 5243.159, 5224.115, 5205.436, 5190.842, 5176.163, 5173.021, 
    5161.126, 5164.323, 5167.118, 5180.706, 5199.467, 5220.223, 5235.371, 
    5242.957,
  5256.303, 5233.58, 5210.993, 5190.243, 5172.388, 5159.778, 5148.768, 
    5151.468, 5148.305, 5152.404, 5167.424, 5189.584, 5214.994, 5232.446, 
    5243.522,
  5247.747, 5221.231, 5194.365, 5170.6, 5149.87, 5135.923, 5129.278, 
    5126.814, 5133.641, 5141.512, 5154.261, 5182.346, 5210.685, 5232.355, 
    5245.451,
  5239.517, 5210.895, 5180.397, 5153.459, 5130.851, 5115.242, 5107.884, 
    5113.172, 5120.819, 5129.738, 5146.018, 5176.952, 5208.963, 5233.021, 
    5250.121,
  5233.101, 5201.188, 5166.983, 5138.645, 5113.185, 5098.039, 5092.789, 
    5097.172, 5109.604, 5123.26, 5140.583, 5175.293, 5210.367, 5236.512, 
    5257.461,
  5228.859, 5195.715, 5160.672, 5130.939, 5106.15, 5090.942, 5086.288, 
    5095.247, 5107.999, 5119.76, 5140.681, 5178.631, 5214.098, 5242.373, 
    5266.523,
  5228.664, 5192.932, 5158.326, 5129.496, 5105.616, 5091.974, 5089.897, 
    5096.475, 5108.505, 5121.511, 5147.522, 5186.444, 5221.878, 5251.399, 
    5277.694,
  5276.955, 5254.873, 5237.14, 5223.667, 5215.466, 5210.353, 5208.551, 
    5210.5, 5212.99, 5214.692, 5218.232, 5222.7, 5231.211, 5243.055, 5259.118,
  5254.396, 5231.365, 5213.945, 5201.319, 5194.437, 5190.979, 5192.788, 
    5193.454, 5199.039, 5206.227, 5210.262, 5215.374, 5221.488, 5235.073, 
    5250.102,
  5231.849, 5208.621, 5191.687, 5180.691, 5174.095, 5175.317, 5172.923, 
    5182.894, 5186.613, 5194.678, 5201.57, 5207.968, 5214.691, 5225.961, 
    5241.887,
  5209.736, 5186.732, 5170.661, 5158.663, 5153.375, 5150.823, 5159.545, 
    5159.338, 5172.717, 5183.251, 5193.67, 5201.31, 5210.312, 5222.273, 
    5237.581,
  5189.047, 5166.959, 5150.313, 5139.151, 5133.023, 5132.198, 5135.335, 
    5149.923, 5159.583, 5172.228, 5185.868, 5196.082, 5207.686, 5219.961, 
    5235.046,
  5171.162, 5148.982, 5132.425, 5121.261, 5113.801, 5112.474, 5119.006, 
    5129.209, 5146.494, 5165.57, 5178.735, 5193.764, 5207.085, 5222.417, 
    5235.937,
  5154.929, 5134.455, 5118.322, 5108.142, 5101.486, 5099.076, 5104.09, 
    5121.984, 5141.314, 5159.208, 5177.362, 5193.65, 5210.54, 5226.248, 
    5239.161,
  5142.598, 5123.275, 5107.917, 5099.043, 5092.26, 5090.082, 5096.957, 
    5112.189, 5134.776, 5159.228, 5177.665, 5197.679, 5217.291, 5232.719, 
    5245.57,
  5134.191, 5116.488, 5102.655, 5094.751, 5089.499, 5088.377, 5096.137, 
    5117.465, 5141.123, 5162.803, 5183.714, 5206.846, 5225.352, 5240.569, 
    5254.452,
  5130.744, 5113.361, 5101.208, 5094.772, 5090.198, 5092.09, 5103.776, 
    5123.147, 5146.77, 5171.24, 5195.023, 5217.893, 5236.097, 5252.878, 
    5269.723,
  5287.585, 5266.829, 5248.687, 5230.771, 5216.297, 5204.552, 5196.761, 
    5193.228, 5192.77, 5193.437, 5197.703, 5203.401, 5209.928, 5217.183, 
    5228.666,
  5252.384, 5229.483, 5210.3, 5192.422, 5180.141, 5171.99, 5172.007, 
    5171.353, 5175.834, 5183.365, 5191.476, 5200.604, 5209.959, 5221.446, 
    5234.967,
  5215.838, 5192.309, 5173.029, 5158.5, 5150.204, 5151.279, 5148.457, 
    5160.692, 5167.522, 5177.444, 5187.982, 5199.33, 5211.187, 5223.694, 
    5240.842,
  5178.622, 5157.074, 5139.885, 5129.512, 5125.273, 5127.136, 5140.198, 
    5144.607, 5159.021, 5172.564, 5186.871, 5199.385, 5213.384, 5228.508, 
    5246.966,
  5148.264, 5129.918, 5117.253, 5110.398, 5109.526, 5115.888, 5124.687, 
    5143.886, 5157.554, 5170.399, 5186.408, 5200.537, 5215.602, 5230.702, 
    5250.546,
  5126.176, 5111.094, 5099.716, 5096.011, 5096.995, 5104.848, 5120.93, 
    5134.794, 5152.09, 5170.639, 5186.598, 5202.927, 5218.009, 5234.679, 
    5253.57,
  5111.087, 5099.042, 5090.271, 5088.493, 5092.778, 5101.707, 5115.15, 
    5136.638, 5155.225, 5171.062, 5188.873, 5205.126, 5220.414, 5236.318, 
    5255.452,
  5103.031, 5093.073, 5085.504, 5086.122, 5090.073, 5100.525, 5116.13, 
    5133.325, 5152.293, 5173.093, 5191.362, 5208.094, 5223.698, 5240.17, 
    5259.843,
  5100.715, 5092.488, 5087.339, 5088.65, 5094.392, 5104.269, 5118.643, 
    5139.802, 5159.743, 5177.533, 5195.377, 5212.328, 5227.994, 5245.292, 
    5264.9,
  5104.21, 5094.902, 5090.997, 5092.984, 5098.388, 5109.633, 5126.18, 
    5144.527, 5163.55, 5183.566, 5201.722, 5218.393, 5234.759, 5252.943, 
    5273.105,
  5309.006, 5289.173, 5270.894, 5253.311, 5239.026, 5227.052, 5217.771, 
    5212.668, 5209.453, 5207.238, 5208.696, 5214.011, 5223.412, 5235.891, 
    5251.498,
  5272.919, 5250.58, 5230.335, 5211.53, 5197.751, 5186.285, 5182.162, 
    5176.312, 5175.231, 5179.427, 5185.154, 5197.582, 5213.425, 5235.262, 
    5255.602,
  5237.296, 5214.599, 5194.46, 5180.026, 5167.15, 5165.054, 5154.007, 
    5159.743, 5158.715, 5165.433, 5174.961, 5192.354, 5214.169, 5239.083, 
    5263.406,
  5203.46, 5183.266, 5166.997, 5154.261, 5146.231, 5139.738, 5144.372, 
    5140.039, 5147.046, 5158.499, 5174.505, 5195.756, 5222.337, 5250.767, 
    5274.866,
  5178.228, 5160.986, 5146.534, 5136.394, 5131.288, 5129.449, 5130.158, 
    5139.756, 5152.217, 5161.748, 5182.643, 5206.722, 5236.109, 5262.538, 
    5288.084,
  5159.038, 5142.917, 5130.364, 5123.239, 5118.984, 5120.345, 5128.208, 
    5137.292, 5151.68, 5172.806, 5195.245, 5222.688, 5251.097, 5278.217, 
    5302.847,
  5144.494, 5131.855, 5121.995, 5116.931, 5115.949, 5120.125, 5130.072, 
    5148.781, 5167.413, 5187.624, 5211.974, 5239.478, 5266.484, 5293.74, 
    5318.078,
  5136.312, 5126.766, 5118.408, 5115.747, 5116.506, 5126.168, 5141.601, 
    5159.3, 5178.934, 5203.938, 5229.096, 5256.273, 5283.378, 5309.206, 
    5331.913,
  5134.539, 5127.827, 5121.777, 5122.035, 5127.485, 5139.944, 5156.823, 
    5177.023, 5198.699, 5221.249, 5246.299, 5272.776, 5298.465, 5322.784, 
    5342.68,
  5138.573, 5132.167, 5128.967, 5131.841, 5139.648, 5155.515, 5172.895, 
    5191.844, 5213.183, 5237.309, 5262.339, 5287.557, 5312.346, 5334.423, 
    5351.664,
  5384.3, 5360.994, 5338.706, 5313.687, 5291.472, 5270.933, 5253.62, 
    5242.823, 5234.172, 5227.582, 5226.032, 5227.863, 5234.183, 5245.438, 
    5260.401,
  5346.771, 5320.348, 5294.967, 5269.34, 5249.328, 5230.249, 5220.52, 
    5208.048, 5202.094, 5200, 5198.232, 5203.136, 5210.115, 5226.387, 5243.643,
  5305.859, 5279.559, 5254.201, 5234.654, 5214.278, 5205.932, 5186.41, 
    5186.698, 5177.803, 5178.378, 5179.456, 5185.99, 5196.395, 5213.486, 
    5236.349,
  5266.967, 5243.74, 5223.486, 5203.275, 5187.553, 5171.845, 5169.789, 
    5157.484, 5160.313, 5159.654, 5165.48, 5173.985, 5190.094, 5211.78, 
    5239.268,
  5238.415, 5218.819, 5198.215, 5180.302, 5165.344, 5154.945, 5146.251, 
    5148.425, 5147.109, 5151.247, 5159.773, 5172.552, 5194.481, 5220.011, 
    5251.254,
  5217.112, 5197.543, 5177.176, 5161.112, 5146.328, 5139.113, 5135.71, 
    5135.505, 5140.251, 5149.529, 5161.845, 5183.384, 5210.319, 5240.165, 
    5268.443,
  5199.503, 5182.104, 5162.872, 5149.279, 5138.54, 5133.293, 5131.569, 
    5137.914, 5145.379, 5159.151, 5180.437, 5207.423, 5235.863, 5263.587, 
    5289.132,
  5186.954, 5170.731, 5154.234, 5144.138, 5136.283, 5136.074, 5138.773, 
    5147.966, 5162.347, 5185.7, 5210.086, 5237.592, 5263.348, 5288.489, 
    5309.757,
  5179.715, 5167.229, 5156.332, 5151.461, 5149.444, 5151.986, 5159.449, 
    5174.899, 5195.667, 5218.002, 5242.678, 5267.469, 5291.129, 5311.742, 
    5328.487,
  5178.822, 5170.027, 5165.144, 5165.019, 5167.029, 5175.238, 5188.188, 
    5206.441, 5227.558, 5251.727, 5274.444, 5297.2, 5316.075, 5332.08, 
    5343.347,
  5474.637, 5461.804, 5445.409, 5421.892, 5394.461, 5361.68, 5326.402, 
    5298.247, 5271.093, 5248.6, 5235.162, 5229.26, 5228.868, 5231.91, 5237.285,
  5447.49, 5432.745, 5414.06, 5388.1, 5358.372, 5323.553, 5295.965, 5261.84, 
    5238.832, 5225.032, 5211.908, 5210.215, 5210.98, 5218.537, 5224.405,
  5421.681, 5406.626, 5383.939, 5358.043, 5323.728, 5299.894, 5255.244, 
    5240.078, 5210.805, 5199.013, 5190.922, 5192.706, 5195.635, 5203.811, 
    5213.439,
  5392.728, 5376.393, 5352.461, 5323.458, 5292.068, 5255.01, 5236.239, 
    5197.82, 5185.891, 5177.112, 5174.25, 5176.457, 5183.825, 5193.475, 
    5205.602,
  5361.596, 5345.132, 5320.314, 5292.755, 5260.305, 5231.168, 5197.442, 
    5187.198, 5168.871, 5159.746, 5161.974, 5165.372, 5175.424, 5185.902, 
    5201.771,
  5330.67, 5314.461, 5289.952, 5261.835, 5230.603, 5201.899, 5179.517, 
    5158.998, 5152.047, 5152.855, 5153.831, 5161.33, 5171.637, 5185.633, 
    5202.983,
  5303.781, 5288.127, 5262.71, 5236.976, 5208.732, 5184.032, 5164.412, 
    5155.877, 5150.39, 5148.992, 5154.154, 5163.423, 5175.304, 5191.886, 
    5212.307,
  5278.41, 5262.562, 5239.957, 5217.649, 5192.964, 5174.578, 5159.425, 
    5150.852, 5150.531, 5157.187, 5164.932, 5176.586, 5190.471, 5208.425, 
    5229.717,
  5256.57, 5244.238, 5227.986, 5211.17, 5193.869, 5179.997, 5172.261, 
    5172.371, 5175.797, 5181.613, 5190.878, 5202.268, 5215.356, 5231.937, 
    5252.188,
  5240.728, 5233.187, 5223.7, 5214.41, 5207.121, 5202.487, 5201.43, 5203.064, 
    5207.833, 5215.3, 5223.356, 5232.685, 5243.982, 5258.119, 5275.221,
  5385.678, 5394.238, 5405, 5413.973, 5422.636, 5426.488, 5426.658, 5425.574, 
    5418.598, 5403.975, 5387.628, 5367.057, 5345.285, 5325.028, 5309.861,
  5358.406, 5367.269, 5377.566, 5386.174, 5393.436, 5397.981, 5400.55, 
    5392.767, 5381.521, 5370.26, 5350.784, 5332.507, 5312.03, 5299.34, 
    5286.489,
  5335.752, 5345.492, 5355.052, 5365.656, 5371.385, 5378.241, 5366.771, 
    5368.037, 5348.271, 5331.793, 5312.778, 5295.468, 5278.328, 5267.194, 
    5262.961,
  5316.938, 5326.016, 5337.064, 5345.121, 5352.477, 5348.372, 5351.124, 
    5326.131, 5313.073, 5293.539, 5274.469, 5256.492, 5245.835, 5240.185, 
    5241.874,
  5301.464, 5311.081, 5322.125, 5329.995, 5333.278, 5331.806, 5315.25, 
    5306.434, 5281.101, 5250.77, 5238.413, 5221.553, 5217.737, 5216.622, 
    5226.146,
  5292.865, 5301.84, 5309.643, 5314.988, 5314.745, 5307.958, 5294.016, 
    5267.582, 5242.515, 5224.121, 5205.547, 5196.226, 5196.917, 5203.914, 
    5217.709,
  5288.194, 5296.08, 5301.859, 5304.368, 5301.853, 5290.89, 5270.261, 
    5248.936, 5223.606, 5197.774, 5184.484, 5182.534, 5187.766, 5199.766, 
    5218.294,
  5285.994, 5293.075, 5297.56, 5297.865, 5289.947, 5276.151, 5259.71, 
    5236.261, 5209.716, 5189.986, 5180.1, 5181.106, 5190.65, 5205.403, 
    5227.021,
  5287.085, 5294.159, 5296.054, 5291.977, 5283.35, 5276.071, 5262.407, 
    5244.109, 5218.292, 5194.629, 5185.674, 5188.096, 5198.148, 5215.323, 
    5239.834,
  5288.182, 5292.955, 5292.615, 5288.597, 5285.974, 5281.259, 5269.033, 
    5250.568, 5227.952, 5209.249, 5200.296, 5201.662, 5213.502, 5233.014, 
    5259.108,
  5386.936, 5361.53, 5341.679, 5327.037, 5318.035, 5312.896, 5310.941, 
    5313.696, 5317.432, 5321.788, 5328.091, 5336.528, 5345.527, 5356.077, 
    5367.639,
  5355.475, 5332.268, 5317.177, 5305.916, 5298.853, 5295.411, 5296.261, 
    5295.309, 5298.365, 5303.352, 5307.099, 5314.022, 5321.803, 5334.305, 
    5343.652,
  5331.721, 5314.661, 5303.702, 5295.858, 5290.12, 5289.607, 5285.508, 
    5288.785, 5286.969, 5288.105, 5291.642, 5297.098, 5303.642, 5312.667, 
    5324.982,
  5316.669, 5303.933, 5294.948, 5288.153, 5284.657, 5281.311, 5282.597, 
    5274.1, 5276.303, 5276.124, 5277.284, 5281.299, 5288.88, 5297.355, 
    5307.501,
  5307.157, 5297.756, 5291.316, 5286.663, 5281.322, 5277.916, 5270.633, 
    5267.02, 5258.518, 5255.02, 5258.159, 5261.637, 5269.87, 5278.012, 5290.27,
  5300.503, 5294.873, 5289.938, 5285.405, 5279.134, 5271.589, 5260.573, 
    5245.903, 5236.205, 5231.252, 5229.466, 5235.085, 5245.858, 5258.394, 
    5272.229,
  5297.806, 5295.771, 5291.819, 5285.497, 5275.853, 5262.287, 5245.13, 
    5227.379, 5209.206, 5197.67, 5197.397, 5205.446, 5218.663, 5236.327, 
    5254.938,
  5297.712, 5298.327, 5293.738, 5285.961, 5273.578, 5258.014, 5236.56, 
    5210.075, 5185.972, 5173.47, 5170.255, 5179.928, 5198.338, 5219.772, 
    5245.149,
  5302.017, 5303.169, 5297.337, 5287.583, 5274.206, 5255.549, 5230.953, 
    5203.528, 5179.966, 5168.086, 5166.589, 5174.345, 5191.645, 5217.007, 
    5245.904,
  5307.763, 5306.588, 5299.544, 5289.598, 5275.622, 5257.905, 5234.204, 
    5206.369, 5184.479, 5174.369, 5172.756, 5180.516, 5198.868, 5225.965, 
    5258.299,
  5479.059, 5471.021, 5463.071, 5448.407, 5432.143, 5413.135, 5393.068, 
    5375.271, 5355.886, 5334.06, 5316.902, 5303.662, 5294.542, 5289.6, 
    5290.786,
  5438.657, 5434.628, 5430.666, 5419.282, 5406.249, 5387.868, 5374.254, 
    5351.906, 5334.343, 5320.093, 5303.889, 5291.351, 5282.044, 5278.786, 
    5278.129,
  5398.179, 5399.556, 5397.786, 5391.953, 5379.821, 5370.537, 5347.214, 
    5339.759, 5318.329, 5300.69, 5287.047, 5278.915, 5272.829, 5270.516, 
    5270.292,
  5360.004, 5365.698, 5367.339, 5364.881, 5356.655, 5342.344, 5333.558, 
    5305.944, 5292.67, 5279.831, 5267.428, 5262.152, 5263.559, 5265.785, 
    5267.206,
  5340.5, 5345.826, 5347.297, 5344.76, 5336.521, 5325.409, 5304.856, 
    5296.101, 5272.492, 5250.786, 5245.178, 5245.826, 5258.634, 5263.687, 
    5268.719,
  5330.975, 5332.912, 5331.466, 5327.606, 5317.665, 5304.154, 5287.195, 
    5260.735, 5239.241, 5224.668, 5220.725, 5235.089, 5256.338, 5266.046, 
    5273.482,
  5323.754, 5323.821, 5320.544, 5313.549, 5302.989, 5286.319, 5266.58, 
    5245.438, 5222.072, 5200.782, 5205.165, 5231.915, 5256.688, 5271.319, 
    5281.58,
  5318.296, 5315.147, 5308.835, 5299.98, 5286.814, 5269.735, 5248.365, 
    5220.793, 5197.425, 5188.267, 5200.637, 5231.731, 5259.026, 5277.684, 
    5290.097,
  5308.401, 5305.621, 5299.917, 5290.413, 5276.253, 5256.297, 5232.729, 
    5209.198, 5191.869, 5185.639, 5204.176, 5236.571, 5264.884, 5284.749, 
    5299.509,
  5305.76, 5302.371, 5294.757, 5283.202, 5266.32, 5244.307, 5220.856, 
    5197.837, 5184.764, 5191.089, 5214.104, 5244.023, 5272.47, 5293.199, 
    5310.743,
  5362.576, 5337.509, 5318.756, 5305.106, 5300.518, 5302.663, 5313.227, 
    5331.871, 5352.422, 5368.3, 5378.917, 5379.694, 5372.52, 5359.038, 
    5343.454,
  5335.582, 5307.773, 5287.007, 5273.693, 5270.773, 5276.306, 5292.504, 
    5309.852, 5331.65, 5350.976, 5359.058, 5358.371, 5350.042, 5338.204, 
    5320.26,
  5320.191, 5289.967, 5270.112, 5258.859, 5257.144, 5267.487, 5277.131, 
    5302.458, 5320.612, 5334.373, 5340.029, 5337.926, 5328.057, 5313.625, 
    5299.011,
  5313.836, 5286.402, 5267.781, 5257.249, 5259.709, 5261.942, 5283.021, 
    5289.691, 5308.498, 5317.304, 5321.114, 5316.2, 5307.063, 5294.072, 
    5284.466,
  5314.515, 5292.521, 5276.912, 5269.37, 5267.266, 5274.849, 5277.805, 
    5290.587, 5299.013, 5299.026, 5303.798, 5295.686, 5288.41, 5280.583, 
    5277.522,
  5315.346, 5297.097, 5282.381, 5275.561, 5272.785, 5272.875, 5277.622, 
    5279.253, 5282.62, 5286.682, 5283.218, 5278.792, 5276.896, 5276.497, 
    5277.821,
  5313.384, 5298.85, 5286.37, 5277.839, 5272.919, 5272.375, 5271.199, 
    5272.743, 5273.283, 5269.801, 5267.831, 5269.711, 5272.857, 5278.48, 
    5286.002,
  5307.975, 5295.15, 5282.01, 5274.273, 5266.771, 5262.31, 5258.798, 
    5256.754, 5254.477, 5253.957, 5256.546, 5266.651, 5276.247, 5287.333, 
    5297.496,
  5302.019, 5290.731, 5278.442, 5268.885, 5260.093, 5253.836, 5247.884, 
    5246.326, 5242.884, 5243.715, 5255.675, 5272.182, 5285.714, 5299.102, 
    5310.236,
  5297.168, 5284.801, 5271.886, 5261.42, 5249.907, 5240.963, 5234.564, 
    5232.366, 5231.241, 5245.171, 5266.146, 5283.825, 5299.575, 5313.359, 
    5324.346,
  5514.575, 5473.435, 5435.478, 5396.912, 5363.134, 5329.664, 5295.004, 
    5267.668, 5248.63, 5237.238, 5240.592, 5254.625, 5272.016, 5285.569, 
    5298.152,
  5490.775, 5452.045, 5417.809, 5383.102, 5355.478, 5322.469, 5303.61, 
    5276.927, 5264.217, 5262.616, 5269.662, 5282.522, 5292.799, 5302.153, 
    5307.373,
  5467.877, 5433.286, 5401.578, 5373.948, 5347.674, 5329.402, 5305.121, 
    5295.233, 5289.869, 5290.892, 5296.945, 5304.79, 5310.388, 5311.755, 
    5310.01,
  5443.837, 5413.262, 5384.799, 5361.732, 5341.461, 5324.936, 5314.43, 
    5307.056, 5304.649, 5310.619, 5316.539, 5321.343, 5320.42, 5315.941, 
    5306.513,
  5421.105, 5392.693, 5369.666, 5350.363, 5336.487, 5326.688, 5317.075, 
    5315.323, 5321.021, 5324.158, 5329.185, 5331.187, 5326.684, 5315.439, 
    5302.851,
  5396.5, 5371.878, 5351.826, 5337.391, 5326.929, 5319.914, 5318.719, 
    5315.287, 5320.776, 5329.43, 5335.079, 5335.465, 5329.252, 5316.138, 
    5308.003,
  5373.479, 5352.707, 5333.198, 5323.012, 5316.844, 5314.469, 5314.375, 
    5319.038, 5323.619, 5331.387, 5336.248, 5338.481, 5329.688, 5320.302, 
    5318.297,
  5352.28, 5330.549, 5311.905, 5305.042, 5301.39, 5303.626, 5305.077, 
    5312.069, 5317.646, 5328.906, 5335.037, 5338.18, 5330.983, 5328.993, 
    5330.728,
  5332.022, 5308.016, 5289.998, 5283.803, 5284.795, 5291.028, 5295.999, 
    5305.155, 5314.359, 5324.635, 5332.663, 5334.752, 5335.329, 5339.655, 
    5342.173,
  5313.515, 5285.076, 5266.706, 5261.968, 5265.987, 5275.851, 5284.148, 
    5293.964, 5304.979, 5317.568, 5328.646, 5335.419, 5343.452, 5350.717, 
    5355.49,
  5613.039, 5586.1, 5555.892, 5519.273, 5484.822, 5449.135, 5417.746, 
    5395.184, 5381.773, 5369.491, 5356.932, 5331.802, 5307.542, 5288.726, 
    5276.276,
  5593.559, 5564.301, 5531.639, 5494.073, 5459.584, 5422.675, 5401.895, 
    5380.373, 5372.422, 5369.546, 5358.147, 5335.836, 5310.472, 5294.638, 
    5281.413,
  5572.927, 5540.702, 5505.724, 5469.623, 5432.939, 5412.351, 5377.433, 
    5373.022, 5367.359, 5370.544, 5359.209, 5339.812, 5315.451, 5298.926, 
    5285.479,
  5548.67, 5513.758, 5477.166, 5439.461, 5409.188, 5376.788, 5368.013, 
    5354.904, 5362.942, 5368.739, 5362.274, 5344.881, 5324.308, 5307.693, 
    5293.843,
  5522.342, 5485.946, 5448.071, 5413.866, 5382.429, 5360.783, 5346.438, 
    5351.762, 5364.812, 5368.619, 5364.969, 5351.655, 5334.96, 5319.934, 
    5306.434,
  5495.332, 5457.163, 5420.1, 5384.532, 5353.706, 5336.188, 5335.648, 
    5342.371, 5355.365, 5369.924, 5367.662, 5359.281, 5346.535, 5335.024, 
    5322.404,
  5468.865, 5433.178, 5393.964, 5359.35, 5331.47, 5323.044, 5327.333, 
    5344.094, 5360.3, 5370.855, 5372.185, 5366.994, 5358.172, 5349.083, 
    5338.519,
  5448.207, 5411.886, 5370.942, 5335.104, 5312.426, 5311.994, 5326.522, 
    5344.152, 5360.017, 5374.229, 5377.812, 5375.319, 5369.669, 5362.873, 
    5353.788,
  5431.905, 5396.607, 5354.936, 5322.458, 5306.971, 5313.149, 5332.038, 
    5351.484, 5368.048, 5380.505, 5384.781, 5384.636, 5381.169, 5375.781, 
    5367.563,
  5422.004, 5385.24, 5346.433, 5319.204, 5309.92, 5320.954, 5340.196, 
    5357.784, 5373.848, 5387.007, 5393.027, 5394.52, 5393.227, 5388.938, 
    5381.21,
  5616.679, 5587.196, 5557.678, 5520.15, 5480.566, 5437.066, 5397.127, 
    5367.821, 5353.668, 5344.96, 5334.973, 5321.39, 5308.903, 5302.354, 
    5298.731,
  5596.858, 5568.814, 5535.945, 5495.916, 5453.646, 5407.02, 5380.564, 
    5361.039, 5353.778, 5351.628, 5341.415, 5328.787, 5314.727, 5306.918, 
    5301.549,
  5578.498, 5549.083, 5514.515, 5473.597, 5428.292, 5399.504, 5363.83, 
    5364.561, 5361.564, 5360.945, 5350.242, 5339.446, 5324.773, 5313.418, 
    5304.245,
  5560.571, 5530.211, 5493.236, 5449.818, 5409.855, 5376.08, 5369.39, 
    5365.842, 5369.251, 5368.021, 5360.703, 5349.441, 5335.404, 5321.434, 
    5308.706,
  5543.623, 5511.546, 5473.753, 5433.213, 5397.692, 5378.192, 5371.794, 
    5377.469, 5382.284, 5376.528, 5370.516, 5357.995, 5344.701, 5328.246, 
    5313.348,
  5526.556, 5495.164, 5457.87, 5420.718, 5392.08, 5379.756, 5382.646, 
    5387.215, 5387.716, 5386.049, 5378.423, 5366.411, 5351.491, 5334.123, 
    5316.555,
  5511.99, 5481.775, 5446.788, 5417.399, 5398.289, 5394.416, 5395.716, 
    5400.663, 5400.764, 5395.8, 5386.583, 5373.975, 5357.312, 5338.996, 
    5318.626,
  5499.008, 5471.792, 5440.926, 5418.865, 5407.773, 5407.875, 5410.892, 
    5412.395, 5409.951, 5405.255, 5395.263, 5381.177, 5363.128, 5343.072, 
    5321.079,
  5489.453, 5466.182, 5439.704, 5426.326, 5423.171, 5424.098, 5424.725, 
    5424.957, 5422.304, 5415.311, 5403.964, 5388.309, 5368.766, 5347.245, 
    5323.813,
  5483.378, 5462.246, 5441.338, 5434.341, 5434.529, 5435.649, 5436.893, 
    5435.635, 5431.622, 5424.346, 5412.472, 5395.596, 5374.991, 5352.866, 
    5328.963,
  5589.954, 5562.534, 5535.387, 5503.277, 5470.018, 5444.811, 5431.008, 
    5421.411, 5409.024, 5390.622, 5371.287, 5350.359, 5330.02, 5309.993, 
    5294.739,
  5572.844, 5547.697, 5521.528, 5488.636, 5461.495, 5439.537, 5434.237, 
    5418.576, 5405.161, 5389.91, 5369.309, 5346.606, 5323.607, 5304.962, 
    5286.377,
  5558.862, 5533.607, 5509.257, 5479.892, 5454.984, 5445.904, 5429.774, 
    5424.104, 5407.877, 5388.543, 5365.509, 5341.701, 5316.879, 5295.55, 
    5276.694,
  5545.115, 5521.048, 5496.593, 5469.746, 5451.547, 5441.362, 5433.093, 
    5418.374, 5401.903, 5385.532, 5360.678, 5335.972, 5310.536, 5289.302, 
    5268.051,
  5531.379, 5509.062, 5485.407, 5462.406, 5451.979, 5442.297, 5430.753, 
    5421.007, 5405.67, 5380.274, 5357.34, 5330.372, 5306.211, 5281.904, 
    5260.846,
  5518.617, 5497.83, 5474.238, 5457.764, 5448.82, 5440.69, 5431.493, 
    5415.512, 5397.299, 5377.246, 5353.621, 5327.982, 5304.209, 5280.438, 
    5258.169,
  5506.193, 5487.507, 5466.248, 5454.631, 5449.745, 5441.711, 5430.804, 
    5417.791, 5399.43, 5375.627, 5352.455, 5329.276, 5305.95, 5283.386, 
    5260.877,
  5496.355, 5478.761, 5460.01, 5453.299, 5448.773, 5441.724, 5431.144, 
    5414.55, 5394.845, 5374.987, 5354.626, 5333.938, 5313.5, 5292.831, 
    5271.572,
  5489.084, 5472.99, 5457.398, 5453.772, 5450.76, 5443.352, 5431.83, 
    5416.654, 5397.756, 5377.492, 5358.945, 5341.828, 5324.673, 5306.525, 
    5287.753,
  5484.512, 5469.238, 5456.678, 5456.154, 5451.962, 5444.635, 5432.732, 
    5415.848, 5397.521, 5380.271, 5365.017, 5351.271, 5338.127, 5324.15, 5309,
  5566.935, 5534.088, 5501.464, 5470.969, 5446.318, 5425.045, 5408.752, 
    5397.098, 5384.746, 5367.338, 5351.1, 5334.15, 5318.195, 5300.707, 5286.8,
  5551.78, 5517.146, 5483.941, 5455.402, 5433.359, 5413.324, 5404.116, 
    5386.661, 5373.021, 5358.335, 5342.062, 5326.648, 5309.765, 5293.336, 
    5275.566,
  5537.731, 5501.604, 5469.695, 5445.307, 5424.248, 5413.166, 5394.086, 
    5386.449, 5367.823, 5351.049, 5336.302, 5322.708, 5305.504, 5286.792, 
    5267.379,
  5522.445, 5486.606, 5458.556, 5435.859, 5419.136, 5403.75, 5394.693, 
    5373.216, 5358.483, 5346.783, 5334.561, 5321.724, 5304.618, 5285.779, 
    5265.312,
  5508.695, 5475.45, 5451.062, 5431.745, 5418.01, 5404.208, 5385.854, 
    5374.489, 5357.473, 5343.904, 5335.035, 5321.979, 5306.259, 5286.861, 
    5268.087,
  5496.43, 5466.777, 5445.36, 5429.711, 5415.023, 5400.212, 5384.836, 
    5365.19, 5351.771, 5344.939, 5335.643, 5323.78, 5308.298, 5290.992, 
    5272.552,
  5487.138, 5461.989, 5442.95, 5429.63, 5415.91, 5400.044, 5381.989, 
    5367.857, 5354.972, 5344.847, 5335.782, 5324.005, 5308.945, 5293.121, 
    5276.329,
  5480.539, 5458.43, 5441.783, 5429.926, 5413.999, 5398.701, 5381.67, 
    5364.973, 5352.318, 5344.413, 5334.643, 5322.443, 5308.333, 5293.641, 
    5279.444,
  5476.89, 5458.104, 5443.169, 5431.218, 5416.296, 5400.265, 5382.726, 
    5368.563, 5355.029, 5343.08, 5331.689, 5318.905, 5304.974, 5291.422, 
    5279.872,
  5475.894, 5458.243, 5445.698, 5434.133, 5417.895, 5401.991, 5384.782, 
    5367.444, 5352.458, 5339.723, 5327.102, 5314.095, 5301.191, 5289.036, 
    5279.4,
  5569.098, 5531.782, 5494.471, 5462.472, 5441.341, 5421.383, 5400.716, 
    5384.721, 5368.502, 5351.862, 5345.648, 5344.216, 5341.725, 5335.788, 
    5327.692,
  5556.294, 5517.998, 5482.311, 5455.271, 5435.149, 5412.085, 5397.282, 
    5372.42, 5357.811, 5348.636, 5343.025, 5341.519, 5339.131, 5334.434, 
    5326.279,
  5545.083, 5507.402, 5473.926, 5452.106, 5429.163, 5412.386, 5383.464, 
    5374.123, 5353.201, 5341.999, 5337.609, 5336.081, 5333.672, 5330.256, 
    5323.121,
  5533.149, 5496.789, 5467.731, 5445.897, 5423.903, 5399.131, 5382.853, 
    5354.867, 5342.486, 5333.668, 5327.942, 5326.816, 5325.206, 5323.271, 
    5318.209,
  5523.092, 5488.958, 5464.705, 5442.521, 5420.097, 5396.122, 5370.287, 
    5354.833, 5334.663, 5320.202, 5316.169, 5313.302, 5313.496, 5311.874, 
    5310.008,
  5514.015, 5482.58, 5460.928, 5438.289, 5413.617, 5388.616, 5364.654, 
    5338.132, 5319.162, 5307.824, 5299.613, 5298.099, 5298.427, 5298.783, 
    5298.643,
  5507.223, 5479.926, 5459.391, 5436.201, 5411.757, 5384.253, 5356.245, 
    5332.537, 5310.514, 5293.335, 5284.96, 5282.128, 5282.208, 5283.866, 
    5285.089,
  5502.095, 5477.839, 5457.358, 5434.018, 5406.971, 5378.777, 5349.249, 
    5319.902, 5296.345, 5281.315, 5271.62, 5267.542, 5267.502, 5269.749, 
    5272.379,
  5499.949, 5479.095, 5458.456, 5434.757, 5408.078, 5377.019, 5344.99, 
    5316.301, 5291.151, 5272.539, 5262.416, 5257.217, 5254.961, 5256.248, 
    5259.687,
  5500.547, 5480.434, 5460.66, 5437.358, 5408.007, 5377.252, 5345.794, 
    5314.091, 5288.107, 5269.776, 5257.771, 5250.516, 5247.037, 5246.835, 
    5249.836,
  5543.875, 5510.218, 5479.23, 5451.689, 5427.705, 5403.568, 5378.557, 
    5360.312, 5344.108, 5328.703, 5322.453, 5321.354, 5325.769, 5331.902, 
    5334.466,
  5529.141, 5496.139, 5467.322, 5440.252, 5414.755, 5385.305, 5367.532, 
    5340.551, 5325.25, 5315.511, 5309.594, 5310.907, 5317.256, 5327.809, 
    5333.181,
  5517.105, 5486.245, 5459.437, 5433.03, 5403.141, 5381.354, 5345.759, 
    5334.666, 5312.501, 5299.741, 5294.448, 5298.208, 5306.213, 5320.713, 
    5330.299,
  5507.599, 5478.82, 5452.802, 5423.438, 5393.323, 5359.553, 5340.932, 
    5308.103, 5295.257, 5285.329, 5280.728, 5284.943, 5295.468, 5312.937, 
    5327.064,
  5501.166, 5475.378, 5449.755, 5418.761, 5386.269, 5354.071, 5319.608, 
    5303.815, 5284.367, 5269.311, 5266.804, 5271.246, 5284.382, 5303.308, 
    5322.979,
  5497.545, 5473.678, 5446.952, 5414.712, 5378.128, 5342.214, 5310.681, 
    5282.099, 5265.924, 5259.12, 5255.888, 5262.05, 5275.012, 5296.488, 
    5318.125,
  5496.735, 5475.127, 5448.339, 5415.443, 5378.255, 5337.745, 5299.923, 
    5276.308, 5260.981, 5250.21, 5249.165, 5255.75, 5267.804, 5290.396, 
    5314.145,
  5498.084, 5478.28, 5451.298, 5417.752, 5377.036, 5335.003, 5295.647, 
    5265.754, 5250.913, 5246.398, 5245.743, 5253.335, 5265.067, 5287.679, 
    5311.702,
  5501.57, 5483.902, 5458.106, 5426.708, 5387.624, 5342.314, 5298.13, 
    5268.531, 5252.018, 5245.715, 5244.142, 5252.299, 5264.643, 5287.032, 
    5311.613,
  5506.872, 5490.484, 5468.717, 5438.228, 5397.816, 5354.323, 5309.188, 
    5272.83, 5253.589, 5248.045, 5247.619, 5254.287, 5268.391, 5289.766, 
    5313.011,
  5462.864, 5446.002, 5429.719, 5407.245, 5379.789, 5350.747, 5321.835, 
    5302.299, 5292.426, 5290.683, 5296.401, 5307.507, 5320.896, 5337.447, 
    5353.432,
  5455.841, 5439.582, 5419.543, 5391.028, 5357.647, 5320.584, 5296.778, 
    5274.263, 5269.115, 5273.834, 5284.415, 5300.073, 5317.153, 5338.743, 
    5358.036,
  5451.818, 5434.231, 5409.217, 5375.63, 5334.752, 5305.42, 5265.491, 
    5257.553, 5251.96, 5261.542, 5274.986, 5294.522, 5315.296, 5338.702, 
    5360.584,
  5448.095, 5428.365, 5398.725, 5358.681, 5316.726, 5276.234, 5255.343, 
    5234.726, 5240.524, 5252.559, 5271.027, 5290.682, 5314.907, 5341.117, 
    5365.891,
  5445.759, 5423.615, 5390.148, 5346.739, 5304.192, 5266.782, 5237.457, 
    5230.122, 5237.947, 5249.859, 5269.185, 5290.231, 5316.689, 5342.674, 
    5370.325,
  5443.533, 5420.027, 5383.12, 5339.253, 5295.574, 5259.844, 5235.618, 
    5228.306, 5235.204, 5253.533, 5270.187, 5293.059, 5319.226, 5348.14, 
    5374.44,
  5442.681, 5419.03, 5380.662, 5338.072, 5297.517, 5264.669, 5242.412, 
    5238.251, 5247.7, 5259.187, 5275.459, 5298.797, 5324.828, 5353.347, 
    5379.148,
  5443.128, 5419.375, 5381.679, 5341.208, 5302.69, 5273.228, 5255.933, 
    5250.928, 5255.495, 5268.088, 5284.141, 5306.702, 5332.758, 5360.512, 
    5385.054,
  5445.396, 5422.968, 5387.361, 5350.238, 5316.257, 5288.988, 5271.681, 
    5268.093, 5271.641, 5280.989, 5295.722, 5319.079, 5342.988, 5368.745, 
    5390.485,
  5448.779, 5427.535, 5395.819, 5362.99, 5330.507, 5306.112, 5290.969, 
    5284.37, 5286.35, 5296.261, 5311.805, 5332.865, 5354.774, 5377.583, 
    5396.216,
  5452.634, 5426.56, 5400.36, 5371.704, 5342.372, 5314.523, 5292.417, 
    5280.141, 5278.935, 5287.796, 5304.759, 5328.945, 5350.547, 5375.26, 
    5401.013,
  5436.967, 5409.988, 5381.588, 5349.48, 5317.14, 5286.533, 5270.658, 
    5257.717, 5257.46, 5271.62, 5293.427, 5322.344, 5349.25, 5381.481, 5407.55,
  5422.065, 5394.865, 5363.928, 5330.173, 5295.805, 5275.447, 5248.16, 
    5244.768, 5247.372, 5264.573, 5290.052, 5321.814, 5354.564, 5386.842, 
    5415.243,
  5408.03, 5379.545, 5346.617, 5311.264, 5280.702, 5254.026, 5244.352, 
    5232.631, 5241.438, 5264.121, 5294.314, 5327.207, 5363.687, 5398.761, 
    5426.075,
  5394.652, 5365.938, 5332.286, 5298.492, 5271.932, 5250.887, 5237.729, 
    5236.084, 5255.165, 5270.898, 5304.958, 5338.556, 5376.668, 5408.561, 
    5436.705,
  5382.98, 5353.888, 5320.089, 5290.627, 5266.489, 5250.088, 5242.844, 
    5246.053, 5257.738, 5287.232, 5318.782, 5354.88, 5390.883, 5423.246, 
    5448.279,
  5373.317, 5345.102, 5313.621, 5288.756, 5269.357, 5258.274, 5252.759, 
    5260.692, 5281.391, 5305.765, 5337.153, 5372.398, 5405.396, 5435.849, 
    5460.396,
  5366.753, 5339.706, 5311.444, 5290.708, 5274.772, 5267.979, 5268.747, 
    5278.224, 5296.77, 5324.484, 5356.816, 5388.656, 5420.334, 5448.572, 
    5473.768,
  5363.697, 5339.17, 5315.688, 5297.988, 5286.855, 5283.514, 5286.47, 
    5300.473, 5321.414, 5346.015, 5374.425, 5404.183, 5433.536, 5460.974, 
    5486.356,
  5364.663, 5342.596, 5323.053, 5308.528, 5299.791, 5299.248, 5305.901, 
    5318.669, 5337.672, 5362.91, 5390.504, 5418.224, 5446.186, 5473.045, 
    5498.513,
  5467.982, 5458.217, 5446.27, 5429.66, 5412.243, 5392.479, 5369.712, 
    5351.455, 5336.636, 5328.864, 5329.928, 5344.714, 5369.011, 5393.77, 
    5413.461,
  5450.536, 5438.287, 5422.533, 5404.595, 5384.221, 5359.787, 5340.349, 
    5321.404, 5306.559, 5306.299, 5313.825, 5337.179, 5366.596, 5397.502, 
    5417.8,
  5432.166, 5417.253, 5398.42, 5379.806, 5352.643, 5338.311, 5305.169, 
    5297.754, 5286.357, 5291.249, 5305.438, 5336.286, 5371.056, 5400.516, 
    5423.482,
  5412.419, 5393.195, 5373.234, 5348.305, 5326.33, 5298.564, 5290.722, 
    5270.732, 5271.884, 5282.432, 5307.261, 5342.584, 5380.104, 5409.64, 
    5433.459,
  5388.092, 5368.463, 5345.876, 5322.24, 5298.398, 5280.286, 5265.442, 
    5265.487, 5273.406, 5285.489, 5317.813, 5355.512, 5392.335, 5420.509, 
    5445.206,
  5364.258, 5343.751, 5320.465, 5297.185, 5276.437, 5262.768, 5257.731, 
    5260.602, 5271.533, 5298.972, 5334.759, 5372.899, 5407.189, 5435.82, 
    5458.134,
  5342.065, 5323.836, 5300.023, 5280.757, 5264.965, 5257.589, 5256.686, 
    5269.468, 5289.742, 5320.294, 5357.45, 5392.609, 5425.086, 5450.456, 
    5471.601,
  5326.958, 5307.55, 5286.7, 5272.575, 5262.255, 5262.139, 5269.474, 
    5285.714, 5310.786, 5346.818, 5381.799, 5414.549, 5443.154, 5466.078, 
    5486.237,
  5315.792, 5299.74, 5285.566, 5277.222, 5274.454, 5279.148, 5291.121, 
    5314.803, 5344.341, 5376.928, 5407.352, 5436.311, 5460.021, 5481.049, 
    5499.516,
  5313.879, 5300.967, 5293.058, 5290.149, 5292.983, 5304.044, 5323.155, 
    5347.14, 5375.208, 5405.026, 5431.868, 5455.851, 5476.896, 5496.87, 
    5514.28,
  5448.405, 5463.053, 5476.646, 5484.226, 5488.5, 5488.583, 5484.237, 
    5478.823, 5467.724, 5452.21, 5434.208, 5416.461, 5401.555, 5399.384, 
    5409.712,
  5444.398, 5456.942, 5465.997, 5471.131, 5472.476, 5469.891, 5466.438, 
    5454.387, 5442.743, 5429.269, 5411.141, 5394.283, 5387.606, 5398.192, 
    5411.836,
  5438.787, 5447.921, 5452.864, 5456.371, 5453.234, 5452.924, 5437.973, 
    5436.06, 5419.254, 5405.379, 5389.017, 5380.536, 5387.304, 5402.712, 
    5417.416,
  5429.539, 5433.55, 5435.526, 5433.506, 5431.206, 5421.472, 5420.64, 
    5400.576, 5393.021, 5382.847, 5374.791, 5378.263, 5395.937, 5412.302, 
    5427.601,
  5415.954, 5415.698, 5413.373, 5409.595, 5403.024, 5396.85, 5384.293, 
    5384.602, 5374.105, 5365.889, 5370.67, 5386.781, 5408.359, 5422.487, 
    5436.302,
  5393.22, 5389.254, 5382.875, 5376.799, 5368.35, 5362.407, 5357.314, 
    5351.313, 5351.939, 5360.062, 5376.498, 5400.822, 5419.92, 5436.918, 
    5449.748,
  5366.495, 5360.835, 5352.025, 5344.662, 5337.412, 5333.297, 5330.944, 
    5337.931, 5345.31, 5363.061, 5390.601, 5415.578, 5436.859, 5453.693, 
    5467.223,
  5338.708, 5330.479, 5319.347, 5312.1, 5306.72, 5307.657, 5313.269, 
    5322.872, 5344.019, 5377.292, 5408.208, 5434.605, 5456.359, 5472.644, 
    5487.145,
  5312.332, 5302.71, 5293.9, 5289.334, 5288.986, 5294.065, 5306.113, 
    5329.141, 5362.744, 5398.563, 5429.042, 5456.602, 5476.363, 5494.849, 
    5508.987,
  5293.047, 5284.34, 5278.674, 5276.888, 5280.872, 5292.967, 5314.293, 
    5347.364, 5386.815, 5422.751, 5453.19, 5478.375, 5499.184, 5516.495, 
    5530.795,
  5426.039, 5444.271, 5465.355, 5487.668, 5508.745, 5527.082, 5542.301, 
    5555.428, 5561.288, 5558.271, 5543.837, 5522.126, 5494.911, 5466.087, 
    5458.174,
  5417.563, 5438.173, 5460.161, 5483.686, 5504.047, 5522.32, 5538.472, 
    5548.037, 5551.418, 5546.594, 5530.68, 5504.863, 5472.801, 5453.852, 
    5447.3,
  5412.338, 5434.78, 5457.713, 5480.502, 5501.228, 5522.348, 5532.951, 
    5542.91, 5545.255, 5533.398, 5516.665, 5488.378, 5461.317, 5450.912, 
    5447.005,
  5410.537, 5432.18, 5455.644, 5476.368, 5499.414, 5514.665, 5531.41, 
    5532.757, 5531.857, 5521.915, 5502.659, 5476.923, 5464.714, 5458.271, 
    5458.533,
  5411.238, 5431.782, 5454.342, 5474.802, 5494.493, 5515.264, 5522.919, 
    5530.369, 5524.745, 5508.594, 5490.749, 5471.404, 5472.107, 5467.519, 
    5472.194,
  5413.628, 5431.333, 5450.78, 5469.796, 5488.421, 5505.125, 5516.342, 
    5517.707, 5510.334, 5498.258, 5479.837, 5473.161, 5478.385, 5478.804, 
    5483.636,
  5415.488, 5431.167, 5448.604, 5463.831, 5481.9, 5498.556, 5505.715, 
    5508.34, 5501.26, 5485.726, 5474.523, 5477.934, 5482.488, 5486.306, 
    5491.314,
  5414.194, 5428.349, 5441.529, 5455.505, 5470.954, 5486.321, 5494.721, 
    5495.44, 5487.4, 5477.286, 5474.996, 5482.298, 5486.966, 5492.462, 
    5497.805,
  5406.945, 5419.844, 5432.717, 5446.73, 5462.473, 5475.858, 5483.424, 
    5486.031, 5479.296, 5475.92, 5480.731, 5487.184, 5491.672, 5497.616, 
    5504.868,
  5392.877, 5405.096, 5417.356, 5432.644, 5448.59, 5463.668, 5472.472, 
    5475.958, 5475.745, 5481.614, 5489.227, 5494.706, 5500.825, 5507.911, 
    5515.81,
  5406.937, 5414.755, 5430.234, 5453.36, 5477.201, 5500.03, 5523.39, 
    5545.124, 5563.402, 5577.545, 5587.421, 5593.408, 5592.476, 5588.115, 
    5582.315,
  5407.522, 5416.307, 5433.146, 5456.132, 5476.417, 5499.469, 5521.476, 
    5541.873, 5556.807, 5571.01, 5577.521, 5580.235, 5575.106, 5569.204, 
    5558.396,
  5411.984, 5425.224, 5442.443, 5463.228, 5481.565, 5506.56, 5521.435, 
    5539.869, 5553.295, 5562.246, 5567.277, 5565.776, 5557.449, 5546.456, 
    5534.723,
  5421.51, 5434.938, 5452.297, 5468.918, 5490.574, 5503.373, 5526.262, 
    5534.413, 5547.847, 5554.619, 5555.625, 5549.54, 5539.799, 5527.684, 
    5514.284,
  5430.26, 5444.966, 5461.868, 5479.308, 5494.075, 5512.994, 5521.897, 
    5536.763, 5543.647, 5545.458, 5543.564, 5533.87, 5523.672, 5510.185, 
    5497.047,
  5437.338, 5453.265, 5468.518, 5484.374, 5497.305, 5509.458, 5525.514, 
    5533.489, 5538.698, 5537.493, 5529.508, 5518.094, 5509.775, 5498.426, 
    5485.908,
  5444.113, 5460.118, 5474.897, 5487.776, 5500.345, 5514.108, 5524.366, 
    5533.064, 5533.416, 5525.47, 5515.288, 5506.157, 5499.656, 5491.306, 
    5481.346,
  5450.305, 5465.893, 5479.207, 5490.668, 5502.305, 5515.465, 5528.034, 
    5530.2, 5524.591, 5512.957, 5502.979, 5498.655, 5495.773, 5490.653, 
    5484.289,
  5456.899, 5471.999, 5483.923, 5495.346, 5508.687, 5521.45, 5529.043, 
    5527.441, 5516.12, 5505.009, 5499.459, 5498.402, 5495.781, 5493.832, 
    5492.526,
  5464.248, 5476.688, 5487.612, 5499.297, 5513.114, 5526.767, 5532.445, 
    5526.155, 5513.951, 5506.66, 5502.715, 5500.561, 5500.028, 5499.914, 
    5500.975,
  5361.019, 5380.636, 5397.504, 5422.181, 5444.334, 5461.445, 5482.102, 
    5506.573, 5534.5, 5559.386, 5580.388, 5600.555, 5615.636, 5628.015, 
    5637.084,
  5361.899, 5378.096, 5394.929, 5418.898, 5439.244, 5459.111, 5478.438, 
    5499.843, 5524.028, 5550.961, 5570.714, 5588.715, 5602.304, 5614.591, 
    5620.863,
  5362.049, 5377.855, 5395.852, 5418.975, 5439.074, 5460.927, 5474.962, 
    5498.088, 5520.22, 5543.193, 5561.98, 5577.345, 5589.575, 5597.814, 
    5604.367,
  5369.667, 5382.869, 5401.273, 5420.927, 5442.233, 5456.986, 5480.825, 
    5492.414, 5514.264, 5534.634, 5553.298, 5566.314, 5576.529, 5583.267, 
    5586.738,
  5385.372, 5396.239, 5412.023, 5430.419, 5446.973, 5466.287, 5476.57, 
    5496.991, 5513.567, 5525.656, 5542.702, 5553.498, 5561.604, 5564.601, 
    5567.368,
  5409.9, 5417.638, 5427.923, 5442.412, 5455.202, 5468.043, 5484.326, 
    5494.769, 5506.602, 5522.364, 5531.232, 5540.575, 5546.306, 5547.453, 
    5546.902,
  5436.089, 5440.993, 5447.406, 5456.773, 5467.637, 5478.028, 5486.992, 
    5500.36, 5509.726, 5514.094, 5519.958, 5524.359, 5526.591, 5525.616, 
    5523.106,
  5457.675, 5460.219, 5464.004, 5470.164, 5476.723, 5485.334, 5493.271, 
    5496.785, 5499.881, 5503.989, 5505.539, 5506.715, 5506.958, 5506.497, 
    5503.699,
  5473.621, 5475.062, 5477.754, 5482.192, 5487.808, 5491.717, 5493.39, 
    5494.915, 5494.417, 5492.69, 5492.421, 5493.207, 5492.792, 5492.34, 
    5491.064,
  5485.208, 5486.519, 5489.419, 5493.212, 5496.323, 5498.69, 5497.949, 
    5494.694, 5490.99, 5490.277, 5490.172, 5489.08, 5487.706, 5487.112, 
    5486.777,
  5361.836, 5362.96, 5366.846, 5368.917, 5377.577, 5391.655, 5424.848, 
    5471.535, 5510.427, 5546.751, 5578.216, 5609.381, 5633.59, 5654.314, 
    5668.46,
  5371.448, 5372.174, 5369.06, 5373.499, 5377.172, 5387.747, 5419.227, 
    5465.429, 5504.069, 5544.107, 5576.463, 5606.23, 5629.959, 5649.714, 
    5662.099,
  5383.583, 5381.027, 5379.615, 5381.646, 5382.286, 5395.158, 5420.1, 
    5468.838, 5506.965, 5541.442, 5572.886, 5601.182, 5623.907, 5641.063, 
    5654.015,
  5402.757, 5399.226, 5396.456, 5394.857, 5398.175, 5398.695, 5433.525, 
    5465.219, 5503.318, 5539.159, 5567.983, 5593.786, 5615.83, 5632.638, 
    5643.375,
  5421.129, 5419.57, 5416.997, 5416.635, 5415.098, 5423.804, 5436.781, 
    5482.153, 5511.8, 5536.358, 5562.772, 5586.08, 5606.183, 5620.687, 
    5630.872,
  5437.405, 5437.588, 5435.81, 5434.973, 5435.447, 5437.663, 5457.307, 
    5480.312, 5503.351, 5535.11, 5555.523, 5578.274, 5594.77, 5608.288, 
    5615.958,
  5448.107, 5447.899, 5447.663, 5446.982, 5449.766, 5455, 5465.208, 5490.287, 
    5511.846, 5529.86, 5549.479, 5568.142, 5582.272, 5593.646, 5598.979,
  5456.977, 5456.002, 5455.486, 5456.673, 5458.646, 5465.314, 5476.094, 
    5488.084, 5502.713, 5523.695, 5541.171, 5556.033, 5569.295, 5578.255, 
    5582.762,
  5467.206, 5465.667, 5464.936, 5465.4, 5469.105, 5473.703, 5481.726, 
    5494.764, 5508.9, 5520.347, 5532.509, 5544.486, 5554.297, 5561.051, 
    5564.711,
  5478.273, 5474.992, 5473.703, 5473.382, 5474.646, 5478.656, 5484.949, 
    5490.954, 5499.979, 5511.528, 5522.104, 5530.709, 5538.701, 5543.931, 
    5546.688,
  5412.146, 5403.84, 5396.208, 5393.956, 5396.852, 5408.846, 5427.097, 
    5451.517, 5476.692, 5501.026, 5529.867, 5559.441, 5589.355, 5617.569, 
    5643.765,
  5410.001, 5399.517, 5389.437, 5385.593, 5384.546, 5395.87, 5414.981, 
    5437.572, 5463.785, 5495.922, 5528.971, 5560.798, 5592.051, 5622.405, 
    5647.263,
  5406.566, 5393.266, 5381.484, 5375.012, 5374.31, 5385.538, 5400.782, 
    5433.563, 5463.712, 5493.247, 5529.104, 5562.413, 5596.394, 5623.305, 
    5649.188,
  5399.403, 5384.528, 5370.56, 5360.728, 5358.308, 5366.289, 5395.825, 
    5416.807, 5453.149, 5490.244, 5530.741, 5564.482, 5600.159, 5627.825, 
    5651.361,
  5392.874, 5376.389, 5358.106, 5345.046, 5338.695, 5355.953, 5374.368, 
    5422.259, 5459.748, 5490.8, 5532.561, 5567.611, 5602.748, 5627.922, 
    5650.001,
  5388.642, 5369.047, 5345.142, 5324.691, 5318.634, 5336.52, 5374.274, 
    5409.354, 5449.338, 5495.811, 5534.732, 5572.231, 5603.802, 5629.387, 
    5648.449,
  5387.554, 5365.484, 5336.482, 5312.609, 5310.618, 5334.553, 5369.424, 
    5422.621, 5465.873, 5499.167, 5540.781, 5574.603, 5604.473, 5626.705, 
    5643.685,
  5392.349, 5369.982, 5341.478, 5321.411, 5319.843, 5346.5, 5384.313, 
    5423.703, 5462.23, 5506.031, 5544.531, 5575.938, 5603.839, 5623.532, 
    5638.035,
  5402.519, 5383.988, 5361.854, 5347.399, 5350.079, 5371.344, 5404.827, 
    5446.755, 5482.254, 5514.897, 5547.699, 5576.866, 5600.322, 5617.13, 
    5628.753,
  5417.17, 5403.766, 5389.383, 5380.603, 5382.771, 5402.051, 5428.114, 
    5456.324, 5485.736, 5519.447, 5550.626, 5575.474, 5595.682, 5609.678, 
    5618.475,
  5452.635, 5446.671, 5441.157, 5435.812, 5431.708, 5427.032, 5424.797, 
    5428.084, 5433.674, 5438.922, 5448.679, 5463.88, 5482.802, 5509.118, 
    5541.27,
  5434.813, 5427.14, 5420.651, 5415.624, 5413.446, 5412.555, 5413.357, 
    5414.546, 5421.801, 5432.445, 5443.509, 5461.111, 5481.518, 5509.593, 
    5540.54,
  5416.41, 5406.679, 5399.704, 5396.129, 5396.068, 5399.601, 5399.786, 
    5408.212, 5417.622, 5428.177, 5441.57, 5462.215, 5486.464, 5512.646, 
    5545.29,
  5397.676, 5385.52, 5377.192, 5373.303, 5377.287, 5382.579, 5393.827, 
    5394.607, 5408.534, 5424.815, 5442.77, 5466.454, 5492.489, 5522.408, 
    5554.297,
  5380.34, 5364.089, 5352.789, 5350.279, 5356.728, 5368.905, 5379.203, 
    5394.36, 5409.04, 5424.896, 5446.469, 5473.128, 5501.538, 5530.487, 
    5562.752,
  5362.155, 5339.356, 5319.648, 5316.632, 5331.21, 5351.679, 5372.124, 
    5384.479, 5402.14, 5428.185, 5451.812, 5481.657, 5510.186, 5542.589, 
    5572.542,
  5346.576, 5316.23, 5290.591, 5286.402, 5306.577, 5338.107, 5362.252, 
    5386.007, 5409.036, 5432.257, 5460.513, 5490.459, 5520.021, 5552.283, 
    5581.746,
  5340.014, 5306.636, 5279.729, 5275.145, 5297.396, 5333.125, 5361.697, 
    5382.445, 5408.003, 5440.102, 5469.612, 5500.195, 5531.054, 5563.757, 
    5591.463,
  5344.358, 5315.37, 5293.156, 5289.907, 5312.425, 5341.143, 5366.576, 
    5392.772, 5420.913, 5449.808, 5479.16, 5511.004, 5542.174, 5573.532, 
    5599.164,
  5359.032, 5336.87, 5321.943, 5320.689, 5335.076, 5355.729, 5377.85, 
    5399.563, 5427.497, 5458.517, 5489.846, 5521.851, 5553.228, 5582.393, 
    5606.17,
  5492.014, 5486.07, 5481.481, 5475.573, 5471.494, 5466.345, 5461.291, 
    5458.947, 5455.503, 5451.255, 5449.902, 5449.803, 5451.177, 5454.226, 
    5468.586,
  5468.798, 5462.3, 5456.706, 5450.757, 5445.871, 5442.185, 5441.823, 
    5437.242, 5436.445, 5437.05, 5435.686, 5438.497, 5441.986, 5448.349, 
    5462.79,
  5445.734, 5438.489, 5430.8, 5425.213, 5420.219, 5420.604, 5414.96, 
    5422.909, 5418.992, 5421.204, 5423.257, 5427.663, 5433.767, 5441.671, 
    5460.065,
  5423.504, 5413.83, 5404.55, 5396.788, 5393.001, 5391.761, 5400.256, 
    5396.392, 5405.384, 5407.467, 5413.102, 5419.262, 5428.314, 5440.243, 
    5463.138,
  5401.711, 5388.404, 5375.173, 5365.734, 5362.171, 5366.162, 5370.361, 
    5386.617, 5388.779, 5396.795, 5405.643, 5414.502, 5426.699, 5442.93, 
    5471.03,
  5380.753, 5363.344, 5345.722, 5332.588, 5328.523, 5337.69, 5353.074, 
    5364.518, 5378.609, 5391.281, 5401.823, 5415.548, 5430.328, 5453.854, 
    5483.422,
  5363.528, 5342.759, 5319.074, 5302.151, 5299.964, 5312.61, 5334.167, 
    5357.848, 5373.748, 5388.695, 5404.568, 5421.157, 5439.874, 5468.767, 
    5501.84,
  5352.317, 5329.472, 5302.008, 5283.924, 5283.695, 5302.951, 5329.85, 
    5352.272, 5373.76, 5393.848, 5412.934, 5430.892, 5456.479, 5488.96, 
    5521.901,
  5349.738, 5330.056, 5304.96, 5291.606, 5296.03, 5314.833, 5338.458, 
    5362.326, 5384.327, 5404.347, 5424.722, 5447.359, 5478.646, 5511.894, 
    5540.952,
  5355.122, 5341.597, 5325.729, 5317.181, 5321.208, 5335.26, 5354.5, 
    5374.928, 5398.105, 5420.735, 5442.036, 5469.926, 5502.75, 5533.768, 
    5561.142,
  5495.188, 5508.374, 5521.623, 5531.501, 5540.712, 5545.746, 5548.486, 
    5550.325, 5547.07, 5539.999, 5532.076, 5520.872, 5508.052, 5492.939, 
    5477.792,
  5483.209, 5492.945, 5502.664, 5511.696, 5517.979, 5523.907, 5527.602, 
    5526.561, 5526.091, 5525.08, 5517.184, 5509.955, 5499.499, 5489.692, 
    5474.432,
  5473.873, 5479.521, 5485.576, 5492.95, 5496.763, 5503.813, 5500.521, 
    5509.393, 5505.051, 5505.167, 5502.887, 5499.771, 5494.442, 5489.256, 
    5478.58,
  5460.929, 5464.018, 5466.448, 5468.872, 5472.27, 5472.822, 5482.261, 
    5475.273, 5486.287, 5486.859, 5489.447, 5490.474, 5492.022, 5490.813, 
    5487.254,
  5440.45, 5443.042, 5443.297, 5443.729, 5444.4, 5446.567, 5445.553, 
    5459.583, 5459.387, 5467.548, 5476.03, 5483.438, 5490.729, 5493.925, 
    5497.29,
  5420.557, 5419.532, 5417.017, 5414.825, 5411.055, 5411.992, 5416.811, 
    5421.477, 5437.323, 5452.604, 5463.913, 5478.811, 5490.835, 5499.956, 
    5506.917,
  5400.792, 5397.99, 5392.637, 5386.662, 5381.173, 5378.602, 5382.539, 
    5398.544, 5415.224, 5434.865, 5455.835, 5475.978, 5493.468, 5507.049, 
    5518.202,
  5385.817, 5381.149, 5373.277, 5364.375, 5354.423, 5350.833, 5354.395, 
    5368.67, 5394.004, 5424.755, 5449.791, 5475.423, 5498.514, 5516.267, 
    5529.236,
  5375.952, 5371.971, 5362.349, 5351.746, 5341.884, 5335.584, 5337.733, 
    5355.98, 5383.706, 5416.404, 5447.791, 5479.146, 5505.311, 5526.955, 
    5539.274,
  5374.031, 5368.532, 5359.068, 5349.349, 5338.916, 5332.304, 5332.82, 
    5348.638, 5379.098, 5416.776, 5452.47, 5486.277, 5516.598, 5538.865, 
    5549.656,
  5446.109, 5445.508, 5452.254, 5460.607, 5467.627, 5485.546, 5506.056, 
    5522.703, 5538.79, 5552.389, 5563.392, 5568.724, 5565.35, 5551.586, 
    5537.022,
  5449.068, 5447.619, 5455.409, 5465.531, 5472.492, 5488.425, 5504.127, 
    5518.568, 5533.942, 5549.296, 5559.642, 5563.379, 5557.123, 5544.998, 
    5530.363,
  5453.736, 5451.877, 5460.308, 5470.827, 5478.489, 5494.12, 5503.646, 
    5519.705, 5533.257, 5546.231, 5556.146, 5557.104, 5548.754, 5535.28, 
    5524.922,
  5457.645, 5457.201, 5465.375, 5472.814, 5485.377, 5491.574, 5509.578, 
    5517.119, 5533.453, 5544.446, 5551.5, 5548.484, 5540.146, 5529.465, 
    5520.918,
  5457.993, 5462.552, 5469.646, 5477.692, 5485.343, 5499.435, 5505.185, 
    5521.438, 5531.165, 5538.6, 5544.091, 5538.928, 5531.911, 5522.396, 
    5517.036,
  5451.312, 5462.084, 5470.415, 5477.924, 5485.941, 5493.935, 5508.793, 
    5515.587, 5525.393, 5533.729, 5534.296, 5529.813, 5524.195, 5518.69, 
    5514.457,
  5444.203, 5455.52, 5468.015, 5475.399, 5483.385, 5493.616, 5501.473, 
    5513.874, 5520.54, 5523.324, 5523.311, 5520.897, 5517.788, 5515.198, 
    5511.337,
  5431.915, 5442.558, 5457.662, 5469.002, 5475.039, 5486.028, 5495.098, 
    5502.007, 5507.255, 5512.354, 5512, 5512.165, 5513.017, 5514.112, 5509.816,
  5419.229, 5429.28, 5444.317, 5457.226, 5464.915, 5475.253, 5483.393, 
    5492.262, 5496.658, 5499.433, 5502.014, 5506.749, 5511.484, 5513.714, 
    5508.663,
  5408.248, 5415.851, 5427.995, 5442.07, 5451.922, 5462.231, 5471.194, 
    5477.959, 5483.86, 5490.713, 5497.506, 5505.674, 5512.685, 5514.975, 
    5509.331,
  5568.248, 5538.429, 5513.756, 5491.227, 5476.259, 5475.69, 5477.102, 
    5483.97, 5489.793, 5501.746, 5511.904, 5523.655, 5534.474, 5542.906, 
    5543.799,
  5566.415, 5542.133, 5520.6, 5503.062, 5492.374, 5489.096, 5488.631, 
    5492.294, 5497.891, 5509.049, 5519.029, 5532.104, 5541.75, 5545.379, 
    5539.066,
  5561.635, 5543.514, 5526.705, 5512.389, 5502.993, 5505.033, 5498.316, 
    5500.489, 5507.129, 5517.27, 5529.028, 5541.665, 5545.85, 5542.145, 
    5531.093,
  5552.032, 5539.029, 5528.463, 5515.549, 5510.527, 5504.608, 5508.632, 
    5508.164, 5515.912, 5527.078, 5539.828, 5546.87, 5545.705, 5536.663, 
    5520.71,
  5538.727, 5530.363, 5525.089, 5517.949, 5510.529, 5511.882, 5512.165, 
    5514.927, 5527.129, 5537.393, 5546.006, 5547.928, 5540.882, 5525.754, 
    5509.402,
  5520.726, 5516.688, 5515.503, 5513.74, 5511.477, 5511.237, 5516.349, 
    5524.283, 5532.737, 5544.133, 5548.631, 5544.481, 5532.521, 5515.777, 
    5499.964,
  5502.381, 5502.178, 5505.398, 5506.802, 5508.539, 5513.435, 5518.116, 
    5528.288, 5540.019, 5547.17, 5547.856, 5538.787, 5522.635, 5506.292, 
    5493.646,
  5482.623, 5484.735, 5491.869, 5497.94, 5502.494, 5509.798, 5520.601, 
    5531.084, 5541.7, 5548.546, 5544.07, 5530.088, 5513.877, 5502.407, 5491.96,
  5463.722, 5467.296, 5479.078, 5490.619, 5498.906, 5508.846, 5520.243, 
    5534.459, 5545.493, 5546.079, 5537.358, 5522.115, 5510.272, 5502.713, 
    5493.577,
  5443.897, 5449.028, 5463.233, 5480.205, 5493.014, 5507.477, 5521.261, 
    5534.733, 5542.395, 5541.946, 5530.674, 5519.29, 5512.735, 5506.556, 
    5501.323,
  5661.018, 5652.478, 5642.845, 5627.917, 5612.383, 5597.251, 5582.411, 
    5573.143, 5565.336, 5556.574, 5551.308, 5549.704, 5551.439, 5554.346, 
    5555.788,
  5643.371, 5637.388, 5631.542, 5619.564, 5607.515, 5593.781, 5584.814, 
    5573.624, 5566.501, 5562.425, 5559.742, 5560.22, 5560.605, 5559.101, 
    5554.509,
  5620.963, 5617.119, 5613.439, 5607.022, 5597.578, 5592.245, 5577.028, 
    5574.743, 5566.792, 5562.535, 5562.526, 5563.779, 5561.357, 5555.834, 
    5545.306,
  5590.722, 5590.206, 5589.167, 5587.219, 5583.44, 5577.07, 5575.086, 
    5563.39, 5561.659, 5561.172, 5562.013, 5562.113, 5557.562, 5546.979, 
    5531.561,
  5554.913, 5557.687, 5560.176, 5563.438, 5565.504, 5566.034, 5561.146, 
    5561.14, 5556.556, 5556.389, 5559.617, 5556.391, 5548.335, 5533.042, 
    5515.671,
  5513.226, 5518.16, 5524.327, 5534.501, 5541.951, 5548.731, 5550.442, 
    5549.704, 5550.774, 5553.269, 5553.57, 5548.893, 5537.163, 5520.023, 
    5503.21,
  5469.917, 5477.187, 5487.227, 5503.198, 5518.652, 5530.815, 5537.317, 
    5541.98, 5544.033, 5547.416, 5547.521, 5540.549, 5525.144, 5509.026, 
    5495.171,
  5439.719, 5448.063, 5458.749, 5476.841, 5496.045, 5514.027, 5524.585, 
    5530.932, 5536.569, 5543.034, 5541.214, 5530.834, 5515.516, 5502.408, 
    5489.514,
  5421.265, 5431.255, 5445.422, 5463.756, 5483.453, 5500.801, 5513.293, 
    5523.884, 5532.308, 5538.053, 5535.068, 5523.613, 5509.824, 5497.471, 
    5484.027,
  5404.596, 5414.667, 5431.811, 5452.109, 5472.466, 5489.835, 5504.442, 
    5516.887, 5528.31, 5535.348, 5529.816, 5518.841, 5507.875, 5494.702, 
    5482.426,
  5656.5, 5653.018, 5651.109, 5646.511, 5641.773, 5634.523, 5625.911, 
    5618.838, 5609.273, 5598.986, 5591.771, 5584.76, 5580.06, 5575.5, 5572.59,
  5636.984, 5633.116, 5630.188, 5625.049, 5619.132, 5612.368, 5607.753, 
    5598.126, 5593.007, 5587.935, 5580.43, 5575.617, 5571.29, 5568.435, 
    5563.413,
  5610.271, 5605.128, 5599.51, 5593.896, 5587.915, 5585.535, 5576.546, 
    5580.582, 5571.28, 5568.186, 5564.231, 5561.499, 5557.68, 5554.499, 
    5548.985,
  5580.783, 5573.085, 5565.011, 5557.726, 5551.872, 5547.396, 5551.609, 
    5541.893, 5548.667, 5547.503, 5545.943, 5544.503, 5542.576, 5540.232, 
    5533.506,
  5550.031, 5539.078, 5526.822, 5517.241, 5510.089, 5507.323, 5505.342, 
    5519.085, 5515.631, 5520.231, 5524.546, 5525.421, 5525.868, 5523.033, 
    5518.024,
  5512.523, 5495.996, 5478.27, 5466.077, 5457.513, 5458.795, 5465.024, 
    5470.355, 5484.481, 5496.894, 5500.934, 5507.493, 5508.435, 5507.523, 
    5502.203,
  5470.387, 5449.933, 5429.945, 5415.34, 5406.578, 5408.219, 5419.319, 
    5439.538, 5454.727, 5468.356, 5481.703, 5489.775, 5492.85, 5492.803, 
    5487.468,
  5428.436, 5404.575, 5378.326, 5362.051, 5354.197, 5363.508, 5382.45, 
    5404.407, 5428.134, 5450.715, 5465.077, 5475.358, 5479.777, 5478.493, 
    5475.087,
  5389.245, 5363.873, 5343.401, 5329.433, 5325.184, 5337.024, 5361.371, 
    5391.211, 5416.69, 5437.354, 5453.524, 5464.526, 5467.745, 5467.649, 
    5464.843,
  5359.455, 5342.927, 5332.187, 5320.009, 5312.565, 5327.594, 5354.391, 
    5383.197, 5410.711, 5434.267, 5448.941, 5457.293, 5459.004, 5459.439, 
    5464.192,
  5605.525, 5608.707, 5611.403, 5611.518, 5612.655, 5611.546, 5610.555, 
    5610.334, 5605.985, 5599.038, 5593.559, 5587.322, 5579.935, 5571.795, 
    5564.409,
  5582.136, 5585.456, 5587.214, 5586.618, 5584.847, 5582.833, 5581.122, 
    5573.474, 5570.404, 5568.755, 5562.646, 5558.51, 5553.427, 5549.014, 
    5542.616,
  5556.902, 5560.739, 5562.287, 5561.657, 5558.252, 5556.152, 5546.039, 
    5549.676, 5539.402, 5536.307, 5533.266, 5531.274, 5527.439, 5524.646, 
    5521.254,
  5531.831, 5534.147, 5533.872, 5531.435, 5526.411, 5521.657, 5521.035, 
    5506.888, 5507.633, 5504.583, 5501.154, 5499.845, 5499.923, 5499.235, 
    5497.605,
  5508.759, 5510.287, 5509.449, 5506.991, 5502.465, 5494.723, 5483.658, 
    5483.389, 5469.812, 5462.545, 5464.596, 5462.928, 5467.054, 5468.318, 
    5472.047,
  5492.751, 5491.072, 5485.671, 5477.915, 5465.743, 5454.161, 5441.334, 
    5425.002, 5418.831, 5416.069, 5414.232, 5419.376, 5426.955, 5435.33, 
    5443.317,
  5471.043, 5466.077, 5456.156, 5444.482, 5429.476, 5410.399, 5391.689, 
    5379.865, 5368.144, 5362.755, 5368.753, 5378.002, 5390.971, 5405.578, 
    5418.932,
  5450.317, 5440.869, 5426.836, 5409.129, 5387.293, 5365.933, 5345.025, 
    5328.329, 5322.884, 5327.018, 5334.833, 5348.931, 5367.189, 5386.541, 
    5404.072,
  5422.393, 5411.158, 5395.508, 5376.181, 5355.736, 5333.94, 5314.352, 
    5302.14, 5296.199, 5301.542, 5315.656, 5334.405, 5355.291, 5377.153, 
    5396.771,
  5400.318, 5388.382, 5373.575, 5358.151, 5339.932, 5318.831, 5296.733, 
    5281.059, 5280.803, 5292.971, 5311.029, 5331.991, 5355.401, 5377.725, 
    5397.352,
  5522.362, 5525.948, 5532.148, 5537.558, 5544.329, 5550.561, 5556.087, 
    5563.685, 5570.106, 5574.431, 5578.95, 5580.989, 5580.188, 5577.816, 
    5575.258,
  5489.116, 5490.65, 5493.911, 5498.773, 5502.764, 5510.58, 5519.47, 
    5524.283, 5532.744, 5542.84, 5547.864, 5552.55, 5553.422, 5554.362, 
    5549.582,
  5466.389, 5462.383, 5459.779, 5462.372, 5466.901, 5477.071, 5477.979, 
    5493.833, 5495.777, 5506.521, 5514.507, 5521.33, 5523.282, 5523.714, 
    5522.5,
  5452.137, 5449.02, 5446.683, 5444.68, 5446.21, 5447.436, 5458.419, 
    5454.344, 5466.993, 5474.009, 5481.031, 5486.825, 5491.506, 5492.211, 
    5489.874,
  5437.756, 5434.335, 5432.107, 5431.8, 5432.451, 5434.216, 5433.792, 
    5441.234, 5443.055, 5443.513, 5451.622, 5453.153, 5457.375, 5457.222, 
    5458.472,
  5424.225, 5422.032, 5419.927, 5419.229, 5418.716, 5419.631, 5422.25, 
    5419.209, 5420.602, 5422.971, 5421.314, 5422.052, 5424.043, 5424.422, 
    5425.005,
  5413.688, 5412.339, 5410.996, 5409.081, 5408.119, 5406.117, 5403.221, 
    5402.281, 5397.674, 5391.573, 5389.758, 5388.403, 5388.798, 5390.854, 
    5393.7,
  5404.23, 5403.99, 5402.606, 5400.824, 5397.461, 5393.808, 5388.19, 
    5379.161, 5370.582, 5363.692, 5357.863, 5355.71, 5358.209, 5362.432, 
    5369.203,
  5391.953, 5390.498, 5387.814, 5384.761, 5380.116, 5374.062, 5365.824, 
    5356.32, 5343.176, 5331.351, 5325.01, 5326.121, 5331.094, 5341.608, 
    5353.836,
  5381.535, 5378.357, 5374.622, 5370.564, 5364.542, 5357.848, 5348.613, 
    5334.16, 5317.629, 5306.425, 5302.291, 5306.002, 5317.541, 5332.683, 
    5351.854,
  5572.342, 5576.714, 5582.497, 5585.302, 5587.961, 5585.773, 5579.62, 
    5573.836, 5562.922, 5546.793, 5533.692, 5521.067, 5509.807, 5501.652, 
    5498.804,
  5545.964, 5551.485, 5555.909, 5557.082, 5555.794, 5552.059, 5547.985, 
    5532.769, 5521.979, 5510.34, 5494.33, 5481.907, 5471.193, 5466.719, 
    5460.753,
  5518.629, 5524.211, 5526.853, 5527.609, 5525.124, 5524.542, 5509.206, 
    5509.588, 5489.334, 5474.697, 5460.217, 5448.558, 5437.545, 5432.675, 
    5431.297,
  5490.993, 5494.487, 5496.5, 5496.47, 5494.001, 5486.876, 5486.742, 
    5466.065, 5460.943, 5448.104, 5434.286, 5423.547, 5416.651, 5413.329, 
    5412.42,
  5462.943, 5465.151, 5465.887, 5464.382, 5461.584, 5456.643, 5446.687, 
    5447.768, 5434.744, 5424.177, 5418.778, 5410.097, 5406.018, 5402.208, 
    5404.134,
  5435.491, 5435.121, 5434.202, 5432.761, 5429.422, 5426.254, 5422.308, 
    5413.446, 5411.658, 5411.032, 5406.631, 5404.245, 5402.791, 5402.388, 
    5404.124,
  5415.122, 5413.772, 5411.608, 5409.905, 5407.765, 5404.754, 5401.738, 
    5401.721, 5398.349, 5395.904, 5397.118, 5399.21, 5400.577, 5402.589, 
    5405.838,
  5399.136, 5396.449, 5393.905, 5392.296, 5389.432, 5387.38, 5384.115, 
    5380.59, 5381.032, 5384.655, 5388.631, 5392.22, 5397.647, 5401.716, 
    5405.266,
  5386.372, 5384.426, 5381.47, 5379.114, 5375.802, 5371.553, 5367.439, 
    5365.297, 5363.889, 5365.559, 5372.187, 5381.824, 5389.631, 5398.109, 
    5404.91,
  5376.821, 5373.534, 5370.443, 5367.324, 5362.021, 5356.101, 5349.257, 
    5343.043, 5341.004, 5345.299, 5354.217, 5367.491, 5381.288, 5393.539, 
    5403.577,
  5537.889, 5562.251, 5586.783, 5608.752, 5629.493, 5644.991, 5656.654, 
    5665.619, 5669.41, 5666.881, 5661.52, 5650.232, 5632.618, 5608.641, 
    5580.224,
  5519.409, 5542.928, 5566.01, 5587.895, 5605.727, 5622.166, 5635.156, 
    5640.416, 5644.254, 5646.331, 5638.183, 5626.166, 5606.908, 5585.479, 
    5555.832,
  5501.444, 5524.376, 5546.336, 5567.702, 5584.255, 5602.482, 5605.387, 
    5621.459, 5618.279, 5617.859, 5611.731, 5600.04, 5580.755, 5557.797, 
    5534.724,
  5482.505, 5501.556, 5521.534, 5539.731, 5558.22, 5568.178, 5587.995, 
    5582.09, 5593.098, 5590.561, 5583.873, 5571.163, 5555.407, 5536.93, 
    5518.732,
  5464.037, 5480.039, 5496.196, 5513.182, 5528.317, 5544.999, 5547.909, 
    5565.041, 5561.267, 5557.104, 5554.934, 5543.287, 5532.121, 5517.887, 
    5506.266,
  5448.034, 5458.889, 5471.199, 5486.098, 5498.685, 5510.439, 5522.217, 
    5521.818, 5527.405, 5530.215, 5524.67, 5518.865, 5511.965, 5503.841, 
    5497.089,
  5433.242, 5440.411, 5449.348, 5459.43, 5471.406, 5481.465, 5489.224, 
    5498.996, 5500.961, 5499.633, 5500.523, 5498.638, 5495.19, 5492.029, 
    5489.159,
  5416.73, 5421.277, 5427.31, 5435.22, 5443.214, 5452.368, 5460.388, 
    5465.668, 5472.149, 5478.528, 5480.103, 5481.091, 5481.966, 5482.605, 
    5484.518,
  5401.541, 5404.771, 5408.545, 5413.575, 5419.528, 5426.46, 5433.84, 
    5442.938, 5450.008, 5455.594, 5461.991, 5467.514, 5471.881, 5475.601, 
    5482.149,
  5389.282, 5390.084, 5391.823, 5395.414, 5399.274, 5404.575, 5410.768, 
    5417.829, 5427.073, 5438.26, 5447.945, 5456.827, 5465.672, 5473.183, 
    5483.969,
  5527.392, 5550.096, 5574.014, 5598.701, 5622.871, 5646.336, 5669.091, 
    5690.646, 5707.166, 5717.697, 5724.575, 5726.814, 5722.753, 5712.345, 
    5696.849,
  5510.066, 5533.08, 5556.267, 5580.498, 5603.711, 5627.641, 5651.551, 
    5670.118, 5687.008, 5702.733, 5709.37, 5712.413, 5708.062, 5700.399, 
    5683.761,
  5492.04, 5513.464, 5536.81, 5561.712, 5584.876, 5612.011, 5628.207, 
    5657.179, 5670.106, 5682.999, 5691.754, 5695.88, 5692.307, 5683.553, 
    5668.735,
  5474.625, 5492.076, 5514.979, 5538.622, 5564.362, 5584.244, 5616.086, 
    5624.02, 5649.461, 5663.672, 5673.063, 5676.699, 5675.828, 5667.29, 
    5652.696,
  5456.89, 5471.892, 5491.35, 5516.008, 5540.408, 5567.873, 5583.924, 
    5616.371, 5627.824, 5640.519, 5653.016, 5656.719, 5656.958, 5648.434, 
    5637.564,
  5440.808, 5452.138, 5468.13, 5490.195, 5514.267, 5539.455, 5567.602, 
    5582.11, 5603.168, 5624.054, 5630.663, 5637.971, 5638.661, 5633.361, 
    5621.518,
  5425.775, 5435.035, 5447.914, 5466.537, 5490.157, 5515.274, 5538.858, 
    5567.913, 5587.937, 5598.473, 5611.548, 5618.9, 5619.398, 5614.274, 
    5602.047,
  5411.417, 5419.083, 5429.473, 5444.479, 5464.208, 5489.527, 5515.048, 
    5535.213, 5556.976, 5577.721, 5589.46, 5596.025, 5599.055, 5594.744, 
    5585.717,
  5396.502, 5404.404, 5414.696, 5427.413, 5444.687, 5465.487, 5490.417, 
    5517.137, 5538.27, 5553.12, 5565.546, 5574.471, 5577.853, 5575.751, 
    5569.439,
  5383.057, 5389.123, 5398.747, 5411.802, 5426.792, 5446.968, 5468.769, 
    5490.066, 5510.794, 5529.835, 5544.158, 5553.583, 5558.411, 5558.188, 
    5555.864,
  5541.181, 5558.196, 5584.181, 5608.087, 5631.09, 5651.756, 5671.36, 
    5691.652, 5709.109, 5722.837, 5733.923, 5741.023, 5743.425, 5741.109, 
    5733.476,
  5529.958, 5544.889, 5564.712, 5590.523, 5613.532, 5634.869, 5655.896, 
    5672.926, 5690.394, 5708.2, 5719.337, 5727.184, 5730.492, 5729.97, 
    5723.448,
  5516.544, 5531.435, 5548, 5569.179, 5594.772, 5619.919, 5634.521, 5660.312, 
    5674.459, 5689.23, 5702.331, 5711.758, 5716.392, 5715.974, 5712.005,
  5501.123, 5515.326, 5530.17, 5547.18, 5569.687, 5590.881, 5620.911, 
    5630.126, 5654.799, 5671.159, 5684.922, 5694.622, 5701.403, 5702.43, 
    5698.918,
  5481.007, 5496.381, 5511.071, 5527.15, 5545.333, 5569.69, 5586.777, 
    5618.754, 5633.646, 5648.74, 5666.38, 5676.364, 5684.855, 5686.471, 
    5685.38,
  5457.808, 5472.163, 5487.232, 5504.177, 5519.728, 5539.755, 5564.437, 
    5582.201, 5605.936, 5629.595, 5643.654, 5657.696, 5666.374, 5670.724, 
    5670.457,
  5432.396, 5445.95, 5461.537, 5478.748, 5497.081, 5515.142, 5534.068, 
    5561.443, 5583.031, 5600.109, 5621.234, 5636.346, 5646.783, 5653.119, 
    5654.748,
  5405.854, 5418.119, 5432.024, 5449.437, 5467.014, 5487.382, 5507.39, 
    5526.255, 5548.999, 5575.257, 5595.712, 5612.209, 5626.037, 5634.548, 
    5639.146,
  5381.199, 5392.423, 5405.705, 5421.891, 5439.747, 5458.699, 5478.868, 
    5502.846, 5525.698, 5545.949, 5567.429, 5588.166, 5603.661, 5615.294, 
    5621.574,
  5358.048, 5368.957, 5381.127, 5395.143, 5410.828, 5429.622, 5449.747, 
    5470.439, 5494.052, 5519.32, 5542.419, 5562.86, 5580.797, 5595.359, 
    5603.769,
  5509.694, 5520.297, 5537.893, 5558.469, 5582.671, 5607.169, 5633.249, 
    5661.984, 5687.927, 5711.893, 5731.241, 5747.594, 5756.333, 5761.317, 
    5759.467,
  5512.596, 5525.945, 5542.604, 5561.885, 5581.826, 5605.808, 5630.747, 
    5656.003, 5679.848, 5706.207, 5724.787, 5739.925, 5749.014, 5754.388, 
    5753.614,
  5508.929, 5528.155, 5543.389, 5563.565, 5582.074, 5606.237, 5625.989, 
    5654.276, 5676.911, 5697.362, 5715.737, 5730.16, 5739.567, 5744.789, 
    5745.797,
  5501.242, 5521.682, 5539.205, 5557.081, 5578.912, 5594.53, 5624.56, 
    5639.009, 5664.837, 5686.787, 5704.277, 5717.617, 5727.978, 5733.636, 
    5735.425,
  5490.308, 5509.513, 5528.073, 5549.131, 5567.716, 5592.811, 5605.958, 
    5635.186, 5655.605, 5671.451, 5690.065, 5702.61, 5713.631, 5719.625, 
    5723.84,
  5476.699, 5492.876, 5511.367, 5531.396, 5552.695, 5571.933, 5597.376, 
    5611.437, 5633.432, 5655.995, 5670.965, 5685.963, 5696.63, 5704.291, 
    5708.992,
  5455.648, 5471.745, 5490.386, 5510.757, 5532.761, 5554.917, 5573.676, 
    5598.157, 5617.098, 5632.121, 5650.276, 5664.675, 5676.469, 5685.743, 
    5691.875,
  5429.038, 5444.765, 5462.686, 5483.785, 5504.547, 5527.481, 5549.777, 
    5567.293, 5585.914, 5607.588, 5624.893, 5639.553, 5652.927, 5663.329, 
    5671.168,
  5397.377, 5412.625, 5431.261, 5452.886, 5475.451, 5497.52, 5518.747, 
    5542.122, 5562.327, 5578.203, 5594.021, 5609.581, 5623.306, 5635.366, 
    5645.554,
  5363.188, 5377.875, 5396.352, 5417.268, 5439.202, 5462.576, 5484.222, 
    5504.086, 5523.956, 5544.335, 5561.943, 5576.873, 5590.675, 5603.486, 
    5614.688,
  5408.028, 5419.442, 5446.003, 5477.659, 5514.65, 5552.683, 5597.686, 
    5638.625, 5675.561, 5703.415, 5725.379, 5746.485, 5761.916, 5772.467, 
    5776.045,
  5411.137, 5420.767, 5445.417, 5477.868, 5511.896, 5551.624, 5593.919, 
    5631.834, 5665.537, 5698.242, 5722.015, 5742.607, 5759.643, 5772.018, 
    5777.113,
  5421.917, 5427.236, 5450.024, 5480.077, 5514.241, 5553.752, 5589.912, 
    5630.569, 5662.995, 5690.575, 5716.021, 5736.927, 5755.062, 5767.35, 
    5775.548,
  5433.847, 5437.218, 5456.779, 5481.948, 5516.816, 5544.103, 5591.43, 
    5615.563, 5651.09, 5682.58, 5709.109, 5729.818, 5748.682, 5762.132, 
    5771.006,
  5439.868, 5448.761, 5463.998, 5488.978, 5515.747, 5551.524, 5574.601, 
    5619.096, 5645.806, 5672.152, 5699.401, 5720.399, 5739.496, 5752.688, 
    5762.951,
  5440.914, 5453.403, 5469.386, 5491.637, 5517.186, 5541.967, 5577.207, 
    5599.94, 5628.933, 5663.683, 5685.991, 5709.888, 5727.255, 5742.289, 
    5752.356,
  5437.691, 5451.588, 5469.012, 5491.993, 5517.234, 5541.6, 5564.616, 
    5600.216, 5626.759, 5646.34, 5672.606, 5694.476, 5712.186, 5727.104, 
    5737.579,
  5429.852, 5443.745, 5460.39, 5483.959, 5507.943, 5533.263, 5557.566, 
    5577.703, 5602.523, 5632.395, 5656.204, 5676.137, 5694.626, 5709.125, 
    5720.563,
  5415.236, 5430.332, 5448.017, 5470.228, 5496.291, 5521.221, 5545.981, 
    5572.968, 5596.373, 5615.952, 5636.307, 5656.538, 5673.407, 5687.785, 
    5699.013,
  5397.384, 5410.092, 5428.725, 5450.337, 5474.186, 5502.118, 5527.446, 
    5549.447, 5571.657, 5595.394, 5616.254, 5634.802, 5650.968, 5665.247, 
    5676.419,
  5404.65, 5403.135, 5419.979, 5450.5, 5489.672, 5533.583, 5576.719, 
    5625.407, 5659.897, 5688.709, 5709.652, 5725.387, 5734.022, 5738.012, 
    5737.481,
  5406.057, 5407.406, 5422.15, 5452.005, 5488.996, 5532.574, 5576.658, 
    5623.18, 5655.694, 5690.769, 5714.301, 5732.509, 5743.137, 5751.069, 
    5753.121,
  5412.553, 5414.897, 5430.263, 5456.935, 5492.436, 5537.222, 5575.712, 
    5627.452, 5662.13, 5692.034, 5717.365, 5737.093, 5751.757, 5760.404, 
    5765.929,
  5419.683, 5423.277, 5439.359, 5461.266, 5496.098, 5527.093, 5582.402, 
    5616.008, 5656.245, 5691.343, 5719.606, 5739.688, 5757.065, 5767.821, 
    5776.326,
  5424.325, 5432.067, 5447.258, 5469.455, 5495.626, 5535.97, 5568.122, 
    5624.852, 5660.607, 5690.212, 5718.829, 5740.646, 5759.832, 5771.952, 
    5781.827,
  5428.276, 5436.341, 5452.966, 5472.618, 5497.04, 5527.063, 5572.395, 
    5608.159, 5646.229, 5688.525, 5714.897, 5739.683, 5758.176, 5773.825, 
    5783.824,
  5430.993, 5439.127, 5457.127, 5475.078, 5501.107, 5529.501, 5561.773, 
    5610.656, 5650.911, 5679.822, 5710.258, 5734.68, 5754.391, 5770.634, 
    5781.626,
  5429.673, 5439.189, 5455.014, 5474.701, 5497.096, 5525.79, 5555.95, 
    5590.56, 5627.926, 5669.342, 5701.035, 5725.693, 5747.07, 5763.964, 
    5776.479,
  5425.033, 5435.014, 5451.103, 5470.939, 5494.188, 5519.694, 5546.684, 
    5585.947, 5624.792, 5657.452, 5686.898, 5714.002, 5735.478, 5753.079, 
    5765.774,
  5417.957, 5426.553, 5442.476, 5461.519, 5482.801, 5509.432, 5535.228, 
    5564.243, 5599.817, 5637.387, 5670.22, 5697.847, 5720.287, 5738.356, 
    5751.433,
  5479.718, 5481.107, 5488.431, 5504.18, 5529.154, 5555.154, 5584.204, 
    5609.91, 5633.073, 5647.614, 5656.79, 5657.728, 5657.523, 5663.001, 
    5667.58,
  5465.314, 5462.721, 5463.733, 5478.108, 5501.983, 5533.909, 5570.214, 
    5599.594, 5624.052, 5646.159, 5657.919, 5662.224, 5665.564, 5673.874, 
    5679.915,
  5453.689, 5446.487, 5444.036, 5455.768, 5479.546, 5516.961, 5552.235, 
    5595.968, 5625.075, 5645.041, 5659.697, 5667.946, 5677.248, 5687.367, 
    5696.752,
  5444.784, 5434.116, 5429.521, 5436.65, 5462.075, 5493.674, 5546.424, 
    5578.739, 5616.211, 5643.372, 5662.942, 5674.95, 5689.932, 5703.103, 
    5713.485,
  5438.935, 5427.644, 5421.082, 5427.835, 5449.27, 5488.757, 5527.917, 
    5582.706, 5618.131, 5643.149, 5665.611, 5683.075, 5702.464, 5715.777, 
    5728.181,
  5436.272, 5426.208, 5418.317, 5424.889, 5444.428, 5478.907, 5530.178, 
    5569.25, 5608.033, 5645.468, 5668.402, 5691.584, 5711.317, 5727.913, 
    5739.963,
  5435.583, 5428.937, 5423.148, 5429.476, 5449.617, 5482.372, 5526.282, 
    5577.025, 5616.714, 5645.009, 5672.665, 5697.864, 5718.828, 5736.195, 
    5749.721,
  5436.776, 5434.271, 5429.913, 5437.867, 5455.665, 5487.989, 5530.926, 
    5569.875, 5607.125, 5645.813, 5674.979, 5701.549, 5723.835, 5742.274, 
    5757.529,
  5438.482, 5440.57, 5441.062, 5450.152, 5468.556, 5496.96, 5535.219, 
    5578.668, 5615.239, 5647.17, 5675.274, 5703.439, 5725.616, 5745.341, 
    5761.595,
  5441.221, 5444.859, 5448.723, 5459.921, 5476.8, 5504.863, 5538.565, 
    5573.746, 5607.497, 5643.789, 5673.902, 5701.696, 5724.543, 5745.139, 
    5762.324,
  5545.29, 5546.539, 5556.211, 5567.605, 5582.409, 5594.658, 5605.561, 
    5614.878, 5622.538, 5627.171, 5628.45, 5621.37, 5613.774, 5603.717, 
    5599.71,
  5530.135, 5528.733, 5531.978, 5545.73, 5560.468, 5579.433, 5595.292, 
    5605.585, 5615.816, 5625.171, 5628.579, 5625.264, 5619.879, 5613.956, 
    5612.302,
  5511.664, 5509.488, 5509.79, 5518.745, 5535.044, 5560.454, 5577.426, 
    5601.581, 5611.379, 5621.229, 5627.396, 5628.226, 5626.618, 5623.203, 
    5624.141,
  5493.101, 5488.391, 5488.142, 5491.744, 5506.279, 5525.759, 5561.383, 
    5579.466, 5603.035, 5616.663, 5626.403, 5630.091, 5633.612, 5633.148, 
    5638.432,
  5475.103, 5468.584, 5465.946, 5469.107, 5477.75, 5500.819, 5527.197, 
    5568.9, 5593.481, 5609.093, 5623.235, 5631.776, 5639.497, 5641.969, 
    5650.723,
  5458.706, 5452.196, 5448.202, 5449.185, 5454.858, 5470.183, 5503.19, 
    5537.273, 5573.283, 5602.904, 5618.149, 5633.047, 5643.578, 5651.88, 
    5662.021,
  5448.741, 5443.75, 5438.291, 5435.115, 5438.536, 5450.225, 5475.217, 
    5520.301, 5562.059, 5591.337, 5613.433, 5632.555, 5647.435, 5658.252, 
    5672.167,
  5444.053, 5438.005, 5428.434, 5422.489, 5419.775, 5431.422, 5454.365, 
    5493.233, 5540.838, 5581.603, 5607.995, 5631.153, 5650.772, 5664.667, 
    5681.969,
  5441.152, 5433.953, 5422.723, 5412.405, 5406.382, 5415.146, 5438.101, 
    5481.094, 5531.908, 5572.422, 5601.913, 5630.293, 5652.305, 5670.091, 
    5689.145,
  5440.277, 5430.946, 5419.586, 5406.917, 5396.005, 5403.396, 5427.391, 
    5465.472, 5516.88, 5564.132, 5597.576, 5628.915, 5653.962, 5675.017, 
    5696.373,
  5588.331, 5595.296, 5603.701, 5609.851, 5618.247, 5625.691, 5631.091, 
    5637.016, 5640.856, 5642.736, 5645.695, 5649.95, 5657.368, 5667.718, 
    5677.605,
  5573.541, 5580.96, 5589.277, 5597.749, 5606.213, 5614.849, 5624.781, 
    5631.167, 5637.325, 5644.799, 5649.392, 5655.947, 5664.484, 5678.406, 
    5690.374,
  5551.892, 5561.047, 5569.316, 5580.312, 5588.186, 5603.262, 5608.857, 
    5625.625, 5633.891, 5641.909, 5649.509, 5657.607, 5669.111, 5683.747, 
    5699.406,
  5532.219, 5535.888, 5543.946, 5552.398, 5566.219, 5574.464, 5596.56, 
    5602.916, 5621.265, 5634.426, 5646.473, 5655.185, 5668.792, 5686.111, 
    5704.951,
  5519.109, 5519.318, 5520.137, 5525.837, 5534.826, 5551.794, 5564.005, 
    5591.088, 5608.62, 5621.929, 5638.081, 5650.755, 5665.065, 5684.159, 
    5705.475,
  5504.312, 5502.191, 5500.796, 5503.777, 5507.587, 5518.257, 5536.57, 
    5555.218, 5579.542, 5607.327, 5626.543, 5643.267, 5658.073, 5679.944, 
    5703.349,
  5491.157, 5487.263, 5484.389, 5484.213, 5487.855, 5494.489, 5505.218, 
    5528.583, 5559.094, 5585.386, 5611.666, 5633.123, 5650.229, 5671.449, 
    5697.395,
  5478.543, 5472.021, 5467.444, 5467.493, 5468.701, 5473.976, 5483.063, 
    5496.056, 5522.776, 5561.188, 5592.836, 5620.362, 5640.892, 5662.103, 
    5689.627,
  5467.597, 5458.656, 5451.012, 5447.518, 5448.034, 5453.254, 5461.732, 
    5477.27, 5500.902, 5535.929, 5571.86, 5605.297, 5629.871, 5651.916, 
    5679.335,
  5459.104, 5445.741, 5436.412, 5432.373, 5429.586, 5431.49, 5439.973, 
    5452.312, 5474.295, 5511.124, 5550.888, 5589.096, 5617.957, 5641.862, 
    5669.23 ;
}
