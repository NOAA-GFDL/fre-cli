netcdf \00010101.atmos_daily.tile3.pr {
dimensions:
	time = UNLIMITED ; // (182 currently)
	phalf = 66 ;
	grid_xt = 15 ;
	grid_yt = 10 ;
	scalar_axis = 1 ;
	nv = 2 ;
	pfull = 65 ;
variables:
	double average_DT(time) ;
		average_DT:_FillValue = 1.e+20 ;
		average_DT:missing_value = 1.e+20 ;
		average_DT:units = "days" ;
		average_DT:long_name = "Length of average period" ;
	double average_T1(time) ;
		average_T1:_FillValue = 1.e+20 ;
		average_T1:missing_value = 1.e+20 ;
		average_T1:units = "days since 0001-01-01 00:00:00" ;
		average_T1:long_name = "Start time for average period" ;
	double average_T2(time) ;
		average_T2:_FillValue = 1.e+20 ;
		average_T2:missing_value = 1.e+20 ;
		average_T2:units = "days since 0001-01-01 00:00:00" ;
		average_T2:long_name = "End time for average period" ;
	float bk(phalf) ;
		bk:_FillValue = 1.e+20f ;
		bk:missing_value = 1.e+20f ;
		bk:long_name = "vertical coordinate sigma value" ;
		bk:cell_methods = "time: point" ;
	double grid_xt(grid_xt) ;
		grid_xt:units = "degrees_E" ;
		grid_xt:long_name = "T-cell longitude" ;
		grid_xt:axis = "X" ;
	double grid_yt(grid_yt) ;
		grid_yt:units = "degrees_N" ;
		grid_yt:long_name = "T-cell latitude" ;
		grid_yt:axis = "Y" ;
	float height10m(scalar_axis) ;
		height10m:_FillValue = 1.e+20f ;
		height10m:missing_value = 1.e+20f ;
		height10m:units = "m" ;
		height10m:long_name = "Height" ;
		height10m:cell_methods = "time: point" ;
		height10m:axis = "Z" ;
		height10m:positive = "up" ;
		height10m:standard_name = "height" ;
	float height2m(scalar_axis) ;
		height2m:_FillValue = 1.e+20f ;
		height2m:missing_value = 1.e+20f ;
		height2m:units = "m" ;
		height2m:long_name = "Height" ;
		height2m:cell_methods = "time: point" ;
		height2m:axis = "Z" ;
		height2m:positive = "up" ;
		height2m:standard_name = "height" ;
	double nv(nv) ;
		nv:long_name = "vertex number" ;
	double pfull(pfull) ;
		pfull:units = "mb" ;
		pfull:long_name = "ref full pressure level" ;
		pfull:axis = "Z" ;
		pfull:positive = "down" ;
	double phalf(phalf) ;
		phalf:units = "mb" ;
		phalf:long_name = "ref half pressure level" ;
		phalf:axis = "Z" ;
		phalf:positive = "down" ;
	float pk(phalf) ;
		pk:_FillValue = 1.e+20f ;
		pk:missing_value = 1.e+20f ;
		pk:units = "pascal" ;
		pk:long_name = "pressure part of the hybrid coordinate" ;
		pk:cell_methods = "time: point" ;
	float pr(time, grid_yt, grid_xt) ;
		pr:_FillValue = 1.e+20f ;
		pr:missing_value = 1.e+20f ;
		pr:units = "kg m-2 s-1" ;
		pr:long_name = "Precipitation" ;
		pr:cell_methods = "time: mean" ;
		pr:cell_measures = "area: area" ;
		pr:time_avg_info = "average_T1,average_T2,average_DT" ;
		pr:standard_name = "precipitation_flux" ;
		pr:interp_method = "conserve_order1" ;
	double scalar_axis(scalar_axis) ;
		scalar_axis:long_name = "none" ;
	double time(time) ;
		time:units = "days since 0001-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "NOLEAP" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bnds" ;
	double time_bnds(time, nv) ;
		time_bnds:long_name = "time axis boundaries" ;

// global attributes:
		:title = "cm5_c96_am5f7c1r0_b06_piC_galb_noiceinit_alb" ;
		:associated_files = "area: 00010101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:history = "Wed Apr 30 14:48:00 2025: ncks -d grid_xt,0,14 -d grid_yt,0,9 -d time,0,181 /home/cew/Code/cmip7-sprint/testfiles/input/00010101.atmos_daily.tile3.nc -O /home/cew/Code/cmip7-sprint/testfiles/00010101.atmos_daily.tile3.nc\nFri Apr 25 14:15:06 2025: ncks -x -v sphum,psl 00010101.atmos_daily.tile3.nc -o reduce/00010101.atmos_daily.tile3.nc\nFri Apr 25 13:47:12 2025: ncks -d grid_xt,35,55 -d grid_yt,30,45 00010101.atmos_daily.tile3.nc var_select/00010101.atmos_daily.tile3.nc" ;
		:NCO = "netCDF Operators version 5.1.9 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 average_DT = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 average_T1 = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 
    18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 
    36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 
    54, 55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 
    72, 73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 
    90, 91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 
    106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 
    120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 
    134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 
    148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 
    162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 
    176, 177, 178, 179, 180, 181 ;

 average_T2 = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 
    19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 
    37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 
    55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 
    73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 
    91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 106, 
    107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 
    121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 
    135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 
    149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 
    163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 
    177, 178, 179, 180, 181, 182 ;

 bk = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.00193294, 0.00749994, 0.01640714, 0.02841953, 
    0.04334756, 0.06103661, 0.0813586, 0.1042054, 0.1294836, 0.1571101, 
    0.1870091, 0.2191095, 0.2533426, 0.2896406, 0.3279357, 0.3681587, 
    0.4102391, 0.454293, 0.5001689, 0.5468886, 0.5935643, 0.6397641, 
    0.6851825, 0.729505, 0.7723162, 0.8125153, 0.8492141, 0.8817441, 
    0.909788, 0.9332725, 0.9524949, 0.9678352, 0.9798011, 0.9889621, 0.99575, 1 ;

 grid_xt = 36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50 ;

 grid_yt = 31, 32, 33, 34, 35, 36, 37, 38, 39, 40 ;

 height10m = 10 ;

 height2m = 2 ;


 nv = 1, 2 ;

 pfull = 0.0252729048206747, 0.0885404738757409, 0.213072411383256, 
    0.41190537807884, 0.671080828691593, 0.987471468515016, 1.36790961365676, 
    1.82562112064242, 2.38097588033244, 3.06218961364243, 3.90121721567151, 
    4.9296281825995, 6.18008131929323, 7.68875807563375, 9.49537809361575, 
    11.643153995098, 14.1786857151188, 17.1517875598959, 20.6152476986609, 
    24.6245259348741, 29.237386591333, 34.5134757786445, 40.5138467378254, 
    47.3004421634272, 54.9355325495126, 63.4811392623337, 72.9984371159701, 
    83.5471442618119, 95.1849171805989, 107.966767294215, 121.944503506415, 
    137.166169497631, 153.675572970355, 171.511834307961, 190.708985325578, 
    211.295632932361, 233.294677858721, 256.723099608772, 281.591803639405, 
    307.905555737256, 335.66293113824, 364.856338389786, 395.47216160598, 
    427.490864234311, 460.887168786725, 495.630391513078, 531.761718445649, 
    569.289185351388, 607.768705103107, 646.445374671436, 684.792067788697, 
    722.468679913451, 759.124006783627, 794.401045766566, 827.769968639223, 
    858.597822486016, 886.389109609622, 910.841030891388, 931.860653469283, 
    949.549679924174, 964.159924710431, 976.012345333387, 985.470174132691, 
    992.77226220014, 997.948601287575 ;

 phalf = 0.01, 0.0513470268, 0.1404240036, 0.3072783852, 0.5379505539, 
    0.8245489502, 1.170559845, 1.5862843323, 2.0879000854, 2.700272522, 
    3.4550848389, 4.3841940308, 5.5185266113, 6.8925054932, 8.5440936279, 
    10.5147802734, 12.8495031738, 15.5965148926, 18.8071691895, 
    22.5356542969, 26.8386547852, 31.7749560547, 37.4049951172, 
    43.7903613281, 50.9932617188, 59.0759326172, 68.100078125, 78.1262353516, 
    89.2131933594, 101.4173632812, 114.7922466406, 129.3878501562, 
    145.2501478125, 162.4206823438, 180.9360560938, 200.8276451562, 
    222.1212074219, 244.8367185938, 268.9881007812, 294.5831945312, 
    321.6236510156, 350.1049399219, 380.0163883594, 411.3414303125, 
    444.0575547656, 478.1367280469, 513.5456339062, 550.403556875, 
    588.6019571094, 627.3470909766, 665.9273852344, 704.0097012891, 
    741.2475327734, 777.2856108203, 811.7659041211, 843.9830114648, 
    873.3803854492, 899.5263707422, 922.2501762402, 941.5376650684, 
    957.6070185254, 970.7426572876, 981.30107, 989.65107, 995.9000099865, 1000 ;

 pk = 1, 5.134703, 14.0424, 30.72784, 53.79506, 82.4549, 117.056, 158.6284, 
    208.79, 270.0273, 345.5085, 438.4194, 551.8527, 689.2505, 854.4094, 
    1051.478, 1284.95, 1559.651, 1880.717, 2253.565, 2683.865, 3177.496, 
    3740.5, 4379.036, 5099.326, 5907.593, 6810.008, 7812.624, 8921.319, 
    10141.74, 11285.93, 12188.79, 12884.3, 13400.12, 13758.85, 13979.1, 
    14076.26, 14063.13, 13950.46, 13747.31, 13461.45, 13099.54, 12667.38, 
    12170.08, 11612.19, 10997.8, 10330.65, 9611.055, 8843.304, 8045.85, 
    7236.312, 6424.557, 5606.509, 4778.059, 3944.972, 3146.775, 2416.634, 
    1778.226, 1246.215, 826.5195, 511.2139, 290.7407, 150, 68.893, 14.999, 0 ;

 pr =
  1.541242e-05, 2.149244e-05, 1.789696e-05, 3.449073e-05, 2.898845e-05, 
    1.512394e-05, 1.853227e-05, 2.058743e-05, 1.964916e-05, 5.417909e-06, 
    6.469748e-06, 8.294474e-06, 4.556026e-06, 4.174302e-06, 8.112652e-07,
  3.304964e-05, 2.855557e-05, 2.48103e-05, 3.996154e-05, 2.033398e-05, 
    1.540473e-05, 2.119337e-05, 1.839629e-05, 2.010591e-05, 1.204061e-05, 
    9.248628e-06, 1.643999e-05, 1.432952e-05, 3.740712e-06, 6.340566e-07,
  2.534045e-05, 2.754723e-05, 3.171658e-05, 3.572768e-05, 2.471734e-05, 
    2.096064e-06, 1.998213e-05, 1.67057e-05, 1.929956e-05, 1.896231e-05, 
    1.636189e-05, 2.006903e-05, 2.098643e-05, 1.281043e-05, 5.704926e-06,
  3.098029e-05, 2.329577e-05, 2.966183e-05, 3.702644e-05, 3.815746e-05, 
    1.704895e-05, 2.312034e-06, 1.615273e-05, 2.379888e-05, 1.880619e-05, 
    1.717348e-05, 2.036215e-05, 2.227437e-05, 1.931813e-05, 1.215085e-05,
  5.019759e-05, 3.128999e-05, 3.013168e-05, 3.177963e-05, 3.684043e-05, 
    3.744761e-05, 2.050868e-05, 3.039537e-06, 6.722388e-06, 9.672612e-06, 
    1.475029e-05, 1.818954e-05, 2.200485e-05, 2.437644e-05, 1.912651e-05,
  5.403291e-05, 4.348331e-05, 3.468652e-05, 3.491564e-05, 3.3709e-05, 
    3.53848e-05, 3.447505e-05, 2.461184e-05, 1.636995e-05, 1.600544e-05, 
    1.260528e-05, 1.895299e-05, 2.190742e-05, 2.607091e-05, 2.208986e-05,
  5.01689e-05, 4.673811e-05, 3.903202e-05, 3.838182e-05, 3.828103e-05, 
    3.800392e-05, 3.834345e-05, 3.748023e-05, 3.334786e-05, 3.21458e-05, 
    2.53297e-05, 2.12881e-05, 2.228568e-05, 2.52427e-05, 2.482493e-05,
  5.790083e-05, 4.494716e-05, 3.954942e-05, 4.051331e-05, 3.755954e-05, 
    3.961224e-05, 4.153988e-05, 3.96587e-05, 3.895505e-05, 3.826829e-05, 
    3.429255e-05, 2.26958e-05, 2.379993e-05, 2.567318e-05, 2.399821e-05,
  4.721759e-05, 4.113105e-05, 3.815673e-05, 4.024105e-05, 3.708599e-05, 
    3.644662e-05, 3.709995e-05, 4.082697e-05, 4.040192e-05, 4.171166e-05, 
    3.637889e-05, 2.57895e-05, 2.530864e-05, 2.473353e-05, 1.735654e-05,
  3.364938e-05, 3.401121e-05, 3.603425e-05, 3.531952e-05, 3.373628e-05, 
    3.501731e-05, 3.616545e-05, 3.476049e-05, 2.928733e-05, 1.872777e-05, 
    2.544651e-05, 2.473375e-05, 2.280703e-05, 2.2938e-05, 1.901704e-05,
  1.76077e-05, 2.864065e-05, 1.776834e-05, 3.148875e-05, 1.508937e-05, 
    7.106938e-06, 2.181913e-05, 2.782342e-05, 3.137803e-05, 3.520778e-05, 
    4.732734e-05, 6.401946e-05, 5.233364e-05, 2.89776e-05, 2.358943e-05,
  4.307582e-05, 4.057435e-05, 4.180562e-05, 2.543804e-05, 5.837779e-06, 
    3.058517e-06, 2.23636e-05, 2.730484e-05, 2.95197e-05, 3.580458e-05, 
    4.368949e-05, 6.172113e-05, 5.117038e-05, 2.675562e-05, 1.987387e-05,
  5.131335e-05, 5.417901e-05, 5.288439e-05, 4.300658e-05, 1.343086e-05, 
    3.457004e-07, 1.25697e-05, 2.788672e-05, 3.400298e-05, 3.627205e-05, 
    4.337105e-05, 5.520205e-05, 4.9348e-05, 2.86029e-05, 1.637547e-05,
  4.812831e-05, 5.133654e-05, 5.419298e-05, 5.286975e-05, 4.325551e-05, 
    1.41237e-05, 1.120472e-06, 1.395564e-05, 2.853648e-05, 3.594159e-05, 
    4.130859e-05, 4.7857e-05, 4.391781e-05, 3.278372e-05, 1.785635e-05,
  4.53042e-05, 5.034003e-05, 4.927324e-05, 4.875718e-05, 4.662075e-05, 
    4.112302e-05, 1.465915e-05, 1.945829e-06, 1.149936e-05, 2.568054e-05, 
    3.628296e-05, 4.258106e-05, 3.871245e-05, 2.953047e-05, 1.993626e-05,
  4.317964e-05, 4.63599e-05, 4.774864e-05, 4.832307e-05, 4.654443e-05, 
    4.591968e-05, 4.397864e-05, 3.67497e-05, 2.601861e-05, 2.856782e-05, 
    2.572462e-05, 3.661433e-05, 3.543294e-05, 2.57325e-05, 1.911987e-05,
  4.269351e-05, 4.499312e-05, 4.432832e-05, 4.543574e-05, 4.369643e-05, 
    4.319287e-05, 4.12421e-05, 3.823872e-05, 4.36662e-05, 4.025041e-05, 
    3.021921e-05, 3.083509e-05, 3.223219e-05, 2.487799e-05, 1.796996e-05,
  4.032556e-05, 4.450034e-05, 4.252103e-05, 4.576749e-05, 4.338922e-05, 
    4.022404e-05, 3.970858e-05, 3.855252e-05, 4.279742e-05, 4.217462e-05, 
    2.867606e-05, 2.352637e-05, 2.6028e-05, 2.34745e-05, 1.773227e-05,
  3.680445e-05, 3.8561e-05, 3.932453e-05, 4.008911e-05, 4.10592e-05, 
    4.242024e-05, 4.183842e-05, 4.25545e-05, 4.257812e-05, 4.113019e-05, 
    2.809104e-05, 1.796148e-05, 1.856431e-05, 1.771724e-05, 1.29635e-05,
  2.843303e-05, 3.07888e-05, 3.418518e-05, 3.619152e-05, 3.659911e-05, 
    3.608476e-05, 3.940264e-05, 4.082692e-05, 3.383959e-05, 2.009884e-05, 
    2.079521e-05, 1.416753e-05, 1.292397e-05, 1.170525e-05, 8.398287e-06,
  7.106108e-06, 3.670168e-05, 2.88846e-05, 2.202875e-05, 5.372665e-06, 
    1.350819e-06, 7.190079e-06, 1.132825e-05, 6.466976e-06, 3.321941e-06, 
    4.574737e-06, 5.205121e-06, 2.596597e-06, 2.163669e-06, 1.301985e-06,
  4.009838e-05, 3.509641e-05, 3.697587e-05, 2.820417e-05, 6.392709e-06, 
    6.295394e-07, 1.232776e-05, 1.453577e-05, 6.511846e-06, 7.562039e-06, 
    6.278542e-06, 1.045935e-05, 9.465883e-06, 1.30805e-06, 6.833992e-07,
  3.503971e-05, 3.417911e-05, 3.774076e-05, 3.748374e-05, 1.579207e-05, 
    1.184036e-06, 5.742508e-06, 1.46137e-05, 1.241755e-05, 1.337688e-05, 
    1.188243e-05, 1.271275e-05, 1.296508e-05, 4.735341e-06, 5.874992e-07,
  3.529558e-05, 3.386871e-05, 3.967529e-05, 4.145858e-05, 4.401032e-05, 
    1.389758e-05, 2.564483e-06, 8.944627e-06, 1.747162e-05, 1.942495e-05, 
    1.542892e-05, 1.26918e-05, 1.172026e-05, 8.336124e-06, 1.337085e-06,
  3.723596e-05, 3.666956e-05, 3.789528e-05, 4.137732e-05, 4.707062e-05, 
    4.249486e-05, 7.523884e-06, 2.050615e-06, 5.395336e-06, 1.15063e-05, 
    1.527645e-05, 1.421404e-05, 1.145178e-05, 7.691116e-06, 2.805901e-06,
  3.648175e-05, 3.707033e-05, 3.878397e-05, 4.180503e-05, 4.775535e-05, 
    4.881659e-05, 3.888029e-05, 2.997961e-05, 1.846556e-05, 2.206802e-05, 
    1.332975e-05, 1.529024e-05, 1.224978e-05, 6.190134e-06, 2.958833e-06,
  3.925908e-05, 4.129323e-05, 4.056869e-05, 4.317392e-05, 4.581196e-05, 
    4.981386e-05, 4.843214e-05, 4.989196e-05, 4.048089e-05, 3.314703e-05, 
    2.424715e-05, 1.76877e-05, 1.319223e-05, 6.311184e-06, 2.774854e-06,
  4.088867e-05, 4.21737e-05, 4.627809e-05, 4.676771e-05, 4.444002e-05, 
    4.957293e-05, 4.8714e-05, 5.927267e-05, 5.232033e-05, 4.109531e-05, 
    3.365188e-05, 2.267609e-05, 1.833405e-05, 7.386638e-06, 3.835118e-06,
  3.886756e-05, 4.237497e-05, 4.564897e-05, 4.671698e-05, 4.964941e-05, 
    4.870181e-05, 4.883225e-05, 5.750599e-05, 5.689275e-05, 4.763461e-05, 
    3.870661e-05, 2.895994e-05, 2.243406e-05, 1.501851e-05, 7.439327e-06,
  3.417029e-05, 4.132056e-05, 4.452689e-05, 4.569264e-05, 4.866045e-05, 
    5.059425e-05, 5.060138e-05, 5.159399e-05, 4.085731e-05, 3.639381e-05, 
    3.66254e-05, 2.962897e-05, 2.69435e-05, 2.110098e-05, 9.786656e-06,
  1.412738e-05, 3.444016e-05, 1.635069e-05, 2.225159e-05, 7.356462e-06, 
    8.719302e-07, 2.014427e-06, 3.486881e-06, 3.841482e-06, 2.111431e-06, 
    7.175692e-07, 9.108653e-07, 5.561317e-07, 1.272681e-07, 2.690871e-07,
  3.631439e-05, 3.37885e-05, 2.48995e-05, 1.747194e-05, 6.427564e-06, 
    2.510525e-07, 2.213334e-06, 3.22136e-06, 4.88044e-06, 3.200353e-06, 
    1.247699e-06, 2.836145e-06, 3.682734e-06, 3.42205e-08, 2.658369e-07,
  3.351846e-05, 2.381559e-05, 1.586314e-05, 1.812548e-05, 1.985387e-05, 
    7.334171e-07, 4.118428e-06, 7.266663e-06, 8.08518e-06, 7.848668e-06, 
    3.929903e-06, 3.392017e-06, 5.330818e-06, 3.87821e-06, 8.943454e-07,
  2.953811e-05, 1.496253e-05, 1.609937e-05, 1.831245e-05, 1.645817e-05, 
    5.183783e-06, 4.002048e-06, 5.362692e-06, 9.015164e-06, 9.118558e-06, 
    5.044044e-06, 4.002778e-06, 4.895315e-06, 5.037329e-06, 3.294717e-06,
  2.186925e-05, 1.425226e-05, 1.705011e-05, 1.835076e-05, 1.859686e-05, 
    2.50432e-05, 5.595197e-06, 2.7204e-06, 9.917804e-06, 3.8406e-06, 
    4.141937e-06, 4.583349e-06, 4.039588e-06, 3.886976e-06, 4.157724e-06,
  1.979912e-05, 1.518336e-05, 1.828795e-05, 1.711965e-05, 1.453967e-05, 
    2.846233e-05, 3.653477e-05, 1.00077e-05, 6.513677e-06, 1.137004e-05, 
    5.253334e-06, 4.09401e-06, 5.057036e-06, 3.682434e-06, 3.60486e-06,
  1.880611e-05, 1.776303e-05, 2.077824e-05, 1.521339e-05, 1.3767e-05, 
    2.771851e-05, 5.454841e-05, 3.307261e-05, 1.870485e-05, 1.397699e-05, 
    8.859436e-06, 5.220707e-06, 5.089776e-06, 4.91151e-06, 3.609422e-06,
  1.919027e-05, 2.068648e-05, 2.025739e-05, 1.960491e-05, 2.162403e-05, 
    3.15303e-05, 4.929882e-05, 3.467216e-05, 3.201815e-05, 2.176693e-05, 
    1.196053e-05, 5.668135e-06, 4.68384e-06, 5.203618e-06, 3.816795e-06,
  2.018142e-05, 2.152686e-05, 2.57855e-05, 2.41367e-05, 3.20894e-05, 
    3.495532e-05, 5.013483e-05, 3.623669e-05, 3.930576e-05, 1.867432e-05, 
    1.438282e-05, 6.87781e-06, 5.442775e-06, 5.600813e-06, 2.671478e-06,
  2.019565e-05, 2.283523e-05, 2.839691e-05, 3.400622e-05, 3.5409e-05, 
    3.545139e-05, 4.125768e-05, 3.571088e-05, 3.149284e-05, 2.456321e-05, 
    1.221603e-05, 7.44139e-06, 7.482104e-06, 5.503097e-06, 5.564933e-06,
  1.752341e-05, 2.099896e-05, 1.537613e-05, 2.173466e-05, 1.152757e-05, 
    4.971685e-06, 8.514819e-06, 3.574243e-06, 4.631477e-06, 2.614068e-06, 
    5.756787e-09, 1.016617e-06, 1.46572e-07, 7.788366e-08, 4.55008e-07,
  3.061757e-05, 2.768067e-05, 3.024626e-05, 3.695185e-05, 8.30832e-06, 
    5.380177e-06, 3.86527e-06, 3.439745e-06, 3.274955e-06, 3.304777e-06, 
    1.389057e-06, 2.84804e-06, 3.301066e-06, 4.41918e-07, 4.752208e-07,
  3.105542e-05, 2.622523e-05, 3.109545e-05, 4.069283e-05, 8.007421e-06, 
    6.22273e-06, 4.159048e-06, 5.101505e-06, 5.051807e-06, 4.263374e-06, 
    3.349738e-06, 2.779153e-06, 3.054392e-06, 2.109542e-06, 8.564373e-07,
  3.300374e-05, 2.806824e-05, 3.036661e-05, 3.879301e-05, 1.479754e-05, 
    7.166243e-07, 2.507696e-06, 5.116882e-06, 5.82435e-06, 4.166865e-06, 
    4.020592e-06, 2.532243e-06, 2.008002e-06, 1.417135e-06, 1.42629e-06,
  2.952376e-05, 3.114973e-05, 2.870732e-05, 4.113417e-05, 3.194893e-05, 
    6.580437e-06, 3.053424e-06, 1.463493e-07, 4.589897e-07, 2.77236e-07, 
    2.504381e-06, 2.519391e-06, 1.699709e-06, 1.717649e-06, 8.326155e-07,
  3.040198e-05, 3.231596e-05, 2.802285e-05, 3.641824e-05, 3.444136e-05, 
    2.795694e-05, 1.914651e-05, 2.357668e-06, 1.994413e-06, 7.307915e-06, 
    2.920713e-06, 2.248071e-06, 1.920849e-06, 1.234466e-06, 6.787951e-07,
  3.705618e-05, 3.34023e-05, 2.648386e-05, 3.159286e-05, 2.955497e-05, 
    3.914058e-05, 4.522553e-05, 2.220027e-05, 1.431991e-05, 1.110772e-05, 
    7.127015e-06, 2.768784e-06, 1.492566e-06, 1.24927e-06, 1.350831e-06,
  4.43046e-05, 3.436562e-05, 2.547515e-05, 2.70438e-05, 2.904631e-05, 
    3.622569e-05, 5.217173e-05, 3.874659e-05, 2.584917e-05, 2.092771e-05, 
    7.549831e-06, 2.63617e-06, 1.563876e-06, 1.645815e-06, 1.122549e-06,
  4.909705e-05, 3.40258e-05, 2.259159e-05, 2.231401e-05, 3.134281e-05, 
    3.785728e-05, 4.238695e-05, 3.91304e-05, 3.061182e-05, 2.232408e-05, 
    8.190901e-06, 2.533904e-06, 1.856204e-06, 2.396991e-06, 3.132101e-06,
  3.687808e-05, 1.86409e-05, 1.733961e-05, 2.4629e-05, 3.290036e-05, 
    3.397434e-05, 4.087497e-05, 3.626336e-05, 3.247584e-05, 1.804245e-05, 
    6.740474e-06, 2.608029e-06, 2.544454e-06, 3.917464e-06, 6.270015e-06,
  1.06478e-05, 1.431573e-05, 1.048107e-05, 1.287163e-05, 8.986055e-06, 
    3.892292e-06, 5.378562e-06, 5.099647e-06, 3.920752e-06, 1.090905e-06, 
    3.419457e-08, 4.124352e-07, 7.587582e-07, 6.906409e-07, 8.059101e-07,
  2.322648e-05, 2.387119e-05, 2.105791e-05, 2.240594e-05, 7.293786e-06, 
    4.666224e-06, 1.010588e-05, 5.663745e-06, 2.341855e-06, 1.705447e-06, 
    1.930042e-07, 1.168953e-06, 2.023119e-06, 8.371455e-07, 9.026458e-07,
  2.722425e-05, 2.825668e-05, 2.752863e-05, 3.183777e-05, 1.555354e-05, 
    4.297801e-06, 6.535015e-06, 4.288318e-06, 2.284601e-06, 1.688399e-06, 
    1.023505e-06, 9.42911e-07, 2.250051e-06, 2.393114e-06, 1.134731e-06,
  2.423591e-05, 2.654565e-05, 2.616609e-05, 3.669896e-05, 3.767787e-05, 
    6.328013e-06, 4.746244e-07, 2.228652e-06, 2.463529e-06, 1.141557e-06, 
    7.768962e-07, 4.356372e-07, 1.210966e-06, 1.795753e-06, 1.612568e-06,
  2.541812e-05, 2.563124e-05, 2.424826e-05, 3.129381e-05, 5.206249e-05, 
    2.070494e-05, 4.979934e-06, 3.150046e-07, 9.220792e-08, 2.429744e-08, 
    4.534852e-07, 2.158743e-07, 2.189301e-07, 1.826514e-06, 1.97209e-06,
  2.623544e-05, 2.377849e-05, 2.629076e-05, 3.276596e-05, 5.077579e-05, 
    3.031946e-05, 1.871367e-05, 4.494448e-06, 8.86356e-07, 2.825796e-06, 
    6.070585e-07, 2.16035e-07, 1.053637e-06, 2.217998e-06, 2.640924e-06,
  2.611388e-05, 2.659559e-05, 2.698322e-05, 3.540641e-05, 4.149429e-05, 
    3.658383e-05, 2.976739e-05, 2.127413e-05, 6.560479e-06, 7.505824e-06, 
    3.391236e-06, 4.457638e-07, 1.212298e-06, 2.147879e-06, 3.505626e-06,
  2.536511e-05, 2.712699e-05, 2.609855e-05, 3.842176e-05, 4.020065e-05, 
    3.068848e-05, 3.327176e-05, 3.605329e-05, 1.481386e-05, 1.677567e-05, 
    4.358502e-06, 6.029626e-07, 8.503265e-07, 3.121112e-06, 4.146217e-06,
  2.986007e-05, 2.917002e-05, 2.750625e-05, 4.146071e-05, 3.331664e-05, 
    2.649478e-05, 3.601538e-05, 3.18672e-05, 2.210747e-05, 2.143873e-05, 
    4.501671e-06, 6.521493e-07, 1.623643e-06, 3.246793e-06, 5.409243e-06,
  2.728973e-05, 2.489198e-05, 2.680654e-05, 3.519013e-05, 2.789481e-05, 
    2.304223e-05, 3.286481e-05, 3.442131e-05, 3.024768e-05, 1.269489e-05, 
    3.570869e-06, 9.656679e-07, 1.508252e-06, 2.905624e-06, 7.819478e-06,
  4.998793e-06, 7.65902e-06, 3.412169e-06, 5.245841e-06, 1.887118e-06, 
    3.041168e-06, 2.700231e-06, 1.53128e-06, 2.201577e-06, 1.532195e-06, 
    2.772602e-06, 2.358015e-06, 1.968987e-06, 1.393593e-06, 1.307008e-06,
  1.048298e-05, 1.494318e-05, 8.433472e-06, 1.12313e-05, 3.928435e-06, 
    2.583957e-06, 3.48558e-06, 1.506647e-06, 1.299753e-06, 1.85045e-06, 
    1.890599e-06, 3.966035e-06, 2.525848e-06, 1.577959e-06, 1.676463e-06,
  1.574986e-05, 1.802609e-05, 1.966399e-05, 1.5598e-05, 7.55392e-06, 
    2.757856e-06, 2.666781e-06, 1.407077e-06, 1.142679e-06, 2.308755e-06, 
    3.943802e-06, 5.13705e-06, 4.847727e-06, 3.3568e-06, 2.285886e-06,
  2.000883e-05, 2.696049e-05, 2.660057e-05, 2.720395e-05, 1.49541e-05, 
    7.735958e-06, 1.541842e-06, 6.129939e-08, 2.055062e-07, 1.060487e-06, 
    3.512821e-06, 3.0753e-06, 4.193606e-06, 3.231095e-06, 2.976665e-06,
  3.209926e-05, 3.366826e-05, 3.286461e-05, 3.452356e-05, 2.742427e-05, 
    1.319695e-05, 8.371133e-06, 2.66236e-06, 1.021162e-07, 8.98469e-07, 
    2.482654e-06, 3.033358e-06, 2.114281e-06, 4.35885e-06, 2.454068e-06,
  4.051539e-05, 3.744676e-05, 3.468842e-05, 3.213275e-05, 2.28083e-05, 
    2.252959e-05, 1.985927e-05, 3.177517e-06, 3.540291e-07, 1.222648e-06, 
    1.473193e-06, 2.277684e-06, 5.624359e-06, 5.522311e-06, 3.157246e-06,
  4.382286e-05, 4.7232e-05, 4.083032e-05, 3.308685e-05, 2.111509e-05, 
    2.485146e-05, 2.244575e-05, 1.488162e-05, 4.853005e-06, 2.868445e-06, 
    3.056387e-06, 2.302619e-06, 5.624697e-06, 5.441173e-06, 4.637694e-06,
  4.151858e-05, 4.808913e-05, 4.182328e-05, 3.613642e-05, 2.255305e-05, 
    2.105529e-05, 2.2509e-05, 1.880564e-05, 1.032971e-05, 9.882336e-06, 
    2.043281e-06, 1.114972e-06, 4.888148e-06, 6.157805e-06, 4.842219e-06,
  3.775155e-05, 4.475031e-05, 4.698021e-05, 3.4487e-05, 2.676021e-05, 
    1.937849e-05, 2.003453e-05, 1.896481e-05, 1.745352e-05, 9.744554e-06, 
    9.523638e-07, 5.158356e-07, 3.645368e-06, 6.140134e-06, 7.993112e-06,
  3.182033e-05, 3.316294e-05, 3.472876e-05, 3.111656e-05, 2.43347e-05, 
    1.740456e-05, 1.843311e-05, 2.499783e-05, 1.114864e-05, 1.293708e-06, 
    1.353442e-06, 2.360391e-07, 2.384027e-06, 5.382725e-06, 6.969449e-06,
  2.201507e-05, 1.809655e-05, 6.276631e-06, 4.392483e-06, 1.773554e-06, 
    3.522572e-07, 2.985092e-06, 3.576798e-06, 3.250454e-06, 1.637118e-06, 
    6.088225e-07, 5.360899e-07, 3.553882e-07, 3.413656e-07, 3.519811e-07,
  3.060243e-05, 2.574447e-05, 8.256703e-06, 7.890771e-06, 4.376517e-07, 
    2.342886e-07, 2.353646e-06, 3.394885e-06, 3.146197e-06, 3.260209e-06, 
    9.100903e-07, 6.487885e-07, 6.094171e-07, 2.671719e-07, 3.834202e-07,
  4.093137e-05, 3.442397e-05, 2.035385e-05, 1.302207e-05, 8.551165e-06, 
    1.589394e-06, 4.515638e-07, 2.731658e-06, 3.210897e-06, 3.269002e-06, 
    2.351889e-06, 9.835214e-07, 9.463446e-07, 8.064054e-07, 4.170828e-07,
  5.214785e-05, 5.47898e-05, 2.735289e-05, 1.727798e-05, 9.651163e-06, 
    5.410365e-06, 9.002266e-07, 1.128709e-06, 3.122523e-06, 3.695787e-06, 
    2.372291e-06, 2.122253e-06, 1.566494e-06, 1.36032e-06, 1.479317e-06,
  5.418365e-05, 5.748347e-05, 4.547316e-05, 3.379874e-05, 1.807458e-05, 
    1.40257e-05, 3.988113e-06, 1.506978e-06, 1.02718e-06, 2.171234e-06, 
    1.89155e-06, 2.688308e-06, 1.763245e-06, 1.491348e-06, 1.757153e-06,
  3.756225e-05, 4.828137e-05, 4.496732e-05, 2.878976e-05, 2.324308e-05, 
    1.919061e-05, 1.539657e-05, 3.142015e-06, 3.77586e-06, 6.24622e-06, 
    1.4737e-06, 3.344171e-06, 2.063058e-06, 1.89221e-06, 1.441565e-06,
  2.610262e-05, 3.746607e-05, 3.324546e-05, 2.733076e-05, 2.37115e-05, 
    1.929271e-05, 1.602088e-05, 1.237449e-05, 1.2518e-05, 1.268021e-05, 
    7.825873e-06, 4.13014e-06, 2.702758e-06, 2.788162e-06, 1.222801e-06,
  2.029222e-05, 2.43429e-05, 3.141717e-05, 2.648073e-05, 2.091228e-05, 
    1.893462e-05, 1.608677e-05, 1.236809e-05, 1.574148e-05, 1.338636e-05, 
    5.001908e-06, 4.503632e-06, 3.543877e-06, 3.268252e-06, 1.967328e-06,
  8.996947e-06, 2.023147e-05, 2.726487e-05, 2.325203e-05, 2.016671e-05, 
    2.030799e-05, 1.67495e-05, 1.475029e-05, 1.595659e-05, 1.249616e-05, 
    3.418822e-06, 4.661791e-06, 4.598432e-06, 4.292406e-06, 4.844431e-06,
  2.144176e-05, 1.019784e-05, 1.625401e-05, 2.199205e-05, 2.184052e-05, 
    1.500472e-05, 1.59726e-05, 1.647582e-05, 1.311972e-05, 6.501938e-06, 
    4.372801e-06, 4.185934e-06, 5.550366e-06, 5.267158e-06, 6.328429e-06,
  1.552007e-05, 3.279196e-05, 1.370485e-05, 8.230774e-06, 2.403046e-06, 
    8.947109e-07, 1.663719e-06, 8.984823e-07, 1.229593e-06, 1.472535e-07, 
    3.174239e-07, 2.630269e-07, 5.619775e-07, 2.567926e-07, 7.792533e-07,
  2.421359e-05, 3.86815e-05, 2.454916e-05, 1.695308e-05, 1.341209e-06, 
    1.254033e-06, 2.704043e-06, 1.537179e-06, 7.978408e-07, 4.93708e-07, 
    1.059226e-07, 2.118677e-07, 6.316327e-07, 3.901215e-07, 1.216401e-06,
  2.741767e-05, 4.107391e-05, 3.547553e-05, 2.119417e-05, 8.721006e-06, 
    1.180394e-06, 2.486973e-06, 1.630487e-06, 1.247308e-06, 8.813684e-07, 
    3.092141e-07, 4.067542e-07, 8.323493e-07, 2.190784e-06, 7.534626e-07,
  2.744207e-05, 4.211738e-05, 4.095511e-05, 2.377037e-05, 1.835674e-05, 
    5.369346e-06, 1.370283e-06, 3.709432e-07, 1.667814e-06, 6.972698e-07, 
    5.018362e-07, 2.880515e-07, 5.973994e-07, 1.463312e-06, 9.065301e-07,
  2.284937e-05, 3.670134e-05, 4.997773e-05, 4.136192e-05, 2.322079e-05, 
    1.769195e-05, 7.016017e-06, 2.258523e-06, 4.250411e-07, 4.471919e-08, 
    3.521147e-08, 2.757708e-07, 3.592066e-07, 7.00389e-07, 1.468963e-06,
  2.335516e-05, 3.570079e-05, 4.022707e-05, 3.551592e-05, 2.828414e-05, 
    2.462839e-05, 1.969481e-05, 4.573005e-06, 8.507042e-07, 1.222012e-06, 
    4.956352e-07, 7.572601e-07, 4.662857e-07, 6.920789e-07, 1.485584e-06,
  2.261596e-05, 3.085616e-05, 3.557306e-05, 2.797346e-05, 2.644337e-05, 
    2.269312e-05, 2.088257e-05, 1.707859e-05, 1.13213e-05, 4.805464e-06, 
    2.944914e-06, 7.601024e-07, 4.24443e-07, 8.518285e-07, 1.064457e-06,
  1.988127e-05, 2.709284e-05, 2.639515e-05, 2.546435e-05, 2.357973e-05, 
    2.106262e-05, 1.666488e-05, 1.682527e-05, 1.765642e-05, 1.282993e-05, 
    1.899801e-06, 1.1608e-06, 7.788253e-07, 5.764144e-07, 1.000481e-06,
  1.376657e-05, 2.070619e-05, 2.594516e-05, 1.944798e-05, 1.980348e-05, 
    1.977199e-05, 1.586107e-05, 1.47847e-05, 1.512546e-05, 1.247751e-05, 
    8.04066e-07, 1.315696e-06, 1.701364e-06, 1.089701e-06, 1.391836e-06,
  3.671504e-06, 1.172106e-05, 1.630736e-05, 1.800432e-05, 1.712807e-05, 
    1.66588e-05, 1.598885e-05, 1.19165e-05, 1.022398e-05, 1.910326e-06, 
    4.367544e-06, 3.755144e-06, 2.373468e-06, 2.344985e-06, 2.321552e-06,
  6.763263e-06, 1.193236e-05, 4.016117e-06, 5.889353e-06, 2.006802e-06, 
    1.824046e-07, 1.653464e-06, 1.690532e-06, 2.986036e-06, 1.192861e-06, 
    2.274012e-06, 2.820745e-06, 3.623316e-06, 2.152836e-06, 2.280014e-06,
  1.507645e-05, 1.987646e-05, 1.448813e-05, 1.055448e-05, 6.766785e-07, 
    3.750407e-08, 1.038627e-06, 1.217686e-06, 1.708718e-06, 1.056225e-06, 
    1.646769e-06, 1.809791e-06, 3.045232e-06, 3.113802e-06, 4.344904e-06,
  2.854803e-05, 2.438236e-05, 2.519524e-05, 1.568382e-05, 7.015562e-06, 
    7.744748e-07, 3.287183e-07, 6.237069e-07, 6.195275e-07, 8.705326e-07, 
    8.790709e-07, 1.731053e-06, 3.850345e-06, 8.319124e-06, 6.266853e-06,
  2.974493e-05, 2.911567e-05, 2.081978e-05, 2.096066e-05, 1.544463e-05, 
    5.639313e-06, 1.076971e-06, 5.464229e-08, 1.409378e-07, 4.800496e-07, 
    6.21204e-07, 1.140652e-06, 2.09036e-06, 3.95188e-06, 5.831717e-06,
  2.417445e-05, 2.594568e-05, 3.245455e-05, 2.746467e-05, 1.945025e-05, 
    1.164788e-05, 7.303208e-06, 1.635235e-06, 1.241921e-06, 4.352215e-07, 
    2.099072e-07, 7.629641e-07, 2.811809e-06, 3.222392e-06, 5.185057e-06,
  2.326039e-05, 2.246878e-05, 2.423201e-05, 2.413371e-05, 2.001474e-05, 
    1.708748e-05, 1.441458e-05, 7.062131e-06, 3.527574e-07, 5.240665e-08, 
    5.170422e-08, 4.927804e-07, 2.434387e-06, 3.86817e-06, 4.873932e-06,
  2.139024e-05, 2.055767e-05, 2.072162e-05, 1.950318e-05, 1.982272e-05, 
    1.549715e-05, 1.57318e-05, 1.518067e-05, 9.437919e-06, 4.229087e-06, 
    2.046076e-06, 1.040996e-06, 2.193831e-06, 3.765578e-06, 4.774584e-06,
  1.69181e-05, 1.869241e-05, 1.911675e-05, 2.028047e-05, 2.037645e-05, 
    1.756121e-05, 1.538677e-05, 1.662589e-05, 1.082312e-05, 7.717204e-06, 
    1.214045e-06, 7.056334e-07, 1.491254e-06, 3.159153e-06, 5.621006e-06,
  9.246479e-06, 1.707221e-05, 2.131385e-05, 1.804964e-05, 1.809993e-05, 
    1.867384e-05, 1.666229e-05, 1.303839e-05, 1.443538e-05, 6.680256e-06, 
    1.866727e-07, 1.458878e-06, 1.334596e-06, 2.027285e-06, 3.585908e-06,
  9.913512e-06, 1.039814e-05, 1.431267e-05, 1.641205e-05, 1.797968e-05, 
    1.775134e-05, 1.67597e-05, 1.452126e-05, 7.855944e-06, 3.512758e-07, 
    1.781435e-06, 9.459179e-07, 5.452825e-07, 8.063911e-07, 2.016058e-06,
  2.77858e-06, 9.419674e-06, 2.142617e-06, 2.541194e-06, 1.89134e-06, 
    1.493924e-07, 1.037957e-06, 1.316604e-06, 2.918207e-06, 3.523624e-06, 
    4.458025e-06, 4.154181e-06, 4.087705e-06, 2.058804e-06, 2.825804e-06,
  1.023586e-05, 1.42337e-05, 1.245857e-05, 8.123897e-06, 1.162887e-06, 
    7.344101e-07, 2.430932e-07, 8.809419e-07, 1.705374e-06, 2.201768e-06, 
    3.744961e-06, 3.802121e-06, 1.829889e-06, 1.834353e-06, 3.39151e-06,
  2.081403e-05, 1.777669e-05, 1.532809e-05, 1.088033e-05, 2.15391e-06, 
    1.316271e-06, 4.087682e-07, 9.756868e-07, 2.420961e-06, 2.750422e-06, 
    2.691783e-06, 2.678114e-06, 5.093994e-06, 7.743492e-06, 5.120096e-06,
  1.788367e-05, 1.616439e-05, 1.473468e-05, 1.127074e-05, 1.139116e-05, 
    3.990029e-06, 1.548335e-06, 6.877104e-07, 1.793219e-06, 2.044437e-06, 
    3.00058e-06, 3.223289e-06, 2.705224e-06, 6.07837e-06, 3.919945e-06,
  1.672238e-05, 1.412579e-05, 1.355057e-05, 1.13089e-05, 1.068416e-05, 
    1.32228e-05, 2.66206e-06, 1.851501e-06, 2.677953e-06, 2.751166e-06, 
    4.567738e-06, 4.180816e-06, 2.142131e-06, 1.130754e-06, 6.58646e-06,
  1.304478e-05, 1.41927e-05, 1.432241e-05, 1.290115e-05, 1.213267e-05, 
    1.227119e-05, 1.035767e-05, 6.177894e-06, 2.799416e-07, 2.981608e-06, 
    6.013041e-06, 4.284357e-06, 3.238332e-06, 2.675579e-06, 2.933871e-06,
  1.318736e-05, 1.355458e-05, 1.397682e-05, 1.39412e-05, 1.412605e-05, 
    1.340062e-05, 1.066852e-05, 6.673246e-06, 8.591696e-06, 7.852006e-06, 
    4.248632e-06, 7.661565e-06, 6.757009e-06, 4.037841e-06, 3.630639e-06,
  1.30427e-05, 1.397821e-05, 1.415083e-05, 1.51775e-05, 1.649977e-05, 
    1.531894e-05, 1.175805e-05, 8.198056e-06, 8.165056e-06, 8.254695e-06, 
    3.11807e-06, 7.598513e-06, 5.741099e-06, 5.305281e-06, 5.286512e-06,
  5.634334e-05, 6.461261e-05, 5.697446e-05, 3.629631e-05, 1.920628e-05, 
    1.465611e-05, 1.419324e-05, 1.307266e-05, 7.863641e-06, 8.484423e-06, 
    6.945814e-07, 4.438205e-06, 4.735038e-06, 4.875713e-06, 4.020088e-06,
  8.764693e-05, 9.081877e-05, 7.929967e-05, 5.120238e-05, 2.561474e-05, 
    1.086447e-05, 1.1126e-05, 1.095444e-05, 5.071305e-06, 8.579331e-07, 
    1.310499e-06, 5.619085e-06, 4.340158e-06, 3.291143e-06, 1.183014e-05,
  2.225269e-06, 2.892379e-06, 1.524403e-07, 2.587593e-07, 1.4203e-06, 
    4.082505e-07, 7.31055e-07, 1.978219e-06, 2.103851e-06, 3.176472e-06, 
    4.301305e-06, 5.661399e-06, 6.743454e-06, 6.832377e-06, 1.163252e-05,
  6.275816e-06, 1.153149e-05, 1.233574e-05, 9.573107e-06, 3.546137e-06, 
    1.007009e-06, 1.127512e-07, 7.43574e-07, 1.108131e-06, 1.508472e-06, 
    3.397086e-06, 4.136726e-06, 5.733872e-06, 5.125845e-06, 1.056169e-05,
  1.398998e-05, 1.686552e-05, 1.240102e-05, 1.395197e-05, 5.842602e-06, 
    3.481336e-06, 1.837889e-07, 8.079307e-07, 1.254941e-06, 1.008941e-06, 
    1.18998e-06, 2.280234e-06, 6.541944e-06, 1.13755e-05, 9.984505e-06,
  1.642843e-05, 1.560874e-05, 1.395927e-05, 1.774874e-05, 1.723473e-05, 
    4.412449e-06, 1.570061e-06, 4.230978e-07, 4.742667e-07, 6.092508e-07, 
    1.160475e-06, 1.199646e-06, 2.543686e-06, 9.145764e-06, 5.537893e-06,
  1.343384e-05, 1.610334e-05, 2.10746e-05, 1.955415e-05, 1.785224e-05, 
    8.190154e-06, 2.515264e-06, 1.601185e-06, 2.78612e-06, 4.826368e-07, 
    7.500761e-07, 4.484262e-07, 7.928239e-07, 1.734219e-06, 7.445217e-06,
  6.418928e-06, 1.359723e-05, 2.084397e-05, 2.069545e-05, 2.023797e-05, 
    1.348001e-05, 5.161909e-06, 1.313146e-06, 9.728076e-08, 1.206034e-06, 
    2.032461e-06, 1.084246e-07, 3.531841e-07, 8.079149e-07, 5.904346e-06,
  2.030655e-05, 1.592009e-05, 1.266675e-05, 1.38811e-05, 1.582172e-05, 
    1.279312e-05, 9.994381e-06, 1.198962e-05, 4.209625e-06, 6.300318e-06, 
    2.737486e-08, 3.153783e-08, 1.358806e-07, 2.956658e-07, 7.475192e-07,
  4.62646e-05, 4.615689e-05, 4.006907e-05, 2.395116e-05, 1.465185e-05, 
    1.483932e-05, 9.728508e-06, 5.051705e-06, 9.058657e-06, 5.880824e-06, 
    7.000906e-09, 2.054156e-08, 5.71902e-08, 9.548418e-08, 1.915701e-07,
  2.893395e-05, 4.288947e-05, 4.876393e-05, 2.644561e-05, 2.074928e-05, 
    1.257386e-05, 7.321855e-06, 9.229324e-06, 9.628874e-06, 1.031796e-05, 
    1.032004e-07, 9.538481e-09, 3.657588e-08, 1.171627e-07, 9.138574e-07,
  3.507137e-06, 6.316194e-06, 8.916379e-06, 1.373738e-05, 1.765994e-05, 
    9.046523e-06, 5.955465e-06, 9.681086e-06, 8.563119e-06, 7.126378e-07, 
    4.589815e-07, 2.777547e-08, 1.406318e-08, 1.534899e-07, 3.418753e-06,
  2.361968e-06, 3.679297e-06, 2.085587e-06, 3.434955e-06, 1.410155e-06, 
    1.70226e-06, 3.074804e-06, 1.657314e-06, 3.391615e-07, 1.906705e-06, 
    3.151204e-06, 4.471759e-06, 6.487726e-06, 7.042913e-06, 1.132477e-05,
  5.276638e-06, 9.756613e-06, 1.247526e-05, 1.653389e-05, 4.717509e-06, 
    2.333068e-06, 1.183522e-06, 2.662659e-06, 2.372444e-07, 2.39283e-07, 
    1.819876e-06, 2.833425e-06, 3.935127e-06, 6.545625e-06, 9.150286e-06,
  1.39207e-05, 1.50208e-05, 1.410074e-05, 2.709829e-05, 1.042501e-05, 
    5.898223e-06, 1.091277e-06, 5.368198e-07, 2.822784e-08, 4.807691e-08, 
    2.407708e-07, 1.355583e-06, 7.46391e-06, 8.867955e-06, 1.162883e-05,
  2.274672e-05, 1.789954e-05, 1.490572e-05, 1.252749e-05, 1.834064e-05, 
    3.37133e-06, 4.493654e-06, 9.762273e-08, 2.547351e-08, 2.409576e-08, 
    4.38705e-07, 6.636859e-07, 6.102874e-06, 1.285677e-05, 9.443009e-06,
  2.284157e-05, 2.201252e-05, 1.832084e-05, 1.23559e-05, 1.784549e-05, 
    1.392559e-05, 3.124778e-06, 2.783818e-06, 1.426091e-06, 6.602233e-07, 
    1.407351e-06, 1.405652e-07, 6.726287e-07, 3.153521e-06, 8.483963e-06,
  1.815807e-05, 1.964586e-05, 2.132296e-05, 1.423461e-05, 1.491237e-05, 
    1.445729e-05, 9.55023e-06, 9.831979e-07, 1.648672e-06, 7.1541e-08, 
    9.583993e-07, 2.696834e-07, 3.577169e-07, 8.888104e-07, 5.442631e-06,
  1.40147e-05, 1.849571e-05, 1.84875e-05, 1.516381e-05, 1.237466e-05, 
    9.604869e-06, 1.064506e-05, 1.108241e-05, 4.955933e-06, 1.563534e-06, 
    1.997664e-07, 5.593478e-07, 7.249608e-07, 2.865512e-07, 1.055049e-06,
  1.777885e-05, 2.076536e-05, 1.941081e-05, 1.364058e-05, 1.273982e-05, 
    9.239765e-06, 1.195238e-05, 1.058354e-05, 7.609872e-06, 6.026878e-06, 
    2.968357e-06, 1.642873e-06, 1.740739e-06, 5.166535e-07, 6.40182e-07,
  2.041461e-05, 2.299178e-05, 1.754985e-05, 1.447968e-05, 9.408461e-06, 
    9.41249e-06, 8.721047e-06, 8.900474e-06, 8.728232e-06, 4.757491e-06, 
    2.414378e-06, 2.254914e-06, 1.993671e-06, 1.325261e-06, 2.110409e-06,
  1.013169e-05, 1.205676e-05, 1.29036e-05, 1.10453e-05, 7.653897e-06, 
    4.354697e-06, 4.902782e-06, 4.732983e-06, 5.208041e-07, 9.67793e-08, 
    1.361636e-06, 1.846944e-06, 1.388528e-06, 1.041733e-06, 8.092092e-07,
  1.679785e-05, 1.295379e-05, 4.541805e-06, 2.673489e-06, 3.623758e-06, 
    3.10659e-06, 3.240261e-06, 2.89048e-06, 1.864396e-07, 1.887635e-06, 
    2.698043e-06, 1.879677e-06, 3.736282e-06, 4.596312e-06, 8.190429e-06,
  1.778411e-05, 1.503239e-05, 9.274941e-06, 9.292849e-06, 1.732097e-06, 
    2.774492e-06, 2.820868e-06, 2.870109e-06, 5.473509e-07, 3.807248e-07, 
    1.508642e-06, 1.584461e-06, 2.310973e-06, 5.929754e-06, 8.255264e-06,
  2.834806e-05, 2.55667e-05, 2.716348e-05, 1.71766e-05, 6.664808e-06, 
    1.691246e-06, 3.884079e-07, 3.474756e-06, 5.310843e-07, 5.584491e-07, 
    7.826204e-07, 1.856303e-06, 3.733137e-06, 7.965262e-06, 1.032341e-05,
  3.623783e-05, 3.662251e-05, 3.352518e-05, 2.847776e-05, 1.51221e-05, 
    3.517984e-06, 3.094873e-06, 7.119495e-07, 2.181694e-07, 3.51844e-07, 
    3.508667e-07, 2.338775e-06, 4.633009e-06, 8.765182e-06, 9.793521e-06,
  4.321398e-05, 3.531141e-05, 2.605879e-05, 1.969615e-05, 1.853898e-05, 
    1.429836e-05, 5.719566e-06, 9.184429e-06, 7.521792e-06, 1.453436e-06, 
    8.814479e-07, 3.578764e-06, 6.279165e-06, 9.542036e-06, 1.164057e-05,
  4.115492e-05, 3.426007e-05, 2.410801e-05, 1.625662e-05, 1.280413e-05, 
    1.002139e-05, 9.484224e-06, 6.920191e-06, 2.248738e-06, 3.626084e-06, 
    3.923686e-06, 5.483984e-06, 8.837703e-06, 1.00932e-05, 1.176014e-05,
  3.794126e-05, 3.155717e-05, 2.443832e-05, 1.784052e-05, 1.34026e-05, 
    1.019956e-05, 1.010665e-05, 7.963862e-06, 2.957097e-06, 3.776676e-06, 
    5.659197e-06, 6.578452e-06, 9.363164e-06, 9.934309e-06, 1.176835e-05,
  2.879559e-05, 2.663204e-05, 2.356624e-05, 1.919951e-05, 1.440352e-05, 
    1.111596e-05, 9.514882e-06, 9.452988e-06, 6.545205e-06, 1.674366e-06, 
    2.841098e-06, 3.948043e-06, 5.329572e-06, 1.005735e-05, 1.258036e-05,
  2.08936e-05, 2.035832e-05, 2.101844e-05, 1.667817e-05, 1.388909e-05, 
    1.172051e-05, 9.25818e-06, 7.254724e-06, 6.270389e-06, 5.410525e-07, 
    3.376672e-07, 6.817547e-07, 2.54626e-06, 7.395258e-06, 1.251245e-05,
  1.259752e-05, 1.474983e-05, 1.407852e-05, 1.204776e-05, 9.447641e-06, 
    7.271488e-06, 7.311155e-06, 4.853964e-06, 9.683804e-07, 4.104438e-07, 
    5.032321e-07, 2.907997e-06, 6.463425e-06, 7.351309e-06, 1.016837e-05,
  1.019132e-05, 1.429162e-05, 7.18898e-06, 4.190149e-06, 2.855155e-06, 
    4.730629e-07, 8.679834e-07, 6.944843e-07, 1.480787e-06, 1.767908e-06, 
    2.002815e-06, 3.654836e-06, 1.133303e-05, 2.055789e-05, 1.681869e-05,
  1.971646e-05, 2.52029e-05, 1.563731e-05, 8.502132e-06, 1.796802e-06, 
    5.143004e-07, 1.665328e-06, 1.715135e-06, 1.407405e-06, 1.799293e-06, 
    1.969346e-06, 3.838713e-06, 1.116106e-05, 2.34181e-05, 1.536804e-05,
  3.900062e-05, 3.768644e-05, 2.615728e-05, 1.564158e-05, 4.830132e-06, 
    1.119975e-06, 1.112553e-07, 1.926906e-06, 2.876144e-06, 9.439881e-07, 
    2.224371e-06, 5.046015e-06, 1.199461e-05, 2.207496e-05, 1.270153e-05,
  4.952309e-05, 4.725549e-05, 3.580248e-05, 2.157031e-05, 5.419633e-06, 
    3.06757e-06, 1.818912e-06, 2.172987e-06, 2.039958e-06, 2.059983e-06, 
    4.639509e-06, 6.24634e-06, 1.203247e-05, 2.29471e-05, 1.076451e-05,
  5.44633e-05, 5.451138e-05, 4.606473e-05, 2.828587e-05, 1.716509e-05, 
    5.091977e-06, 2.341503e-06, 2.144214e-06, 5.867833e-06, 6.944091e-06, 
    6.395433e-06, 7.277795e-06, 9.896517e-06, 1.829534e-05, 1.094894e-05,
  5.131691e-05, 5.078133e-05, 4.452249e-05, 3.326208e-05, 1.73707e-05, 
    1.08669e-05, 7.237678e-06, 1.171141e-06, 3.042656e-06, 5.521682e-06, 
    5.905438e-06, 6.807515e-06, 8.688965e-06, 1.405308e-05, 1.410963e-05,
  5.229908e-05, 4.786335e-05, 3.821086e-05, 2.862693e-05, 2.051821e-05, 
    1.156676e-05, 1.186177e-05, 1.050138e-05, 5.680392e-06, 2.581159e-06, 
    2.876499e-06, 4.14987e-06, 6.37824e-06, 1.211233e-05, 1.56442e-05,
  4.63158e-05, 4.14145e-05, 3.598603e-05, 2.839445e-05, 2.295552e-05, 
    1.682359e-05, 1.218047e-05, 9.986374e-06, 8.661502e-06, 8.260026e-07, 
    7.839676e-07, 1.221917e-06, 4.202304e-06, 9.894963e-06, 1.623417e-05,
  3.763423e-05, 3.663676e-05, 3.184832e-05, 2.337728e-05, 1.812362e-05, 
    1.500236e-05, 1.120729e-05, 1.089025e-05, 9.619418e-06, 4.656197e-07, 
    5.644252e-07, 1.814748e-06, 6.220171e-06, 8.070889e-06, 1.331984e-05,
  2.805151e-05, 2.205809e-05, 1.853048e-05, 1.738057e-05, 1.329053e-05, 
    1.064093e-05, 1.022843e-05, 9.525797e-06, 2.149165e-06, 1.910092e-07, 
    9.586181e-07, 2.941222e-06, 4.891826e-06, 5.536183e-06, 9.570052e-06,
  2.420271e-06, 1.002945e-06, 3.389465e-07, 3.312222e-07, 7.199221e-07, 
    8.650488e-08, 2.890324e-07, 7.456234e-07, 1.693031e-06, 3.693009e-06, 
    4.518564e-06, 5.597477e-06, 5.721421e-06, 6.457637e-06, 8.82586e-06,
  7.509135e-06, 4.081869e-06, 5.199538e-06, 1.41148e-06, 3.083072e-07, 
    3.392402e-07, 2.539348e-07, 4.442673e-07, 9.218161e-07, 4.043176e-06, 
    6.082799e-06, 7.19323e-06, 6.111098e-06, 7.830624e-06, 1.137367e-05,
  1.621273e-05, 1.184945e-05, 7.478134e-06, 7.02918e-06, 3.037742e-06, 
    8.3124e-07, 3.009641e-07, 4.297036e-07, 1.636061e-06, 4.318609e-06, 
    6.736758e-06, 7.384607e-06, 6.998866e-06, 8.246197e-06, 1.053737e-05,
  2.165582e-05, 1.82455e-05, 1.686122e-05, 1.536254e-05, 7.523749e-06, 
    3.138747e-06, 1.260253e-06, 4.536065e-07, 7.49977e-07, 4.742897e-06, 
    7.113646e-06, 7.291883e-06, 6.750661e-06, 8.621471e-06, 9.830972e-06,
  2.451051e-05, 2.061811e-05, 2.15798e-05, 2.262256e-05, 1.61751e-05, 
    5.451211e-06, 1.864828e-06, 1.197806e-06, 3.939598e-06, 5.73594e-06, 
    6.638948e-06, 6.588614e-06, 6.712099e-06, 6.80788e-06, 9.339647e-06,
  2.789911e-05, 2.295696e-05, 2.283804e-05, 2.638529e-05, 2.591391e-05, 
    1.805915e-05, 7.482464e-06, 4.628711e-07, 5.913032e-07, 5.342659e-06, 
    6.468746e-06, 6.387842e-06, 5.55564e-06, 5.919002e-06, 8.388273e-06,
  2.863616e-05, 2.966729e-05, 2.758128e-05, 2.681372e-05, 2.71814e-05, 
    1.930936e-05, 1.434495e-05, 6.86964e-06, 3.509128e-06, 2.515147e-06, 
    5.752485e-06, 5.646635e-06, 5.189911e-06, 6.28566e-06, 7.515919e-06,
  3.45758e-05, 3.548714e-05, 3.371477e-05, 3.386008e-05, 3.071837e-05, 
    2.488208e-05, 1.673439e-05, 1.553962e-05, 1.550162e-05, 7.05091e-07, 
    1.132615e-06, 2.256493e-06, 2.879923e-06, 4.371236e-06, 7.79269e-06,
  3.332357e-05, 3.648308e-05, 3.961209e-05, 3.514978e-05, 2.816588e-05, 
    2.512722e-05, 2.085533e-05, 1.700093e-05, 1.344615e-05, 2.012654e-06, 
    1.617111e-07, 5.43757e-08, 4.829727e-07, 2.202753e-06, 4.587263e-06,
  2.530439e-05, 2.734741e-05, 2.694391e-05, 2.673512e-05, 2.574527e-05, 
    2.346001e-05, 2.082595e-05, 1.399853e-05, 6.455556e-06, 7.681368e-07, 
    1.901549e-07, 9.609745e-08, 4.16773e-07, 1.674094e-06, 4.197016e-06,
  1.720687e-06, 9.915171e-07, 7.302187e-07, 1.368717e-07, 1.37194e-07, 
    4.226952e-07, 2.212581e-06, 2.699999e-06, 3.959523e-06, 6.292029e-06, 
    7.356979e-06, 9.507394e-06, 1.625483e-05, 1.749035e-05, 1.273559e-05,
  6.986319e-06, 5.907416e-06, 6.189685e-06, 1.186788e-06, 6.586768e-08, 
    2.119105e-07, 2.066933e-07, 1.711378e-06, 1.700322e-06, 4.155101e-06, 
    6.379914e-06, 8.464649e-06, 1.258742e-05, 1.692286e-05, 1.298179e-05,
  1.520141e-05, 1.251777e-05, 9.096638e-06, 5.997574e-06, 3.8975e-06, 
    5.474674e-07, 3.487833e-07, 7.440032e-07, 1.496901e-06, 3.16432e-06, 
    4.747621e-06, 6.217695e-06, 1.223832e-05, 1.62746e-05, 1.427351e-05,
  2.38569e-05, 1.70512e-05, 1.616338e-05, 1.313991e-05, 9.923037e-06, 
    2.743128e-06, 2.994015e-06, 8.409573e-07, 3.322271e-07, 2.384102e-06, 
    3.81233e-06, 6.099342e-06, 1.22123e-05, 1.685415e-05, 1.487616e-05,
  2.950269e-05, 1.479674e-05, 1.403407e-05, 1.651181e-05, 1.785694e-05, 
    1.633741e-05, 5.356012e-06, 5.610401e-06, 1.099156e-06, 1.27361e-06, 
    3.051626e-06, 4.131256e-06, 9.338899e-06, 1.328868e-05, 1.400152e-05,
  2.929006e-05, 2.280487e-05, 2.264352e-05, 2.235397e-05, 2.097896e-05, 
    2.103296e-05, 1.97846e-05, 4.556274e-06, 1.573348e-06, 1.756465e-06, 
    2.055083e-06, 2.385766e-06, 6.028403e-06, 1.243947e-05, 1.431996e-05,
  2.740443e-05, 2.41747e-05, 2.159867e-05, 1.93778e-05, 2.017259e-05, 
    2.126551e-05, 2.263021e-05, 1.524948e-05, 6.542926e-06, 1.949131e-06, 
    1.134831e-06, 1.406908e-06, 3.701305e-06, 1.018199e-05, 1.444127e-05,
  2.743059e-05, 2.302405e-05, 1.950187e-05, 1.988472e-05, 1.851487e-05, 
    1.947337e-05, 1.951334e-05, 1.909185e-05, 1.20168e-05, 2.09389e-06, 
    1.516444e-06, 8.128459e-07, 1.479639e-06, 5.251607e-06, 1.206442e-05,
  2.249177e-05, 2.378021e-05, 2.566028e-05, 2.152541e-05, 1.883411e-05, 
    2.024529e-05, 1.542031e-05, 1.567495e-05, 1.358881e-05, 1.617355e-06, 
    1.13481e-06, 6.243171e-07, 2.510206e-07, 1.657021e-06, 1.122954e-05,
  1.906133e-05, 2.056616e-05, 2.510234e-05, 2.899638e-05, 2.612138e-05, 
    2.378261e-05, 2.301912e-05, 1.739239e-05, 8.930825e-06, 2.990115e-06, 
    2.28923e-06, 8.021394e-07, 2.844052e-07, 2.370533e-07, 7.402016e-06,
  4.38411e-07, 1.67716e-06, 1.665448e-06, 6.461823e-08, 5.82079e-07, 
    6.220338e-07, 9.366979e-07, 1.790739e-06, 1.424283e-06, 1.074343e-06, 
    2.523721e-06, 4.573515e-06, 8.630541e-07, 3.085891e-08, 8.929901e-08,
  7.017721e-06, 1.245286e-05, 9.157158e-06, 1.675363e-06, 1.67544e-07, 
    6.254828e-07, 9.128062e-07, 2.56023e-06, 2.031304e-06, 9.497741e-07, 
    2.631765e-06, 4.530889e-06, 8.548363e-07, 3.588297e-08, 4.757691e-08,
  1.452641e-05, 1.777485e-05, 1.71487e-05, 9.84588e-06, 3.361682e-06, 
    2.107524e-06, 9.163303e-07, 6.84764e-06, 7.822085e-06, 1.084105e-06, 
    1.35635e-06, 3.609963e-06, 8.114611e-07, 9.630833e-07, 1.55404e-07,
  1.802359e-05, 1.767656e-05, 1.507476e-05, 1.465118e-05, 1.751153e-05, 
    8.239923e-06, 2.518504e-06, 7.945687e-06, 9.045046e-06, 4.970079e-06, 
    8.788862e-07, 2.057881e-06, 1.183631e-06, 8.978193e-07, 7.437217e-07,
  2.136916e-05, 1.591574e-05, 1.554368e-05, 1.485878e-05, 1.70911e-05, 
    1.637649e-05, 2.073669e-05, 9.295667e-06, 1.24919e-05, 7.357884e-06, 
    1.060381e-06, 1.413313e-06, 1.412179e-06, 4.965866e-07, 6.253246e-07,
  2.011425e-05, 1.526475e-05, 1.547843e-05, 1.561834e-05, 1.669218e-05, 
    2.338361e-05, 1.689074e-05, 9.387047e-06, 3.330074e-06, 5.865343e-06, 
    1.365608e-06, 8.407962e-07, 2.404515e-06, 4.227545e-07, 3.996568e-07,
  1.980259e-05, 2.156249e-05, 1.862725e-05, 1.628166e-05, 2.117784e-05, 
    2.544279e-05, 2.599592e-05, 1.802276e-05, 1.039455e-05, 2.476559e-06, 
    1.882746e-06, 6.88501e-07, 3.806047e-06, 8.385411e-07, 4.332983e-07,
  1.996472e-05, 2.112027e-05, 1.990349e-05, 2.038105e-05, 2.351382e-05, 
    2.248088e-05, 1.58135e-05, 1.227577e-05, 7.205235e-06, 1.336139e-06, 
    2.985456e-06, 1.00515e-06, 1.650165e-06, 2.606996e-06, 2.200362e-07,
  2.434849e-05, 2.746887e-05, 2.59307e-05, 2.391366e-05, 2.127541e-05, 
    1.754971e-05, 1.049784e-05, 1.011976e-05, 9.440493e-06, 9.332725e-07, 
    1.471202e-06, 6.200959e-07, 4.963056e-07, 4.782186e-06, 1.702597e-06,
  2.321937e-05, 2.001971e-05, 1.694103e-05, 1.445459e-05, 1.010794e-05, 
    7.040107e-06, 8.518131e-06, 1.448038e-05, 5.035609e-06, 3.301286e-06, 
    1.926825e-06, 7.346143e-07, 3.52854e-07, 1.047857e-06, 3.945687e-06,
  1.516913e-06, 8.239923e-08, 2.581756e-10, 2.231725e-09, 2.844952e-07, 
    1.87156e-06, 1.706787e-05, 1.122739e-05, 1.751535e-06, 3.084805e-07, 
    8.003174e-08, 2.520468e-08, 3.045683e-07, 3.413798e-07, 1.390794e-06,
  1.147556e-05, 8.338392e-06, 1.349617e-06, 3.970079e-08, 2.929791e-07, 
    4.31442e-07, 1.133363e-05, 1.252288e-05, 2.075102e-06, 1.306427e-06, 
    3.425369e-07, 5.211479e-07, 2.116771e-07, 6.600342e-07, 1.779291e-06,
  1.957787e-05, 1.13514e-05, 7.043172e-06, 5.108544e-06, 2.202856e-07, 
    1.885953e-06, 4.600724e-06, 1.412171e-05, 9.645621e-06, 2.21012e-06, 
    1.369624e-06, 3.146798e-07, 1.567769e-07, 4.181463e-07, 1.590939e-06,
  1.986166e-05, 1.08413e-05, 9.169778e-06, 1.257795e-05, 1.539692e-05, 
    8.560031e-06, 9.810551e-06, 1.322464e-05, 1.193209e-05, 5.834429e-06, 
    1.52991e-06, 3.820314e-07, 1.179862e-07, 5.333941e-07, 1.130075e-06,
  2.096957e-05, 1.27376e-05, 1.05563e-05, 1.104291e-05, 2.223866e-05, 
    2.857326e-05, 1.900484e-05, 1.507734e-05, 1.128167e-05, 2.60068e-06, 
    7.352668e-07, 5.644448e-08, 6.762643e-08, 3.276992e-07, 1.296354e-06,
  2.309719e-05, 1.834346e-05, 1.597187e-05, 1.409378e-05, 2.445394e-05, 
    2.956753e-05, 2.225094e-05, 7.814523e-06, 9.260028e-07, 1.072765e-06, 
    1.456579e-06, 3.894836e-07, 5.505185e-08, 1.838108e-07, 1.266771e-06,
  2.176537e-05, 1.966818e-05, 1.64994e-05, 1.876371e-05, 2.343288e-05, 
    2.168384e-05, 1.614148e-05, 1.010603e-05, 2.700652e-06, 9.386067e-07, 
    2.299684e-06, 3.646672e-07, 2.784558e-07, 2.251251e-07, 6.935503e-07,
  2.077392e-05, 2.124612e-05, 1.92902e-05, 1.886455e-05, 2.25543e-05, 
    1.753712e-05, 9.46561e-06, 8.829628e-06, 6.347862e-06, 4.441195e-06, 
    5.434812e-06, 2.078072e-06, 6.554079e-07, 6.47703e-07, 5.08523e-07,
  1.609646e-05, 2.016982e-05, 2.068162e-05, 1.765802e-05, 1.85114e-05, 
    1.251905e-05, 7.90888e-06, 6.676141e-06, 9.282283e-06, 6.08155e-06, 
    6.800586e-06, 4.955837e-06, 3.084803e-06, 2.531189e-06, 4.189246e-07,
  2.148743e-05, 1.927221e-05, 1.6584e-05, 1.356815e-05, 1.108919e-05, 
    6.819135e-06, 5.94451e-06, 9.537712e-06, 7.251434e-06, 6.818907e-06, 
    8.850903e-06, 8.929336e-06, 6.051358e-06, 3.252666e-06, 1.049695e-06,
  1.786156e-06, 7.566111e-07, 8.355103e-07, 9.464239e-07, 6.918989e-08, 
    2.448829e-06, 7.757296e-06, 2.240316e-06, 1.634962e-06, 3.870071e-06, 
    6.457278e-06, 8.822904e-06, 7.238436e-06, 5.333779e-06, 5.424189e-06,
  5.092377e-06, 3.45888e-06, 4.764355e-06, 3.207106e-07, 1.936408e-08, 
    6.954681e-07, 1.831928e-06, 8.46382e-07, 9.156275e-07, 2.757125e-06, 
    5.50525e-06, 8.863612e-06, 7.123725e-06, 5.463524e-06, 6.344337e-06,
  1.092712e-05, 1.075936e-05, 1.326279e-05, 1.489504e-05, 7.377046e-07, 
    1.975972e-06, 2.797502e-07, 1.467832e-06, 2.206071e-06, 4.136064e-06, 
    6.302214e-06, 7.975711e-06, 7.387626e-06, 6.120313e-06, 7.618251e-06,
  1.8346e-05, 2.217593e-05, 1.960682e-05, 1.82465e-05, 1.385918e-05, 
    2.671441e-06, 8.612859e-07, 1.786928e-06, 1.501696e-06, 2.601482e-06, 
    8.801257e-06, 8.18821e-06, 7.602389e-06, 5.929284e-06, 7.097375e-06,
  3.143772e-05, 2.657136e-05, 2.126952e-05, 1.702488e-05, 2.053999e-05, 
    2.113798e-05, 1.585999e-05, 8.574366e-06, 9.980178e-06, 3.61523e-06, 
    1.103004e-05, 9.8193e-06, 8.927305e-06, 4.426821e-06, 6.628848e-06,
  3.180317e-05, 2.816008e-05, 2.15683e-05, 1.654928e-05, 1.964123e-05, 
    2.334628e-05, 1.87631e-05, 4.802107e-06, 3.731929e-06, 7.688977e-06, 
    1.302225e-05, 1.148125e-05, 9.571459e-06, 3.779211e-06, 5.849648e-06,
  3.328741e-05, 2.738107e-05, 2.336301e-05, 2.185489e-05, 1.933665e-05, 
    1.666956e-05, 1.961949e-05, 1.368678e-05, 4.006573e-06, 5.541144e-06, 
    1.035405e-05, 1.16807e-05, 8.4745e-06, 3.445447e-06, 4.358356e-06,
  2.519741e-05, 2.835957e-05, 2.568187e-05, 2.343929e-05, 2.146817e-05, 
    1.819345e-05, 1.780016e-05, 1.740474e-05, 5.024447e-06, 5.1125e-06, 
    7.78751e-06, 9.21228e-06, 7.563617e-06, 3.722954e-06, 3.493279e-06,
  2.499749e-05, 2.863413e-05, 2.72618e-05, 2.058027e-05, 2.003493e-05, 
    1.895485e-05, 1.512995e-05, 9.581368e-06, 1.829679e-05, 6.448705e-06, 
    5.458979e-06, 6.154036e-06, 6.142579e-06, 4.730866e-06, 2.635524e-06,
  2.047012e-05, 2.031241e-05, 1.759104e-05, 1.396208e-05, 1.283725e-05, 
    6.678508e-06, 2.990557e-06, 1.032636e-05, 8.04331e-06, 7.877687e-06, 
    7.765108e-06, 5.838626e-06, 5.302623e-06, 6.694871e-06, 1.723812e-06,
  9.294788e-06, 5.740592e-06, 4.055748e-06, 2.263421e-06, 1.17433e-06, 
    8.964182e-07, 7.44204e-07, 9.900297e-07, 1.578103e-06, 2.440797e-06, 
    2.225877e-06, 4.935137e-06, 1.278752e-05, 2.294654e-05, 1.788398e-05,
  1.265502e-05, 8.21773e-06, 7.093321e-06, 2.499281e-06, 9.339585e-07, 
    4.719262e-07, 4.551272e-07, 8.745171e-07, 1.916179e-06, 3.11917e-06, 
    3.160189e-06, 5.471063e-06, 1.343699e-05, 2.306222e-05, 1.874291e-05,
  2.320087e-05, 1.75364e-05, 2.130457e-05, 2.160958e-05, 2.163746e-06, 
    1.688529e-06, 1.712901e-07, 5.582117e-07, 2.265781e-06, 3.315169e-06, 
    4.444675e-06, 6.206546e-06, 1.524769e-05, 2.220246e-05, 2.091346e-05,
  2.57492e-05, 2.550523e-05, 2.67732e-05, 3.095067e-05, 2.720648e-05, 
    1.301551e-06, 8.082632e-07, 2.399517e-07, 4.189421e-07, 1.122515e-06, 
    4.960079e-06, 7.570431e-06, 1.589122e-05, 2.36309e-05, 2.289235e-05,
  2.269676e-05, 2.493074e-05, 2.233956e-05, 2.518628e-05, 2.536989e-05, 
    2.127062e-05, 1.042751e-05, 4.274701e-06, 4.035893e-06, 1.898802e-06, 
    5.725107e-06, 8.600417e-06, 1.702437e-05, 2.53964e-05, 2.366808e-05,
  1.679301e-05, 1.776438e-05, 1.862263e-05, 1.95958e-05, 2.276614e-05, 
    2.425206e-05, 2.854917e-05, 1.864409e-05, 1.464821e-05, 1.071626e-05, 
    1.231022e-05, 1.372182e-05, 2.226736e-05, 3.077446e-05, 2.137819e-05,
  1.748345e-05, 1.764549e-05, 2.085743e-05, 1.908371e-05, 2.383705e-05, 
    2.49619e-05, 3.664997e-05, 3.516992e-05, 2.489639e-05, 1.867622e-05, 
    1.652955e-05, 1.955823e-05, 3.155662e-05, 3.730317e-05, 1.868592e-05,
  1.99654e-05, 2.347804e-05, 2.505792e-05, 2.209529e-05, 2.449393e-05, 
    3.36563e-05, 3.308253e-05, 4.057371e-05, 1.632113e-05, 1.27715e-05, 
    1.422634e-05, 2.380483e-05, 4.114206e-05, 4.372064e-05, 1.602162e-05,
  2.511337e-05, 2.857622e-05, 3.193465e-05, 2.686151e-05, 3.51518e-05, 
    4.290594e-05, 3.39882e-05, 1.652732e-05, 2.204836e-05, 7.94173e-06, 
    9.938655e-06, 2.784829e-05, 4.868542e-05, 4.593512e-05, 1.35518e-05,
  2.00553e-05, 1.682523e-05, 2.159703e-05, 3.509543e-05, 3.799444e-05, 
    2.557807e-05, 1.626788e-05, 2.430983e-05, 1.306464e-05, 9.032186e-06, 
    1.487042e-05, 3.406893e-05, 4.824257e-05, 4.258291e-05, 1.360451e-05,
  3.441804e-06, 2.248602e-06, 2.13347e-06, 1.339033e-06, 5.473066e-07, 
    3.461908e-07, 1.643129e-07, 1.852453e-07, 2.764124e-07, 1.322685e-06, 
    1.797255e-06, 9.53166e-06, 3.270667e-05, 4.797104e-05, 5.487775e-05,
  8.206268e-06, 7.924887e-06, 5.633647e-06, 2.110813e-06, 2.989478e-07, 
    5.600141e-07, 8.136473e-07, 3.463855e-08, 1.412054e-07, 7.810838e-07, 
    9.284461e-06, 3.316314e-05, 4.603568e-05, 5.651926e-05, 6.719239e-05,
  1.536484e-05, 1.228569e-05, 1.521725e-05, 1.617552e-05, 1.44311e-06, 
    5.366752e-06, 2.715583e-07, 1.995776e-07, 2.242061e-06, 1.323949e-05, 
    3.788839e-05, 5.015494e-05, 3.478992e-05, 4.387964e-05, 7.542977e-05,
  1.765446e-05, 1.765128e-05, 1.879385e-05, 2.18802e-05, 1.82896e-05, 
    2.545962e-06, 2.573609e-06, 1.242096e-06, 5.578131e-06, 3.099021e-05, 
    6.561174e-05, 4.511387e-05, 2.278236e-05, 3.438175e-05, 7.172494e-05,
  2.340587e-05, 1.561691e-05, 1.608593e-05, 1.788854e-05, 2.196848e-05, 
    1.842094e-05, 1.476652e-05, 3.160589e-05, 4.142001e-05, 4.240819e-05, 
    5.919157e-05, 3.242374e-05, 1.963552e-05, 2.973429e-05, 5.989166e-05,
  2.972039e-05, 2.500016e-05, 1.635494e-05, 1.066704e-05, 1.228032e-05, 
    1.945243e-05, 3.611052e-05, 5.224088e-05, 7.312319e-05, 5.738284e-05, 
    3.057516e-05, 1.585257e-05, 1.542073e-05, 3.892674e-05, 5.57297e-05,
  2.786353e-05, 2.893061e-05, 2.495116e-05, 1.523405e-05, 1.223975e-05, 
    1.785093e-05, 3.425019e-05, 5.262253e-05, 5.321305e-05, 3.064218e-05, 
    1.596557e-05, 7.882101e-06, 1.427411e-05, 4.558187e-05, 4.708474e-05,
  2.456331e-05, 3.136875e-05, 3.336933e-05, 3.01795e-05, 1.850014e-05, 
    1.571459e-05, 2.214899e-05, 2.846047e-05, 2.450304e-05, 1.730599e-05, 
    1.098878e-05, 5.244992e-06, 1.462732e-05, 4.26252e-05, 3.123375e-05,
  2.613647e-05, 3.212157e-05, 4.024597e-05, 3.979907e-05, 3.202761e-05, 
    2.220535e-05, 1.83707e-05, 2.252407e-05, 1.964896e-05, 1.354765e-05, 
    7.595691e-06, 4.111536e-06, 1.397441e-05, 3.476398e-05, 1.453811e-05,
  3.189611e-05, 3.482134e-05, 4.223435e-05, 4.670258e-05, 4.342954e-05, 
    3.391573e-05, 2.497582e-05, 2.078951e-05, 1.762332e-05, 1.25958e-05, 
    6.32571e-06, 4.054081e-06, 1.797185e-05, 2.416468e-05, 6.888646e-06,
  1.390293e-05, 5.922469e-06, 3.293599e-06, 1.814476e-06, 1.328199e-07, 
    1.01259e-07, 4.813183e-07, 2.42518e-08, 9.602798e-08, 3.086985e-07, 
    3.456261e-07, 8.815678e-07, 1.034376e-05, 2.6197e-05, 4.000246e-05,
  3.665836e-05, 1.686222e-05, 1.248481e-05, 8.154074e-06, 1.032544e-06, 
    1.490382e-06, 9.019711e-07, 1.275445e-08, 1.016865e-08, 1.285926e-07, 
    2.044929e-07, 3.030663e-06, 1.98068e-05, 3.03539e-05, 2.227765e-05,
  4.032458e-05, 2.947237e-05, 1.804263e-05, 1.951051e-05, 7.682414e-06, 
    1.872583e-06, 8.003541e-07, 1.124607e-08, 6.137686e-09, 1.376276e-08, 
    3.556088e-07, 6.392653e-06, 2.275281e-05, 2.565727e-05, 1.427486e-05,
  4.780438e-05, 4.137945e-05, 3.393898e-05, 2.255439e-05, 2.461684e-05, 
    9.73592e-06, 3.390202e-06, 1.631019e-06, 1.914837e-06, 1.798134e-07, 
    2.462024e-06, 8.638266e-06, 1.691965e-05, 1.53267e-05, 9.415715e-06,
  4.863353e-05, 4.947363e-05, 4.025216e-05, 4.310551e-05, 4.486044e-05, 
    3.241612e-05, 1.244216e-05, 9.424442e-06, 1.497496e-06, 2.796873e-07, 
    4.868403e-06, 9.781922e-06, 1.182257e-05, 5.004738e-06, 5.561863e-06,
  4.825626e-05, 5.495115e-05, 4.832256e-05, 4.540909e-05, 4.682012e-05, 
    4.183661e-05, 3.603e-05, 1.219801e-05, 3.475983e-06, 2.356314e-06, 
    5.651351e-06, 1.007941e-05, 8.219785e-06, 5.229451e-06, 3.407461e-06,
  3.744841e-05, 5.453671e-05, 5.752804e-05, 5.830581e-05, 5.442773e-05, 
    4.760119e-05, 4.217146e-05, 4.258644e-05, 2.190766e-05, 9.08081e-06, 
    6.472112e-06, 1.088073e-05, 6.693135e-06, 6.266546e-06, 2.632731e-06,
  2.51399e-05, 2.266732e-05, 2.611514e-05, 3.163944e-05, 4.406465e-05, 
    4.389333e-05, 3.582659e-05, 3.284128e-05, 2.939561e-05, 2.242893e-05, 
    1.165638e-05, 1.094609e-05, 7.316155e-06, 5.311213e-06, 8.855538e-07,
  1.039104e-05, 1.465953e-05, 1.568413e-05, 1.583832e-05, 2.442549e-05, 
    3.608549e-05, 3.994476e-05, 3.569485e-05, 3.310678e-05, 3.459826e-05, 
    1.9844e-05, 1.237048e-05, 7.834827e-06, 3.790357e-06, 5.833718e-07,
  1.15347e-05, 1.529635e-05, 1.504481e-05, 1.388915e-05, 2.364015e-05, 
    3.724746e-05, 4.664895e-05, 4.983898e-05, 4.522369e-05, 4.381343e-05, 
    3.087224e-05, 1.522457e-05, 1.113167e-05, 6.540736e-06, 8.549744e-07,
  5.008507e-05, 2.516355e-05, 5.985595e-06, 4.089868e-06, 2.018773e-07, 
    1.633976e-08, 1.277063e-07, 2.627375e-08, 1.183735e-08, 1.796471e-08, 
    9.892455e-09, 8.199066e-08, 5.190209e-07, 2.157452e-06, 2.456286e-06,
  6.572218e-05, 5.117661e-05, 2.21608e-05, 7.776404e-06, 2.062726e-06, 
    1.901454e-06, 1.068064e-06, 1.216191e-08, 1.255635e-09, 7.366933e-11, 
    3.760066e-10, 9.398064e-08, 3.537266e-07, 1.839663e-06, 1.800069e-06,
  5.256108e-05, 6.051718e-05, 4.837662e-05, 2.648294e-05, 3.394129e-06, 
    5.692092e-07, 2.941088e-06, 1.674436e-06, 6.610885e-09, 9.409886e-12, 
    5.578776e-09, 3.017779e-08, 2.011351e-07, 1.316871e-06, 1.340122e-06,
  4.776864e-05, 6.915266e-05, 6.651314e-05, 3.472735e-05, 2.642589e-05, 
    3.512146e-06, 7.449457e-07, 3.40775e-06, 1.552858e-06, 1.402689e-08, 
    9.464841e-08, 2.332445e-08, 1.505013e-07, 1.047064e-06, 2.205838e-06,
  4.104929e-05, 8.459441e-05, 9.332711e-05, 6.644207e-05, 3.607185e-05, 
    2.517694e-05, 9.052481e-06, 1.295685e-06, 3.422612e-07, 5.395985e-09, 
    1.10703e-07, 5.9478e-08, 6.068162e-07, 1.197715e-06, 1.587351e-06,
  2.721829e-05, 7.468125e-05, 0.0001051132, 9.326907e-05, 6.273211e-05, 
    3.290532e-05, 2.392613e-05, 5.715423e-06, 7.297054e-07, 1.117709e-06, 
    7.503197e-07, 1.365034e-06, 2.023574e-06, 7.784187e-07, 1.132989e-06,
  3.153306e-05, 5.052637e-05, 9.130991e-05, 0.0001031852, 8.340398e-05, 
    4.832354e-05, 3.111623e-05, 2.28002e-05, 1.318877e-05, 5.089928e-06, 
    2.677283e-06, 2.243297e-06, 2.059552e-06, 6.512782e-07, 1.178354e-06,
  4.964078e-05, 4.695082e-05, 5.558258e-05, 7.478884e-05, 7.961268e-05, 
    6.257987e-05, 4.736431e-05, 3.271292e-05, 2.964822e-05, 1.117349e-05, 
    1.028506e-05, 6.259453e-06, 1.287659e-06, 1.066104e-06, 1.004596e-06,
  3.152233e-05, 3.521531e-05, 4.358233e-05, 4.098921e-05, 3.93182e-05, 
    4.250389e-05, 3.725691e-05, 3.041326e-05, 2.140937e-05, 1.661277e-05, 
    1.610321e-05, 9.625493e-06, 1.785761e-06, 2.144602e-06, 1.438753e-06,
  2.001548e-05, 1.71332e-05, 2.427856e-05, 2.056175e-05, 2.059799e-05, 
    1.780399e-05, 1.548716e-05, 1.714022e-05, 1.364261e-05, 1.640029e-05, 
    1.984144e-05, 1.201296e-05, 5.06038e-06, 2.767102e-06, 1.892e-06,
  1.192025e-05, 1.118469e-05, 6.876136e-06, 4.501471e-06, 1.113498e-06, 
    9.16724e-07, 1.6619e-06, 9.654567e-07, 8.24483e-07, 1.481353e-07, 
    3.347818e-07, 3.311857e-07, 3.571999e-07, 2.972883e-07, 3.59013e-07,
  1.687769e-05, 1.562489e-05, 1.098047e-05, 5.462571e-06, 2.060704e-06, 
    2.496768e-06, 2.256316e-06, 6.313729e-07, 1.78022e-07, 5.537667e-07, 
    1.728941e-07, 2.349667e-07, 2.87035e-07, 2.065316e-07, 1.944958e-07,
  2.66876e-05, 2.393276e-05, 2.144577e-05, 1.452289e-05, 4.440001e-07, 
    1.24517e-06, 9.459379e-07, 1.106821e-06, 2.309884e-07, 1.21338e-07, 
    3.707239e-07, 1.062347e-07, 1.060135e-07, 2.302253e-07, 1.091142e-07,
  3.147129e-05, 3.268941e-05, 3.235709e-05, 1.635549e-05, 1.42777e-05, 
    2.29406e-07, 1.269497e-06, 1.144945e-06, 7.2558e-07, 2.323677e-07, 
    1.205476e-07, 6.194976e-08, 6.939617e-08, 1.170986e-07, 5.368636e-07,
  4.072974e-05, 3.640669e-05, 3.574968e-05, 2.538344e-05, 1.821802e-05, 
    7.957979e-06, 2.614119e-06, 1.452516e-07, 3.836137e-08, 1.386532e-08, 
    2.503565e-07, 7.731126e-08, 4.980705e-08, 1.379862e-07, 2.215762e-07,
  5.722153e-05, 5.68361e-05, 4.961972e-05, 3.695234e-05, 2.480486e-05, 
    1.601458e-05, 8.328122e-06, 6.932445e-07, 1.109989e-09, 6.967645e-08, 
    7.664775e-07, 4.046304e-07, 4.333443e-08, 8.932794e-08, 2.828334e-08,
  5.442121e-05, 4.968644e-05, 4.606237e-05, 4.111139e-05, 3.245896e-05, 
    2.337871e-05, 2.20285e-05, 7.275855e-06, 1.201524e-06, 4.275213e-07, 
    1.592233e-07, 2.393513e-08, 3.419503e-08, 7.699099e-08, 4.348799e-08,
  5.882966e-05, 6.276659e-05, 5.913381e-05, 5.74509e-05, 4.122294e-05, 
    3.194021e-05, 2.412949e-05, 1.762999e-05, 1.524436e-05, 2.97157e-06, 
    3.641538e-07, 7.146139e-08, 4.08794e-08, 6.285274e-08, 5.016123e-08,
  5.158884e-05, 5.186469e-05, 5.253405e-05, 5.230794e-05, 5.179057e-05, 
    4.312865e-05, 3.205866e-05, 2.466595e-05, 2.260085e-05, 1.658788e-06, 
    2.07627e-07, 1.166821e-07, 1.270187e-07, 1.195522e-07, 9.099423e-08,
  3.945362e-05, 3.685265e-05, 3.816534e-05, 4.158928e-05, 4.091776e-05, 
    3.605875e-05, 2.696873e-05, 2.181022e-05, 5.577454e-06, 9.116752e-07, 
    2.03774e-06, 2.891715e-06, 1.456368e-06, 2.866678e-07, 3.433331e-07,
  3.073241e-06, 2.366558e-06, 1.513007e-06, 8.516952e-07, 5.995163e-07, 
    3.736895e-07, 1.955763e-07, 1.161762e-06, 1.189717e-06, 3.610666e-07, 
    8.801287e-08, 2.624878e-07, 8.70703e-08, 6.145421e-08, 9.720491e-08,
  5.187781e-06, 1.940839e-06, 2.177657e-06, 9.129253e-07, 4.323082e-07, 
    2.591953e-07, 7.577924e-07, 4.669051e-07, 4.979319e-07, 1.1911e-06, 
    5.982418e-08, 2.624593e-07, 4.138929e-07, 3.535759e-08, 5.840014e-08,
  1.168266e-05, 4.497601e-06, 5.076377e-06, 2.998086e-06, 6.149458e-07, 
    9.007721e-07, 5.028592e-07, 8.547692e-07, 6.800364e-07, 2.233143e-07, 
    1.900817e-07, 5.358361e-07, 3.469773e-08, 1.265555e-07, 4.027825e-08,
  1.454388e-05, 1.05434e-05, 7.835542e-06, 5.008073e-06, 2.347955e-06, 
    1.438945e-06, 4.8838e-07, 5.371515e-07, 2.523361e-07, 4.29697e-07, 
    9.644338e-08, 4.795116e-08, 5.770566e-08, 1.361887e-07, 1.209629e-07,
  2.17361e-05, 1.759371e-05, 1.24456e-05, 9.091703e-06, 7.483006e-06, 
    4.992925e-06, 3.459793e-06, 2.256041e-07, 2.236122e-07, 1.043666e-07, 
    6.728895e-09, 2.544681e-08, 1.023638e-08, 2.503271e-08, 7.734219e-08,
  2.59555e-05, 2.338458e-05, 1.789666e-05, 1.364557e-05, 1.116113e-05, 
    8.394745e-06, 4.250986e-06, 1.929266e-08, 4.877134e-09, 1.328534e-06, 
    5.783215e-08, 6.298198e-09, 2.389151e-09, 1.724529e-08, 8.390368e-09,
  2.974792e-05, 2.780215e-05, 2.352615e-05, 1.813051e-05, 1.398375e-05, 
    1.318976e-05, 7.266092e-06, 1.072143e-06, 2.903366e-07, 6.913799e-07, 
    4.148361e-07, 1.47799e-08, 9.012204e-09, 2.545121e-08, 2.195858e-08,
  3.963355e-05, 3.178267e-05, 2.699436e-05, 2.167427e-05, 1.633227e-05, 
    1.314862e-05, 1.266015e-05, 1.136738e-05, 5.885985e-06, 2.389195e-07, 
    1.185863e-07, 5.247317e-08, 1.474106e-08, 4.049233e-08, 6.313906e-08,
  4.190197e-05, 3.371961e-05, 3.025317e-05, 2.144376e-05, 1.801519e-05, 
    1.595782e-05, 1.356431e-05, 1.111443e-05, 6.96232e-06, 7.474874e-08, 
    3.373891e-08, 1.920361e-08, 2.033487e-08, 3.577927e-08, 6.564395e-08,
  3.296701e-05, 2.684479e-05, 2.593209e-05, 1.668336e-05, 1.848476e-05, 
    1.548354e-05, 1.193177e-05, 1.052453e-05, 8.915218e-07, 4.809379e-08, 
    2.736487e-07, 1.539635e-08, 2.319605e-08, 2.949299e-08, 4.393018e-08,
  7.335825e-06, 2.02987e-06, 1.58116e-06, 1.901392e-06, 4.837169e-07, 
    2.397131e-07, 7.034442e-07, 7.840907e-07, 9.993695e-07, 3.328494e-07, 
    5.465503e-07, 6.989419e-07, 8.008675e-07, 4.564703e-07, 4.134204e-07,
  1.04633e-05, 5.246503e-06, 6.98223e-06, 2.933819e-06, 5.045604e-09, 
    1.281859e-07, 5.505484e-07, 2.736058e-07, 3.176395e-07, 1.014791e-06, 
    6.984603e-07, 3.876747e-07, 1.157049e-06, 2.163073e-07, 4.310191e-07,
  2.280469e-05, 1.071666e-05, 9.202932e-06, 3.853037e-06, 1.116923e-06, 
    3.109111e-07, 1.417894e-07, 2.037499e-07, 2.913e-07, 1.020897e-07, 
    1.38829e-07, 2.030249e-07, 1.723715e-07, 6.239115e-07, 9.100618e-07,
  3.179514e-05, 2.362019e-05, 1.433156e-05, 1.269374e-05, 9.309621e-06, 
    8.299148e-07, 1.605672e-07, 2.922552e-08, 1.952631e-08, 1.393334e-07, 
    1.860825e-07, 3.525809e-07, 4.992326e-07, 8.581627e-07, 1.689423e-06,
  3.070411e-05, 1.971953e-05, 1.723733e-05, 1.798418e-05, 1.516318e-05, 
    8.193481e-06, 1.270704e-06, 7.044861e-09, 1.402071e-07, 5.012828e-07, 
    2.582908e-07, 2.940715e-07, 4.476748e-07, 6.075943e-07, 2.174946e-06,
  3.937306e-05, 3.314107e-05, 1.905828e-05, 1.934116e-05, 1.727497e-05, 
    1.390737e-05, 5.299637e-06, 3.750081e-09, 3.104486e-08, 4.130384e-07, 
    2.15935e-07, 5.240127e-08, 1.995053e-07, 3.161062e-07, 9.322849e-07,
  5.793567e-05, 4.875657e-05, 3.709278e-05, 2.227954e-05, 1.671234e-05, 
    1.366384e-05, 8.546269e-06, 2.95694e-06, 9.126514e-07, 4.193653e-07, 
    3.188558e-07, 6.234861e-08, 2.099005e-07, 2.041399e-07, 5.566478e-07,
  5.075933e-05, 4.012495e-05, 3.315638e-05, 2.603462e-05, 2.338939e-05, 
    1.754119e-05, 1.144027e-05, 7.938213e-06, 5.819967e-07, 5.940872e-07, 
    1.2432e-07, 7.105508e-07, 3.543229e-07, 3.537544e-07, 4.255529e-07,
  4.466638e-05, 4.264106e-05, 3.610233e-05, 2.793587e-05, 2.134959e-05, 
    1.944736e-05, 1.772488e-05, 9.936564e-06, 8.524823e-07, 2.43423e-07, 
    7.076497e-07, 1.344197e-06, 1.22533e-06, 7.964857e-07, 4.855149e-07,
  3.939582e-05, 3.510565e-05, 2.920582e-05, 2.117453e-05, 1.971162e-05, 
    1.741952e-05, 1.491604e-05, 7.813216e-06, 7.797183e-08, 1.144967e-06, 
    1.944267e-06, 5.039594e-07, 1.119898e-06, 1.837563e-06, 7.033552e-07,
  1.252771e-06, 8.375124e-07, 9.3792e-07, 1.503598e-06, 7.599083e-07, 
    3.280479e-07, 1.143104e-06, 1.485617e-06, 2.555762e-06, 9.023498e-07, 
    9.647041e-07, 1.59505e-06, 1.656455e-06, 1.540151e-06, 1.921917e-06,
  2.338542e-06, 1.919642e-06, 1.679138e-06, 2.362573e-06, 2.031077e-08, 
    2.912851e-07, 9.587612e-07, 9.722777e-07, 9.879318e-07, 3.750803e-06, 
    2.809023e-06, 5.20709e-06, 6.776093e-06, 3.939165e-06, 5.880247e-06,
  9.569389e-06, 4.506298e-06, 5.269639e-06, 3.244941e-06, 2.13405e-06, 
    1.967828e-07, 3.779172e-07, 3.531833e-06, 6.911312e-06, 7.568825e-06, 
    8.75402e-06, 1.005502e-05, 1.152926e-05, 1.235299e-05, 1.490097e-05,
  1.677307e-05, 1.185334e-05, 7.969613e-06, 5.816825e-06, 3.251364e-06, 
    1.832129e-06, 4.181825e-07, 2.510408e-06, 6.046925e-06, 1.278769e-05, 
    1.522248e-05, 1.637108e-05, 1.725318e-05, 1.636214e-05, 1.673411e-05,
  2.395245e-05, 1.534704e-05, 1.283377e-05, 1.245132e-05, 7.376029e-06, 
    4.732473e-06, 1.288454e-06, 5.236937e-07, 2.723011e-06, 9.305335e-06, 
    1.458918e-05, 1.661452e-05, 1.806539e-05, 1.242161e-05, 1.091379e-05,
  2.667155e-05, 1.242287e-05, 1.175075e-05, 1.595041e-05, 1.029429e-05, 
    1.147909e-05, 6.743927e-06, 4.692341e-06, 3.900989e-06, 7.821217e-06, 
    8.927003e-06, 1.266375e-05, 1.416046e-05, 1.08354e-05, 9.019418e-06,
  3.295262e-05, 2.141258e-05, 1.76644e-05, 1.398386e-05, 1.360033e-05, 
    1.261355e-05, 1.098141e-05, 1.020948e-05, 5.755858e-06, 5.445556e-06, 
    5.296864e-06, 7.723022e-06, 9.092464e-06, 9.926157e-06, 8.83274e-06,
  4.780712e-05, 3.235445e-05, 1.997912e-05, 2.031132e-05, 1.758835e-05, 
    1.688655e-05, 1.314818e-05, 5.174766e-06, 2.971013e-06, 2.576548e-06, 
    2.946382e-06, 4.040191e-06, 5.664944e-06, 7.620935e-06, 8.764647e-06,
  5.419815e-05, 3.658526e-05, 3.073385e-05, 1.984753e-05, 1.909718e-05, 
    1.852e-05, 1.158098e-05, 5.595784e-06, 1.065061e-06, 4.384083e-07, 
    1.332644e-06, 1.674156e-06, 2.325124e-06, 3.971503e-06, 4.927203e-06,
  4.593025e-05, 3.283632e-05, 2.477263e-05, 2.0165e-05, 1.656241e-05, 
    1.764775e-05, 1.171203e-05, 3.293611e-06, 6.247342e-08, 5.798095e-07, 
    4.933594e-07, 3.970437e-07, 5.934147e-07, 8.263447e-07, 1.484829e-06,
  1.112142e-06, 3.54557e-06, 4.605015e-07, 1.347457e-06, 2.331187e-06, 
    9.062121e-08, 4.828525e-07, 8.532039e-07, 1.1012e-06, 8.320613e-07, 
    2.103137e-06, 4.063877e-06, 3.783547e-06, 3.04504e-06, 2.513623e-06,
  6.126196e-06, 6.069471e-06, 5.665604e-06, 3.32812e-06, 1.184071e-07, 
    7.417203e-07, 1.507697e-06, 1.326708e-06, 1.254134e-06, 1.607961e-06, 
    1.712898e-06, 2.888592e-06, 3.964086e-06, 2.277851e-06, 1.635985e-06,
  1.414197e-05, 1.169379e-05, 9.327058e-06, 5.701193e-06, 4.938374e-06, 
    1.963227e-07, 7.047632e-07, 6.021728e-06, 6.706148e-06, 4.325289e-06, 
    2.558274e-06, 1.773424e-06, 2.48168e-06, 2.588106e-06, 1.509239e-06,
  1.977463e-05, 1.876228e-05, 1.517132e-05, 1.200371e-05, 1.628599e-05, 
    1.035115e-05, 2.416938e-06, 8.543631e-06, 1.070636e-05, 7.303572e-06, 
    3.288449e-06, 1.016724e-06, 1.157626e-06, 2.082306e-06, 2.222744e-06,
  2.086907e-05, 2.005091e-05, 1.94728e-05, 1.780784e-05, 1.92016e-05, 
    2.360513e-05, 2.014606e-05, 2.449528e-06, 4.046029e-06, 7.049384e-06, 
    5.444609e-06, 1.285588e-06, 8.863589e-07, 2.509549e-06, 1.307088e-06,
  2.119036e-05, 1.884613e-05, 2.122908e-05, 2.257399e-05, 2.248086e-05, 
    2.081177e-05, 2.171321e-05, 1.280129e-05, 1.135616e-05, 1.090607e-05, 
    6.94369e-06, 2.897674e-06, 2.602607e-06, 1.877568e-06, 7.656055e-08,
  2.360382e-05, 2.20822e-05, 2.421967e-05, 2.343425e-05, 2.707424e-05, 
    2.434795e-05, 1.958339e-05, 1.90195e-05, 1.718931e-05, 1.598262e-05, 
    1.229451e-05, 6.855072e-06, 3.498935e-06, 1.965772e-06, 2.935236e-07,
  2.959487e-05, 2.745985e-05, 2.672564e-05, 2.300825e-05, 2.468788e-05, 
    2.267422e-05, 1.965038e-05, 1.670421e-05, 1.443252e-05, 1.308129e-05, 
    1.249658e-05, 9.792674e-06, 5.40615e-06, 3.17512e-06, 2.959017e-06,
  2.950479e-05, 2.791048e-05, 3.334332e-05, 2.677176e-05, 2.082134e-05, 
    1.833197e-05, 1.599642e-05, 1.490201e-05, 1.476985e-05, 1.183649e-05, 
    1.063082e-05, 1.078421e-05, 7.229082e-06, 4.800391e-06, 2.698701e-06,
  2.570229e-05, 2.408132e-05, 2.541181e-05, 1.723715e-05, 1.778953e-05, 
    1.584948e-05, 1.265581e-05, 7.782138e-06, 7.052859e-06, 6.477689e-06, 
    8.239122e-06, 6.1356e-06, 4.855363e-06, 2.701922e-06, 1.236199e-06,
  2.552458e-06, 2.15915e-06, 1.798905e-06, 2.365765e-06, 4.843896e-06, 
    7.345443e-06, 9.850912e-06, 1.247477e-05, 1.165399e-05, 7.167692e-06, 
    3.968814e-06, 2.483094e-06, 2.584634e-06, 1.71713e-06, 1.229449e-06,
  7.695605e-06, 5.262685e-06, 4.70759e-06, 4.684219e-06, 6.122481e-06, 
    9.172004e-06, 1.583769e-05, 1.223481e-05, 8.351922e-06, 6.898809e-06, 
    3.270043e-06, 3.587377e-06, 3.107248e-06, 1.651845e-06, 8.097142e-07,
  1.537914e-05, 8.776921e-06, 1.005283e-05, 7.317123e-06, 1.093442e-05, 
    7.540401e-06, 1.357538e-05, 1.548327e-05, 1.108905e-05, 7.927496e-06, 
    4.640857e-06, 2.441388e-06, 2.903883e-06, 2.125654e-06, 4.374718e-07,
  2.155918e-05, 1.598148e-05, 1.708644e-05, 1.13782e-05, 1.569884e-05, 
    1.263227e-05, 6.775562e-06, 8.431654e-06, 8.983206e-06, 9.890299e-06, 
    4.309178e-06, 1.612541e-06, 1.514312e-06, 1.744063e-06, 9.030067e-07,
  2.178261e-05, 1.760431e-05, 1.921961e-05, 1.741105e-05, 1.611788e-05, 
    1.874971e-05, 1.234345e-05, 1.099162e-06, 1.750882e-06, 4.536674e-06, 
    3.689266e-06, 1.926766e-06, 1.355238e-06, 1.272187e-06, 7.951882e-07,
  1.931619e-05, 1.662285e-05, 1.765597e-05, 1.855838e-05, 1.697806e-05, 
    1.50701e-05, 1.358719e-05, 5.955847e-06, 3.331436e-06, 4.310376e-06, 
    2.911676e-06, 2.245661e-06, 2.251877e-06, 9.027752e-07, 1.408403e-07,
  2.308085e-05, 2.226843e-05, 1.991893e-05, 1.8259e-05, 1.767766e-05, 
    1.536686e-05, 1.158688e-05, 9.785806e-06, 7.270974e-06, 4.455776e-06, 
    4.325909e-06, 3.233569e-06, 1.986676e-06, 3.148243e-07, 1.884659e-07,
  2.831535e-05, 2.86454e-05, 2.356997e-05, 2.069365e-05, 1.927904e-05, 
    1.879985e-05, 1.468801e-05, 1.123609e-05, 6.235552e-06, 4.131061e-06, 
    4.314956e-06, 3.284491e-06, 1.641875e-06, 5.555129e-07, 1.749388e-07,
  3.034073e-05, 2.875175e-05, 3.194662e-05, 2.533752e-05, 2.113211e-05, 
    1.921649e-05, 1.644496e-05, 1.153368e-05, 6.250107e-06, 4.253925e-06, 
    4.389092e-06, 3.186372e-06, 1.953152e-06, 9.16301e-07, 1.430723e-07,
  2.405831e-05, 1.997682e-05, 2.47583e-05, 2.443882e-05, 2.144922e-05, 
    1.684965e-05, 1.315336e-05, 1.001868e-05, 6.659676e-06, 4.224592e-06, 
    6.751591e-06, 2.749673e-06, 9.513836e-07, 1.918721e-07, 2.39006e-08,
  1.347232e-06, 1.014448e-06, 2.557354e-07, 1.458039e-06, 4.032937e-07, 
    1.263928e-06, 2.128506e-06, 2.557943e-06, 3.963738e-06, 2.77404e-06, 
    2.673295e-06, 3.436824e-06, 2.091077e-06, 6.008461e-07, 3.483736e-07,
  4.061891e-06, 3.778237e-06, 4.207242e-06, 3.237249e-06, 1.845034e-06, 
    1.895464e-06, 2.777415e-06, 2.63453e-06, 2.728123e-06, 3.256454e-06, 
    1.235441e-06, 2.527102e-06, 1.230744e-06, 4.493284e-08, 1.104442e-07,
  1.256123e-05, 8.516502e-06, 1.110963e-05, 8.409015e-06, 9.539342e-06, 
    2.5892e-06, 2.257342e-06, 4.237612e-06, 4.184744e-06, 3.067157e-06, 
    2.13256e-06, 1.496265e-06, 1.281501e-06, 5.072346e-07, 1.228846e-08,
  2.147782e-05, 1.997599e-05, 2.113416e-05, 1.958014e-05, 1.865577e-05, 
    9.521503e-06, 2.414902e-06, 2.234632e-06, 2.22406e-06, 2.550655e-06, 
    8.7508e-07, 1.595376e-07, 4.614181e-07, 3.125099e-07, 2.100055e-08,
  2.521423e-05, 2.280263e-05, 2.46775e-05, 2.648572e-05, 2.498798e-05, 
    2.298889e-05, 1.136911e-05, 1.026843e-06, 1.157843e-06, 1.397946e-06, 
    6.2328e-07, 1.195163e-07, 2.927995e-08, 3.387267e-08, 2.06562e-11,
  2.460203e-05, 2.22305e-05, 2.50402e-05, 2.884415e-05, 2.869389e-05, 
    2.536679e-05, 2.238742e-05, 5.932524e-06, 1.707397e-06, 5.421876e-06, 
    6.481553e-07, 2.555888e-07, 1.033083e-08, 3.421521e-10, 7.490733e-11,
  2.62968e-05, 2.229375e-05, 2.40784e-05, 2.549287e-05, 3.072757e-05, 
    2.725783e-05, 2.102322e-05, 1.55967e-05, 9.307252e-06, 4.677515e-06, 
    2.796464e-06, 5.754954e-07, 1.140426e-09, 7.17395e-12, 7.941422e-11,
  2.776776e-05, 1.828416e-05, 2.062798e-05, 2.257918e-05, 2.393556e-05, 
    2.515766e-05, 2.065335e-05, 1.498998e-05, 8.437606e-06, 2.945273e-06, 
    2.083955e-06, 2.917063e-07, 1.297842e-09, 6.280661e-11, 2.32873e-10,
  3.045973e-05, 1.835553e-05, 2.214342e-05, 2.20918e-05, 2.077199e-05, 
    2.056131e-05, 1.958847e-05, 1.546222e-05, 6.250671e-06, 2.578156e-06, 
    1.357401e-06, 3.39172e-07, 1.852274e-09, 1.772703e-10, 8.727929e-09,
  2.465724e-05, 1.582496e-05, 1.846385e-05, 1.576286e-05, 1.919098e-05, 
    1.684388e-05, 1.587764e-05, 1.221861e-05, 5.494327e-06, 4.76079e-06, 
    3.144693e-06, 3.268055e-07, 3.082157e-09, 2.344748e-10, 5.643008e-10,
  2.358616e-07, 8.165462e-07, 5.380934e-07, 3.924926e-06, 6.501504e-06, 
    6.183597e-06, 5.321049e-06, 6.272162e-06, 7.25333e-06, 4.014978e-06, 
    2.372261e-06, 1.828642e-06, 8.024061e-07, 1.859351e-07, 1.710504e-07,
  2.558028e-06, 1.589662e-06, 2.056513e-06, 2.050737e-06, 4.153948e-06, 
    4.795448e-06, 6.086398e-06, 4.677413e-06, 5.318506e-06, 5.471278e-06, 
    2.702618e-06, 2.507168e-06, 1.907453e-06, 8.743522e-08, 5.300605e-08,
  9.141938e-06, 7.563072e-06, 7.763216e-06, 3.416749e-06, 4.576954e-06, 
    1.889539e-06, 2.16689e-06, 5.076333e-06, 6.095445e-06, 5.945201e-06, 
    4.007608e-06, 1.682742e-06, 1.491973e-06, 7.605752e-07, 8.250384e-08,
  1.852392e-05, 1.830183e-05, 1.721621e-05, 1.332704e-05, 8.324745e-06, 
    6.477175e-06, 1.612869e-06, 2.127661e-06, 4.59142e-06, 4.593286e-06, 
    2.976635e-06, 1.437665e-07, 2.205412e-08, 5.873448e-07, 2.527457e-07,
  2.367655e-05, 2.212014e-05, 1.776443e-05, 2.069008e-05, 1.947086e-05, 
    1.074002e-05, 1.27926e-05, 1.376854e-06, 8.181371e-07, 2.046013e-06, 
    1.195057e-06, 8.580746e-08, 9.973472e-09, 1.596534e-07, 7.087739e-08,
  2.696196e-05, 2.666415e-05, 2.238567e-05, 2.173985e-05, 2.148462e-05, 
    1.619419e-05, 1.634643e-05, 4.333019e-06, 1.836162e-06, 4.790576e-06, 
    6.573726e-07, 1.4337e-08, 5.633503e-09, 2.283632e-09, 2.073326e-09,
  3.515388e-05, 3.121447e-05, 2.318072e-05, 1.838692e-05, 1.784801e-05, 
    2.121026e-05, 1.826877e-05, 1.284254e-05, 7.944062e-06, 3.86668e-06, 
    1.965474e-06, 4.474676e-07, 1.928864e-09, 1.275504e-09, 9.323098e-10,
  3.504107e-05, 3.170142e-05, 2.609515e-05, 1.931303e-05, 1.729518e-05, 
    2.107061e-05, 2.20039e-05, 1.792671e-05, 7.369346e-06, 1.27106e-06, 
    3.496119e-07, 1.262207e-07, 5.20471e-09, 9.545341e-09, 1.00648e-08,
  3.067935e-05, 3.093492e-05, 2.887694e-05, 1.954079e-05, 1.595342e-05, 
    1.802334e-05, 1.858544e-05, 1.510136e-05, 3.206382e-06, 1.018466e-07, 
    2.497503e-08, 3.393588e-09, 7.038428e-09, 9.34663e-09, 6.292087e-08,
  2.511361e-05, 2.324422e-05, 2.274147e-05, 1.484809e-05, 1.206e-05, 
    1.287164e-05, 1.136386e-05, 5.989634e-06, 1.194798e-06, 3.214727e-07, 
    2.89878e-06, 2.508068e-07, 4.820589e-09, 5.52944e-09, 1.514979e-08,
  3.934951e-07, 6.524153e-07, 2.234211e-07, 2.490402e-06, 2.919966e-06, 
    2.019521e-06, 1.926113e-06, 1.004136e-06, 9.735878e-07, 2.806279e-07, 
    5.691753e-08, 1.121515e-06, 1.311436e-06, 2.905879e-08, 3.016254e-08,
  2.17624e-06, 1.697974e-06, 2.512345e-06, 3.217137e-07, 2.500318e-06, 
    1.971847e-06, 1.072272e-06, 1.163562e-06, 8.787337e-07, 9.577633e-07, 
    3.668963e-07, 1.746148e-06, 2.322454e-06, 6.511851e-08, 6.502736e-08,
  7.84705e-06, 5.687995e-06, 4.559824e-06, 3.074165e-06, 5.536202e-06, 
    2.004235e-06, 4.04592e-07, 1.717216e-06, 1.39425e-06, 1.087664e-06, 
    6.86765e-07, 1.053573e-06, 1.507292e-06, 9.026316e-07, 8.861392e-08,
  1.606399e-05, 1.450124e-05, 1.417532e-05, 1.277952e-05, 8.033511e-06, 
    1.367236e-05, 1.772106e-06, 1.074514e-06, 2.424573e-06, 5.944769e-07, 
    1.176258e-07, 2.723675e-07, 4.531439e-07, 1.480822e-06, 8.903053e-07,
  2.115738e-05, 1.806476e-05, 1.439847e-05, 1.406802e-05, 1.656427e-05, 
    1.286967e-05, 1.951705e-05, 1.454745e-06, 2.762176e-07, 3.018973e-07, 
    4.132153e-08, 2.397336e-08, 2.275477e-07, 6.511359e-07, 8.683891e-07,
  2.931543e-05, 2.125483e-05, 1.910811e-05, 1.7223e-05, 1.608443e-05, 
    1.89952e-05, 1.532852e-05, 7.289399e-06, 3.476653e-07, 2.358852e-06, 
    2.256171e-06, 4.453416e-07, 2.871559e-08, 7.924129e-08, 3.104552e-08,
  4.239439e-05, 4.290642e-05, 2.507352e-05, 1.837322e-05, 1.558391e-05, 
    1.451543e-05, 1.988629e-05, 8.43683e-06, 1.00753e-05, 4.554372e-06, 
    3.094627e-06, 2.928435e-07, 1.485874e-09, 4.729543e-08, 1.632183e-08,
  6.147671e-05, 5.632774e-05, 3.214338e-05, 2.206984e-05, 1.659191e-05, 
    1.522864e-05, 1.506203e-05, 1.915707e-05, 9.749261e-06, 1.820049e-06, 
    2.017071e-07, 1.459645e-07, 3.034831e-08, 1.113901e-07, 6.938789e-08,
  7.563406e-05, 5.382991e-05, 3.638635e-05, 2.306803e-05, 1.802358e-05, 
    1.257249e-05, 1.328666e-05, 1.024797e-05, 3.353842e-06, 1.392007e-06, 
    2.62087e-07, 6.272787e-07, 2.372734e-07, 2.055447e-07, 1.334594e-07,
  6.154044e-05, 4.402497e-05, 2.696583e-05, 2.39472e-05, 1.642149e-05, 
    6.159868e-06, 3.448923e-06, 3.776082e-06, 3.192862e-06, 1.88696e-06, 
    2.60605e-06, 2.69449e-06, 5.120091e-07, 1.092759e-06, 5.619226e-08,
  3.686472e-05, 2.733292e-05, 1.363675e-05, 4.560141e-06, 2.866656e-06, 
    1.184041e-06, 7.614792e-07, 5.597404e-07, 6.211265e-07, 6.142898e-08, 
    1.496363e-07, 1.727356e-07, 2.426687e-07, 1.070902e-07, 8.748647e-08,
  3.906028e-05, 2.919574e-05, 1.919998e-05, 7.50029e-06, 2.114379e-06, 
    1.489987e-06, 5.162856e-07, 2.43053e-07, 7.210308e-07, 7.037502e-07, 
    1.01088e-07, 1.117096e-06, 9.282923e-07, 8.084503e-08, 1.228752e-07,
  4.601111e-05, 3.717118e-05, 2.751089e-05, 1.282675e-05, 3.580954e-06, 
    1.25989e-06, 5.407072e-07, 4.223533e-07, 3.669296e-07, 3.866951e-07, 
    8.344631e-07, 1.934337e-07, 2.929111e-07, 6.599143e-07, 2.465422e-07,
  5.537603e-05, 4.564738e-05, 3.732232e-05, 1.829582e-05, 1.539754e-05, 
    2.033031e-06, 5.787447e-07, 4.094491e-07, 9.331018e-08, 2.583601e-08, 
    6.216057e-08, 2.118923e-07, 1.291421e-06, 1.079532e-06, 7.948938e-07,
  6.473818e-05, 5.806355e-05, 4.112702e-05, 2.62338e-05, 2.331941e-05, 
    1.276604e-05, 7.58483e-06, 4.534107e-07, 2.253688e-08, 1.424144e-09, 
    3.327331e-09, 1.170286e-07, 7.886405e-07, 1.138015e-06, 7.32434e-07,
  7.598235e-05, 7.4142e-05, 5.721115e-05, 3.497636e-05, 2.618595e-05, 
    2.290206e-05, 1.615013e-05, 6.69227e-06, 2.78449e-07, 1.220176e-06, 
    2.727195e-06, 1.184523e-06, 1.801614e-07, 6.880236e-07, 4.459478e-07,
  7.135195e-05, 8.860392e-05, 6.474989e-05, 4.768377e-05, 3.387695e-05, 
    2.207626e-05, 2.106329e-05, 1.130463e-05, 9.950125e-06, 1.854864e-06, 
    1.540732e-06, 1.091959e-08, 1.237548e-08, 5.098772e-07, 2.727248e-07,
  6.901781e-05, 8.672155e-05, 8.351902e-05, 5.343434e-05, 3.436144e-05, 
    3.063527e-05, 2.111181e-05, 2.021228e-05, 7.632048e-06, 3.295808e-06, 
    4.47746e-07, 1.674789e-07, 1.152751e-08, 2.676243e-07, 3.17143e-07,
  7.130524e-05, 9.820643e-05, 7.831037e-05, 5.447262e-05, 4.555431e-05, 
    2.77862e-05, 2.118167e-05, 1.145065e-05, 1.90642e-06, 3.047608e-06, 
    1.981309e-06, 2.081708e-06, 4.196041e-07, 3.27136e-07, 2.862672e-07,
  5.921522e-05, 6.407696e-05, 6.117031e-05, 3.616198e-05, 2.757736e-05, 
    1.666769e-05, 1.356218e-05, 1.83475e-06, 8.002511e-07, 2.039206e-06, 
    3.313122e-06, 4.314722e-06, 3.846195e-06, 1.606849e-06, 3.029924e-07,
  1.727584e-05, 1.783226e-05, 2.151484e-05, 1.766621e-05, 8.247745e-06, 
    1.5377e-06, 1.051282e-06, 9.220714e-07, 1.554286e-06, 1.062714e-06, 
    4.048704e-07, 7.868399e-07, 1.96453e-07, 1.002768e-07, 9.349038e-08,
  2.20351e-05, 2.049738e-05, 1.992336e-05, 1.761146e-05, 7.209318e-06, 
    1.574534e-06, 4.511884e-07, 5.680934e-07, 1.506001e-06, 2.161879e-06, 
    9.131718e-07, 1.397488e-06, 1.071451e-06, 8.888932e-08, 1.87324e-07,
  2.236166e-05, 2.506173e-05, 1.997754e-05, 1.754086e-05, 5.440923e-06, 
    9.418457e-07, 5.361485e-07, 1.326528e-06, 1.952712e-06, 2.79702e-06, 
    2.103157e-06, 1.191515e-06, 1.5544e-06, 5.945546e-07, 2.949643e-07,
  3.605475e-05, 3.27434e-05, 2.538863e-05, 2.365433e-05, 1.367126e-05, 
    7.889697e-07, 3.962339e-07, 7.545084e-07, 9.369029e-07, 2.15505e-06, 
    1.574619e-06, 6.823528e-07, 7.229659e-07, 1.020455e-06, 7.383022e-07,
  3.242931e-05, 3.664857e-05, 3.455882e-05, 2.964278e-05, 3.186969e-05, 
    1.533349e-05, 3.93238e-06, 1.324823e-07, 1.04793e-07, 3.44336e-07, 
    7.935907e-07, 1.023225e-06, 4.110543e-07, 9.040271e-07, 9.481369e-07,
  2.681882e-05, 5.018283e-05, 3.554521e-05, 4.811304e-05, 2.954745e-05, 
    2.11076e-05, 1.714936e-05, 1.968622e-06, 8.026054e-08, 1.698067e-06, 
    2.345081e-06, 1.764408e-06, 3.76234e-07, 4.560492e-07, 6.788222e-07,
  3.128219e-05, 5.530247e-05, 5.172516e-05, 4.173264e-05, 4.930487e-05, 
    2.958704e-05, 3.037651e-05, 1.007337e-05, 3.891791e-06, 2.066825e-06, 
    1.963652e-06, 4.632722e-07, 6.839986e-07, 4.793139e-07, 5.261955e-07,
  3.140712e-05, 4.882808e-05, 6.843861e-05, 3.361714e-05, 5.364511e-05, 
    3.89557e-05, 2.347362e-05, 2.218176e-05, 7.136221e-06, 3.095183e-07, 
    5.021635e-07, 3.805798e-07, 4.186221e-07, 5.666041e-07, 5.682443e-07,
  2.97787e-05, 4.41751e-05, 7.808138e-05, 3.566123e-05, 3.694383e-05, 
    5.154208e-05, 3.183902e-05, 2.133209e-05, 8.109664e-07, 1.923197e-07, 
    2.449694e-07, 8.835124e-07, 4.341543e-07, 4.930349e-07, 4.935568e-07,
  1.505346e-05, 2.628838e-05, 5.054371e-05, 3.035276e-05, 2.541264e-05, 
    3.408323e-05, 3.409186e-05, 9.106197e-06, 4.313129e-07, 2.886059e-07, 
    4.665609e-06, 2.611712e-06, 2.081787e-06, 3.090098e-07, 3.480739e-07,
  9.011866e-06, 1.793589e-05, 2.077088e-05, 2.263558e-05, 1.413072e-05, 
    4.156075e-06, 3.637418e-06, 2.04815e-06, 1.147807e-06, 6.105938e-07, 
    2.837343e-07, 7.971755e-07, 7.00962e-07, 3.847209e-07, 4.301484e-07,
  8.489352e-06, 1.491329e-05, 2.296259e-05, 2.77654e-05, 1.744183e-05, 
    4.993592e-06, 2.608664e-06, 1.283856e-06, 1.62824e-06, 1.742678e-06, 
    9.394223e-07, 1.267733e-06, 9.738752e-07, 6.661848e-08, 2.911068e-07,
  1.083249e-05, 1.299019e-05, 2.084839e-05, 2.845617e-05, 1.479491e-05, 
    3.486934e-06, 1.848393e-06, 2.404198e-06, 2.85022e-06, 3.285332e-06, 
    2.01258e-06, 1.57169e-06, 1.361628e-06, 6.309712e-07, 3.868558e-07,
  2.495086e-05, 2.256849e-05, 2.295624e-05, 2.804057e-05, 2.264438e-05, 
    3.024682e-06, 5.790187e-07, 1.617377e-06, 2.011133e-06, 3.226436e-06, 
    1.892884e-06, 1.18052e-06, 1.139964e-06, 1.226692e-06, 7.949953e-07,
  2.65964e-05, 2.681798e-05, 3.302272e-05, 3.020379e-05, 3.422012e-05, 
    2.125945e-05, 3.826875e-06, 1.129427e-07, 1.776686e-07, 3.225518e-07, 
    6.000564e-07, 1.060113e-06, 8.716748e-07, 1.048126e-06, 1.013789e-06,
  2.939174e-05, 3.039322e-05, 4.157834e-05, 3.505901e-05, 3.847757e-05, 
    3.110303e-05, 2.036248e-05, 3.448411e-06, 6.010942e-07, 3.407709e-06, 
    3.01777e-06, 1.488925e-06, 1.119851e-06, 8.137294e-07, 1.009279e-06,
  2.529943e-05, 2.292465e-05, 4.371961e-05, 3.980236e-05, 4.676701e-05, 
    3.140205e-05, 2.870442e-05, 1.210662e-05, 5.472923e-06, 6.111432e-06, 
    3.88523e-06, 1.321862e-06, 1.109346e-06, 7.006325e-07, 8.806687e-07,
  1.52487e-05, 1.552281e-05, 3.189369e-05, 5.586964e-05, 4.305723e-05, 
    4.191393e-05, 1.986225e-05, 1.928362e-05, 9.035795e-06, 2.7633e-06, 
    1.925863e-06, 1.142101e-06, 7.73368e-07, 6.878609e-07, 9.164867e-07,
  9.701825e-06, 1.503796e-05, 3.037109e-05, 6.073593e-05, 3.734962e-05, 
    3.971306e-05, 4.406432e-05, 2.025502e-05, 4.933118e-06, 9.353214e-08, 
    2.432108e-07, 1.093841e-06, 8.966994e-07, 9.409017e-07, 1.004302e-06,
  1.227696e-05, 2.340704e-05, 2.730312e-05, 4.57008e-05, 2.926296e-05, 
    2.603796e-05, 3.080857e-05, 9.716446e-06, 1.080989e-07, 2.023652e-07, 
    4.729926e-06, 2.057284e-06, 1.66888e-06, 1.624348e-06, 1.362701e-06,
  3.439972e-05, 3.397624e-05, 2.684644e-05, 2.280473e-05, 2.062031e-05, 
    2.033759e-05, 1.461812e-05, 1.043485e-05, 4.143083e-06, 5.538785e-07, 
    2.945768e-08, 3.956561e-07, 2.066254e-07, 1.647521e-07, 4.825998e-07,
  4.205255e-05, 3.320817e-05, 3.279222e-05, 2.67196e-05, 2.682936e-05, 
    2.59862e-05, 1.554594e-05, 1.097291e-05, 5.85083e-06, 2.18375e-06, 
    9.14774e-07, 1.150905e-06, 9.578766e-07, 2.653498e-08, 2.169097e-07,
  5.118552e-05, 3.956469e-05, 3.390251e-05, 3.208868e-05, 3.02592e-05, 
    2.640777e-05, 1.327358e-05, 8.861181e-06, 6.477785e-06, 3.759488e-06, 
    1.466129e-06, 1.283794e-06, 1.138488e-06, 7.62153e-07, 3.868608e-07,
  5.862736e-05, 5.202702e-05, 3.73052e-05, 2.982024e-05, 3.586995e-05, 
    1.828423e-05, 7.936607e-06, 3.378991e-06, 3.522752e-06, 3.61322e-06, 
    2.144294e-06, 1.040322e-06, 8.775048e-07, 1.094588e-06, 8.079011e-07,
  4.65959e-05, 5.286422e-05, 5.120499e-05, 4.041467e-05, 4.009539e-05, 
    3.241794e-05, 9.96052e-06, 1.112204e-06, 8.639267e-07, 8.309071e-07, 
    8.046028e-07, 9.128798e-07, 9.382392e-07, 8.208407e-07, 8.780677e-07,
  2.500949e-05, 4.279265e-05, 6.222274e-05, 5.937513e-05, 5.380376e-05, 
    3.592588e-05, 2.397249e-05, 3.695163e-06, 7.891102e-07, 3.072846e-06, 
    2.46654e-06, 1.450807e-06, 1.193941e-06, 7.647931e-07, 7.005365e-07,
  1.483599e-05, 2.867696e-05, 5.545914e-05, 7.618361e-05, 5.368235e-05, 
    4.23256e-05, 2.559114e-05, 1.048902e-05, 5.327532e-06, 7.509484e-06, 
    3.989585e-06, 1.922968e-06, 1.292183e-06, 6.773727e-07, 4.107363e-07,
  2.681781e-05, 3.750298e-05, 5.957041e-05, 7.313056e-05, 4.638968e-05, 
    3.764127e-05, 2.868476e-05, 1.215743e-05, 6.26225e-06, 4.906891e-06, 
    2.115077e-06, 1.72745e-06, 1.313342e-06, 6.217955e-07, 2.807333e-07,
  3.409578e-05, 4.470529e-05, 6.006728e-05, 5.937005e-05, 3.856579e-05, 
    3.13372e-05, 3.123286e-05, 1.559247e-05, 2.33431e-06, 4.332318e-08, 
    8.337719e-08, 1.344109e-06, 1.064435e-06, 5.713242e-07, 2.889131e-07,
  2.877379e-05, 2.949757e-05, 4.626719e-05, 3.395131e-05, 3.079095e-05, 
    2.480513e-05, 2.192289e-05, 9.878159e-06, 3.808024e-07, 1.140714e-07, 
    3.968062e-06, 1.638429e-06, 1.525093e-06, 1.300395e-06, 1.261077e-06,
  3.489617e-05, 3.76153e-05, 3.64857e-05, 4.214638e-05, 3.955129e-05, 
    3.220703e-05, 2.483277e-05, 2.028901e-05, 1.759011e-05, 1.334821e-05, 
    7.723666e-06, 4.607462e-06, 2.078176e-06, 7.702874e-07, 2.244778e-06,
  4.938705e-05, 3.365944e-05, 3.632316e-05, 3.885182e-05, 3.751439e-05, 
    3.01804e-05, 2.631177e-05, 2.342472e-05, 1.874908e-05, 1.569845e-05, 
    8.212217e-06, 4.613676e-06, 1.434909e-06, 1.70415e-07, 8.029832e-07,
  3.48266e-05, 1.927679e-05, 2.25842e-05, 2.436517e-05, 2.40804e-05, 
    1.855825e-05, 2.596744e-05, 2.783251e-05, 2.232192e-05, 1.814861e-05, 
    8.73673e-06, 3.942042e-06, 1.342691e-06, 1.854465e-07, 3.111084e-07,
  2.054638e-05, 2.139738e-05, 2.390952e-05, 2.345662e-05, 2.521404e-05, 
    1.294438e-05, 1.572842e-05, 1.35932e-05, 1.315301e-05, 1.378168e-05, 
    8.211482e-06, 2.040712e-06, 3.860051e-07, 2.08223e-07, 1.70478e-07,
  2.562251e-05, 2.236375e-05, 3.402064e-05, 3.666865e-05, 2.771881e-05, 
    2.454395e-05, 1.025637e-05, 1.539959e-06, 1.597272e-06, 5.919272e-06, 
    5.022483e-06, 6.332379e-07, 1.283055e-07, 1.028282e-07, 1.211856e-07,
  2.428652e-05, 2.78834e-05, 3.906164e-05, 4.862956e-05, 3.999077e-05, 
    3.487193e-05, 2.06227e-05, 4.739618e-06, 4.375791e-06, 9.755244e-06, 
    5.667634e-06, 2.032888e-06, 6.817284e-07, 5.506618e-08, 6.617213e-08,
  1.588411e-05, 2.451831e-05, 6.551806e-05, 4.307999e-05, 4.267272e-05, 
    3.978976e-05, 3.008568e-05, 1.038271e-05, 1.032227e-05, 1.203132e-05, 
    8.092633e-06, 2.483627e-06, 8.451972e-07, 3.799842e-08, 4.362499e-09,
  2.461108e-05, 3.808535e-05, 6.015057e-05, 5.069119e-05, 4.737731e-05, 
    4.009156e-05, 2.354779e-05, 1.590921e-05, 8.01531e-06, 4.875297e-06, 
    3.281822e-06, 1.843857e-06, 4.592706e-07, 1.241687e-07, 3.542796e-08,
  6.680486e-05, 7.180852e-05, 8.518304e-05, 6.108966e-05, 4.781898e-05, 
    3.368383e-05, 1.934181e-05, 1.567175e-05, 1.85009e-06, 1.522786e-06, 
    1.286063e-06, 1.25735e-06, 8.388487e-07, 4.353774e-07, 1.473516e-07,
  4.943025e-05, 4.836696e-05, 4.701743e-05, 3.97577e-05, 3.565191e-05, 
    3.298939e-05, 1.39644e-05, 9.618408e-06, 3.109581e-06, 1.240445e-06, 
    5.317542e-06, 2.280449e-06, 1.65508e-06, 9.791851e-07, 5.215867e-07,
  1.406451e-05, 1.109358e-05, 1.132208e-05, 1.183235e-05, 1.135346e-05, 
    1.321232e-05, 1.220186e-05, 1.205615e-05, 1.082208e-05, 8.041744e-06, 
    8.592227e-06, 1.28508e-05, 1.62025e-05, 1.655742e-05, 1.624797e-05,
  2.47321e-05, 1.840508e-05, 2.340351e-05, 2.801609e-05, 2.576329e-05, 
    1.364234e-05, 9.737825e-06, 1.244401e-05, 9.844811e-06, 1.057979e-05, 
    1.200492e-05, 1.405387e-05, 1.293133e-05, 8.445063e-06, 1.003183e-05,
  2.123641e-05, 1.292402e-05, 2.71319e-05, 4.069007e-05, 3.450618e-05, 
    1.312558e-05, 1.501109e-05, 2.471553e-05, 1.301798e-05, 8.915944e-06, 
    1.063845e-05, 1.127804e-05, 1.082102e-05, 8.649772e-06, 7.484937e-06,
  1.812652e-05, 1.857316e-05, 2.40834e-05, 2.142298e-05, 3.62408e-05, 
    2.446789e-05, 2.570682e-05, 2.208178e-05, 7.597278e-06, 6.447975e-06, 
    9.0437e-06, 8.554561e-06, 8.48986e-06, 7.41965e-06, 4.173972e-06,
  2.365997e-05, 2.17471e-05, 2.32396e-05, 3.059255e-05, 2.845824e-05, 
    5.389034e-05, 2.960989e-05, 1.125112e-05, 4.18922e-06, 6.943175e-06, 
    8.746532e-06, 6.344747e-06, 5.932595e-06, 2.923701e-06, 1.790649e-06,
  1.831407e-05, 1.90504e-05, 2.241578e-05, 3.864246e-05, 6.308366e-05, 
    4.765758e-05, 2.979364e-05, 1.011425e-05, 5.777769e-06, 8.174936e-06, 
    6.479737e-06, 6.698757e-06, 5.039654e-06, 2.524303e-06, 6.201022e-07,
  2.100928e-05, 3.096402e-05, 4.84101e-05, 7.972237e-05, 5.030916e-05, 
    3.05408e-05, 2.260294e-05, 1.211199e-05, 8.089026e-06, 1.140052e-05, 
    1.112606e-05, 8.535675e-06, 4.532767e-06, 1.954024e-06, 1.810541e-08,
  2.070288e-05, 2.997324e-05, 4.435879e-05, 3.64572e-05, 3.300522e-05, 
    2.350392e-05, 2.041471e-05, 1.436458e-05, 6.440078e-06, 5.023591e-06, 
    9.011676e-06, 7.629958e-06, 3.330706e-06, 1.120391e-06, 9.677117e-09,
  2.973454e-05, 2.526979e-05, 2.859136e-05, 3.118788e-05, 2.204823e-05, 
    2.143289e-05, 1.993034e-05, 1.358394e-05, 1.430732e-06, 1.888889e-06, 
    4.514154e-06, 4.771494e-06, 2.395519e-06, 3.465383e-07, 2.179551e-07,
  2.654372e-05, 3.056698e-05, 3.305851e-05, 3.377455e-05, 3.195368e-05, 
    2.00747e-05, 1.116953e-05, 7.332625e-06, 2.527977e-06, 1.47781e-06, 
    5.32051e-06, 4.285611e-06, 2.070791e-06, 3.210569e-07, 2.85799e-07,
  3.702089e-06, 5.316386e-06, 8.134696e-06, 9.880708e-06, 7.71784e-06, 
    8.378558e-06, 6.056211e-06, 3.094808e-06, 1.87618e-06, 1.442737e-06, 
    1.252986e-06, 3.730044e-06, 6.585742e-06, 7.173988e-06, 8.781169e-06,
  5.491135e-07, 1.297026e-06, 3.645077e-06, 9.370394e-06, 1.434763e-05, 
    1.302154e-05, 9.565899e-06, 6.345537e-06, 3.138733e-06, 2.712168e-06, 
    2.861397e-06, 4.542607e-06, 5.935146e-06, 4.643411e-06, 9.436762e-06,
  7.501195e-06, 4.1526e-06, 1.261207e-06, 3.51954e-06, 1.120214e-05, 
    1.830454e-05, 1.591342e-05, 2.120201e-05, 1.039518e-05, 5.051635e-06, 
    4.566521e-06, 6.242083e-06, 7.528526e-06, 8.074334e-06, 1.118539e-05,
  9.532765e-06, 1.519606e-05, 2.033014e-05, 1.195482e-05, 6.602255e-06, 
    1.76656e-05, 2.815549e-05, 2.05478e-05, 7.683001e-06, 5.195987e-06, 
    6.703314e-06, 6.506468e-06, 7.03689e-06, 8.66882e-06, 8.450774e-06,
  1.051666e-05, 1.502439e-05, 1.770276e-05, 2.006637e-05, 1.093982e-05, 
    3.022703e-05, 3.484886e-05, 1.196552e-05, 3.067248e-06, 8.290608e-06, 
    1.209116e-05, 5.799917e-06, 6.121054e-06, 4.724157e-06, 5.633834e-06,
  1.243222e-05, 1.830521e-05, 1.947173e-05, 2.839124e-05, 2.952539e-05, 
    3.771895e-05, 3.798479e-05, 1.81028e-05, 1.619271e-05, 1.801281e-05, 
    1.357307e-05, 8.645372e-06, 6.685264e-06, 4.34907e-06, 3.475976e-06,
  1.147816e-05, 1.917309e-05, 2.489706e-05, 2.315261e-05, 3.020949e-05, 
    2.570678e-05, 2.454752e-05, 1.456551e-05, 1.121658e-05, 1.44736e-05, 
    1.764078e-05, 1.524612e-05, 8.505617e-06, 4.86495e-06, 2.685023e-06,
  8.670674e-06, 1.35259e-05, 1.824345e-05, 2.02683e-05, 2.216991e-05, 
    2.570376e-05, 2.125676e-05, 1.499697e-05, 3.63184e-06, 8.663346e-06, 
    1.813621e-05, 1.932859e-05, 1.221384e-05, 6.789165e-06, 2.288173e-06,
  8.572915e-06, 1.35397e-05, 1.932437e-05, 2.183153e-05, 2.198497e-05, 
    1.96532e-05, 2.175673e-05, 1.041424e-05, 2.117773e-06, 4.249642e-06, 
    1.2229e-05, 1.682965e-05, 1.508828e-05, 7.77727e-06, 2.064816e-06,
  6.384933e-06, 7.575529e-06, 9.064763e-06, 1.372657e-05, 1.58603e-05, 
    1.402123e-05, 1.35477e-05, 6.030598e-06, 5.063089e-07, 1.367403e-06, 
    7.968646e-06, 1.318931e-05, 1.324243e-05, 7.464216e-06, 1.803955e-06,
  8.289644e-07, 7.007809e-07, 6.888297e-07, 1.615258e-06, 5.666602e-06, 
    8.036859e-06, 6.879828e-06, 5.436042e-06, 7.580825e-06, 7.099869e-06, 
    6.588001e-06, 1.27537e-05, 1.859074e-05, 1.840098e-05, 1.858907e-05,
  1.616263e-06, 8.272864e-07, 1.814098e-07, 6.34089e-07, 3.42037e-06, 
    3.88218e-06, 7.966351e-06, 8.293431e-06, 6.721066e-06, 6.738658e-06, 
    7.115314e-06, 9.549673e-06, 1.168925e-05, 1.10303e-05, 1.483263e-05,
  5.264164e-06, 1.407364e-06, 1.571957e-06, 6.180837e-07, 2.678555e-06, 
    6.83841e-06, 3.898973e-06, 8.143034e-06, 9.400233e-06, 6.307909e-06, 
    9.64041e-06, 8.25882e-06, 8.784646e-06, 1.113661e-05, 1.20989e-05,
  4.482179e-06, 5.934816e-06, 1.203102e-05, 1.073086e-05, 3.782816e-06, 
    5.235527e-06, 8.451763e-06, 5.188392e-06, 5.922101e-06, 9.711183e-06, 
    9.935281e-06, 8.179031e-06, 8.676204e-06, 1.025675e-05, 8.409771e-06,
  5.189285e-06, 3.133978e-06, 7.934519e-06, 1.394247e-05, 1.68763e-05, 
    1.044989e-05, 7.225355e-06, 3.682685e-06, 7.284091e-06, 9.561639e-06, 
    1.208672e-05, 9.404761e-06, 1.006637e-05, 7.937929e-06, 7.326594e-06,
  6.465806e-06, 1.926752e-06, 6.110867e-06, 1.184229e-05, 2.19456e-05, 
    2.13057e-05, 1.470221e-05, 8.452249e-06, 4.949762e-06, 7.644197e-06, 
    1.045898e-05, 1.16133e-05, 1.130219e-05, 7.859155e-06, 7.039637e-06,
  5.032562e-06, 8.666032e-07, 4.619363e-06, 1.524816e-05, 2.731483e-05, 
    2.73635e-05, 1.790781e-05, 9.307273e-06, 4.098586e-06, 4.397996e-06, 
    9.264057e-06, 1.281051e-05, 1.027744e-05, 7.329088e-06, 5.591999e-06,
  1.543892e-06, 4.406258e-07, 5.446673e-06, 2.549504e-05, 2.699219e-05, 
    2.541678e-05, 2.021176e-05, 1.338456e-05, 3.306794e-06, 1.589081e-06, 
    6.699666e-06, 1.168189e-05, 1.049995e-05, 6.630195e-06, 4.514463e-06,
  4.509641e-08, 1.994129e-06, 2.672062e-05, 2.990481e-05, 2.320801e-05, 
    2.24842e-05, 2.220149e-05, 1.218231e-05, 9.086611e-07, 9.100586e-07, 
    4.877825e-06, 1.257866e-05, 1.07143e-05, 6.391929e-06, 3.92431e-06,
  1.392881e-06, 9.823711e-06, 3.464685e-05, 2.867158e-05, 1.883768e-05, 
    1.836418e-05, 1.791954e-05, 9.746563e-06, 7.073533e-07, 9.153269e-07, 
    4.108676e-06, 1.261236e-05, 1.459621e-05, 6.995367e-06, 3.426071e-06,
  2.220159e-07, 9.962987e-09, 1.078995e-06, 1.702152e-07, 1.624054e-07, 
    4.956371e-06, 9.950752e-06, 9.833201e-06, 1.144849e-05, 1.245333e-05, 
    1.06143e-05, 7.033677e-06, 5.96899e-06, 8.989075e-06, 1.163649e-05,
  1.998692e-07, 5.283034e-07, 2.531892e-07, 6.669298e-08, 8.71907e-07, 
    6.06555e-06, 8.207062e-06, 1.095042e-05, 1.442474e-05, 1.167142e-05, 
    9.168855e-06, 6.515394e-06, 5.329205e-06, 7.341366e-06, 1.052793e-05,
  2.555571e-06, 2.120239e-06, 3.229511e-07, 4.010183e-07, 4.71204e-06, 
    1.915889e-05, 1.430923e-05, 1.639514e-05, 2.075566e-05, 1.350837e-05, 
    5.539191e-06, 3.82291e-06, 4.420071e-06, 6.518093e-06, 9.31973e-06,
  8.872266e-06, 3.014391e-06, 5.691183e-06, 8.124619e-06, 2.19815e-05, 
    4.193878e-05, 6.437553e-05, 3.129306e-05, 2.290476e-05, 1.470651e-05, 
    5.254887e-06, 2.648723e-06, 3.594505e-06, 3.782092e-06, 6.184581e-06,
  8.701762e-06, 2.521491e-06, 1.108294e-05, 2.789657e-05, 3.922057e-05, 
    6.04499e-05, 7.471373e-05, 7.350511e-05, 2.497858e-05, 1.116605e-05, 
    5.247013e-06, 2.459394e-06, 2.937269e-06, 2.937628e-06, 4.181695e-06,
  1.013314e-05, 1.205645e-05, 2.909222e-05, 4.553007e-05, 6.344027e-05, 
    6.634876e-05, 6.02891e-05, 3.286357e-05, 9.586854e-06, 4.772727e-06, 
    3.000034e-06, 2.651104e-06, 3.375197e-06, 4.229985e-06, 4.278144e-06,
  8.53138e-06, 2.453381e-05, 4.030217e-05, 5.719629e-05, 6.132155e-05, 
    5.365003e-05, 3.464637e-05, 1.07376e-05, 8.488998e-06, 6.08112e-06, 
    7.752091e-07, 1.804819e-06, 2.366471e-06, 5.652723e-06, 6.059721e-06,
  9.320142e-06, 3.219198e-05, 5.002724e-05, 7.214243e-05, 5.520819e-05, 
    3.62847e-05, 1.815911e-05, 1.231918e-05, 1.011096e-05, 6.388157e-06, 
    4.899663e-07, 4.549615e-07, 2.435181e-06, 5.608891e-06, 6.049672e-06,
  2.082663e-05, 4.797346e-05, 7.172948e-05, 6.336974e-05, 3.825034e-05, 
    2.483939e-05, 1.618033e-05, 8.405081e-06, 8.989292e-06, 3.723625e-06, 
    3.621409e-07, 4.538068e-07, 2.722681e-06, 5.277758e-06, 6.109025e-06,
  1.259752e-05, 4.447536e-05, 6.461157e-05, 3.842339e-05, 2.99312e-05, 
    1.549117e-05, 1.161401e-05, 5.111019e-06, 7.701544e-06, 3.149441e-06, 
    2.786404e-07, 5.794819e-07, 3.596968e-06, 5.539459e-06, 6.128178e-06,
  9.103151e-09, 3.006169e-08, 3.624728e-07, 2.331765e-06, 1.480528e-05, 
    2.823537e-05, 3.443325e-05, 3.335945e-05, 2.458758e-05, 1.432006e-05, 
    1.383314e-05, 2.436355e-05, 3.888299e-05, 3.647128e-05, 2.484101e-05,
  8.253664e-08, 5.902563e-07, 1.352691e-06, 1.186848e-05, 2.749601e-05, 
    3.389488e-05, 3.529957e-05, 3.02077e-05, 1.836705e-05, 1.251079e-05, 
    1.553272e-05, 3.552154e-05, 4.018565e-05, 2.771713e-05, 1.989628e-05,
  1.825735e-06, 3.662918e-06, 8.6978e-06, 2.784856e-05, 4.640118e-05, 
    4.667748e-05, 1.806248e-05, 9.482486e-06, 1.010845e-05, 1.276471e-05, 
    1.90433e-05, 3.308578e-05, 2.516349e-05, 1.577658e-05, 1.10355e-05,
  6.477885e-06, 9.1332e-06, 2.450744e-05, 3.955951e-05, 3.831352e-05, 
    2.423264e-05, 8.379351e-06, 8.105015e-07, 3.150469e-06, 1.52141e-05, 
    2.217358e-05, 1.346944e-05, 9.664843e-06, 8.505643e-06, 4.023127e-06,
  7.504396e-06, 1.259823e-05, 2.570375e-05, 2.772193e-05, 1.745269e-05, 
    8.337417e-06, 9.013831e-07, 4.565653e-06, 1.223369e-05, 1.217714e-05, 
    1.112661e-05, 3.728944e-06, 3.292245e-06, 6.051499e-06, 3.988021e-06,
  8.311964e-06, 1.208483e-05, 1.478451e-05, 1.250235e-05, 1.339184e-05, 
    1.11384e-05, 1.006156e-05, 5.98938e-06, 7.560522e-06, 4.618983e-06, 
    1.69549e-06, 3.78406e-06, 4.138778e-06, 2.690395e-06, 2.523497e-06,
  1.280033e-05, 1.177401e-05, 8.830548e-06, 9.371782e-06, 1.131046e-05, 
    1.258436e-05, 1.668327e-05, 1.093664e-05, 7.339535e-06, 3.045266e-06, 
    1.301797e-06, 2.035781e-06, 4.396074e-06, 2.428345e-06, 2.178498e-06,
  1.298553e-05, 1.111667e-05, 9.631355e-06, 6.564061e-06, 1.389128e-05, 
    1.250935e-05, 1.93537e-05, 2.165386e-05, 1.476224e-05, 7.023774e-06, 
    1.653341e-06, 1.526268e-06, 2.767335e-07, 1.425867e-06, 1.469566e-06,
  1.244257e-05, 9.312165e-06, 1.042935e-05, 4.072294e-06, 6.966881e-06, 
    1.310316e-05, 2.079944e-05, 2.999415e-05, 2.858485e-05, 1.598845e-05, 
    3.848954e-06, 1.57523e-07, 1.192964e-07, 8.706759e-07, 1.426598e-06,
  4.098054e-06, 1.350621e-06, 3.770014e-06, 2.215678e-06, 4.11388e-06, 
    1.134369e-05, 2.075708e-05, 3.230749e-05, 4.208825e-05, 3.489195e-05, 
    1.112414e-05, 9.351494e-07, 7.192879e-08, 7.441059e-07, 1.386478e-06,
  3.136083e-07, 4.36748e-08, 1.123629e-06, 4.831843e-08, 1.361153e-06, 
    2.511899e-06, 4.617649e-06, 1.772212e-05, 1.70348e-05, 3.321075e-06, 
    1.759764e-06, 3.766545e-06, 8.472547e-06, 9.110274e-06, 1.037367e-05,
  3.610735e-07, 1.978539e-08, 2.049245e-08, 1.184164e-06, 2.504539e-06, 
    1.751202e-06, 5.930091e-06, 2.6387e-05, 2.437749e-05, 4.628578e-06, 
    7.527083e-07, 2.129902e-06, 3.567428e-06, 3.405366e-06, 5.395387e-06,
  1.645386e-06, 3.423919e-08, 1.085683e-06, 3.161858e-06, 3.269787e-06, 
    3.553182e-06, 5.994488e-06, 2.948733e-05, 4.029698e-05, 1.203333e-05, 
    1.166112e-06, 3.533545e-07, 8.537708e-07, 2.786932e-06, 2.850941e-06,
  5.616435e-06, 4.849217e-06, 5.915319e-06, 6.983494e-06, 4.299879e-06, 
    2.54512e-06, 1.350179e-05, 1.319488e-05, 2.359855e-05, 2.761132e-05, 
    3.31081e-06, 1.671996e-06, 1.718781e-07, 6.945857e-07, 1.422378e-06,
  1.103956e-05, 7.938179e-06, 7.403465e-06, 1.047274e-05, 7.778284e-06, 
    4.783901e-06, 9.445932e-06, 4.22807e-05, 7.050742e-05, 4.689557e-05, 
    1.366547e-05, 2.687279e-06, 1.659396e-06, 8.921779e-07, 2.652908e-06,
  9.666919e-06, 6.285429e-06, 5.762002e-06, 7.253442e-06, 1.319805e-05, 
    8.687037e-06, 1.203526e-05, 2.375715e-05, 4.751861e-05, 6.43372e-05, 
    2.992956e-05, 6.29281e-06, 7.363496e-07, 7.719977e-07, 2.652049e-07,
  1.291634e-05, 6.832656e-06, 5.61222e-06, 3.45776e-06, 1.050025e-05, 
    8.80537e-06, 1.258555e-05, 2.282569e-05, 4.602762e-05, 5.408252e-05, 
    4.389939e-05, 1.520232e-05, 2.279292e-06, 1.397257e-07, 1.255042e-08,
  1.125615e-05, 5.042686e-06, 3.83943e-06, 2.499133e-06, 8.268416e-06, 
    2.511463e-06, 6.258192e-06, 9.448077e-06, 2.892392e-05, 4.962902e-05, 
    5.160133e-05, 2.475426e-05, 7.540863e-06, 1.530209e-06, 1.517251e-07,
  9.146428e-06, 4.767401e-06, 6.862194e-06, 3.692609e-06, 2.978913e-06, 
    7.994743e-07, 2.981452e-06, 6.310661e-06, 1.898384e-05, 4.280595e-05, 
    4.735558e-05, 3.007516e-05, 1.342045e-05, 3.608221e-06, 4.000964e-07,
  2.872244e-06, 2.254556e-06, 3.771516e-06, 2.982839e-06, 1.366918e-06, 
    3.91797e-07, 1.348262e-06, 4.737565e-06, 1.139685e-05, 3.785559e-05, 
    4.830309e-05, 3.516272e-05, 1.568882e-05, 6.922751e-06, 1.400895e-06,
  5.43162e-06, 4.53087e-07, 1.829019e-06, 1.511549e-06, 3.310053e-06, 
    3.53077e-06, 3.303739e-06, 2.332888e-06, 1.583588e-06, 5.862355e-07, 
    7.961636e-07, 8.909325e-07, 6.417694e-07, 8.469675e-07, 1.238395e-06,
  1.80418e-06, 7.212079e-07, 2.164482e-06, 8.936128e-07, 2.333845e-06, 
    1.946686e-06, 1.358514e-06, 1.377732e-06, 3.993222e-06, 1.452955e-06, 
    7.794916e-07, 1.671092e-06, 1.459907e-06, 7.060956e-07, 1.180569e-06,
  1.443278e-06, 1.086436e-05, 3.280293e-06, 2.306007e-06, 1.819908e-06, 
    4.98378e-06, 4.589315e-07, 2.046529e-06, 5.113882e-06, 6.311802e-06, 
    2.125727e-06, 8.398129e-07, 7.335757e-07, 2.489921e-06, 1.801225e-06,
  7.377897e-06, 2.100001e-05, 1.156159e-05, 1.003322e-05, 5.270091e-06, 
    2.436779e-06, 2.43077e-06, 2.61154e-06, 3.987415e-06, 1.176777e-05, 
    7.254119e-06, 2.221338e-06, 1.757653e-07, 1.135268e-06, 2.075314e-06,
  1.457415e-05, 1.27813e-05, 1.234659e-05, 1.020064e-05, 9.061151e-06, 
    6.931661e-06, 3.924995e-06, 1.194374e-05, 2.39942e-05, 1.374913e-05, 
    1.440314e-05, 8.983438e-06, 2.177754e-06, 3.872221e-07, 2.223245e-07,
  2.041478e-05, 1.157937e-05, 1.098081e-05, 8.521866e-06, 9.062239e-06, 
    1.076616e-05, 8.23723e-06, 6.603816e-06, 6.967476e-06, 8.030245e-06, 
    1.315227e-05, 1.11308e-05, 6.71714e-06, 2.507977e-06, 1.154066e-06,
  1.115361e-05, 9.157489e-06, 8.648502e-06, 5.935877e-06, 8.922526e-06, 
    1.069046e-05, 1.314843e-05, 9.563917e-06, 8.825115e-06, 7.855914e-06, 
    1.013591e-05, 9.838822e-06, 8.425873e-06, 4.045454e-06, 2.416526e-06,
  1.114412e-05, 7.456606e-06, 5.072513e-06, 2.715633e-06, 6.688608e-06, 
    8.360802e-06, 8.330771e-06, 8.135973e-06, 9.476177e-06, 7.909855e-06, 
    8.22871e-06, 8.239339e-06, 8.001903e-06, 6.539075e-06, 3.7467e-06,
  1.031732e-05, 1.018037e-05, 6.647133e-06, 4.811503e-06, 4.77377e-06, 
    6.781916e-06, 7.6956e-06, 5.693767e-06, 6.990095e-06, 6.439692e-06, 
    5.653622e-06, 6.46086e-06, 6.611536e-06, 6.770356e-06, 6.577907e-06,
  7.481814e-06, 3.257478e-06, 2.313796e-06, 2.045518e-06, 4.253384e-06, 
    5.024192e-06, 5.550867e-06, 3.391972e-06, 3.168517e-06, 3.381658e-06, 
    3.969048e-06, 4.108098e-06, 4.705422e-06, 6.540973e-06, 7.487288e-06,
  5.981321e-06, 6.948021e-07, 1.114121e-06, 2.498622e-07, 4.662008e-07, 
    8.280001e-07, 2.729798e-06, 5.41349e-06, 5.702573e-06, 2.852047e-06, 
    1.691639e-06, 1.467793e-06, 1.203987e-06, 1.228763e-06, 1.639641e-06,
  1.382994e-06, 1.585203e-06, 3.747993e-07, 9.418427e-08, 3.10572e-07, 
    1.347702e-06, 2.19812e-06, 3.396134e-06, 4.000971e-06, 4.98609e-06, 
    1.894154e-06, 2.258894e-06, 2.33891e-06, 2.967754e-06, 2.678454e-06,
  1.302903e-05, 1.084788e-05, 7.540336e-07, 9.474717e-08, 1.681247e-07, 
    1.082542e-06, 9.925232e-07, 2.7118e-06, 4.077122e-06, 4.984808e-06, 
    5.309566e-06, 5.250402e-06, 4.054824e-06, 3.47583e-06, 4.243256e-06,
  1.675573e-05, 1.624859e-05, 1.488246e-05, 7.798611e-06, 7.824999e-07, 
    9.237692e-07, 3.370505e-06, 1.839397e-06, 3.469034e-06, 5.265322e-06, 
    6.732447e-06, 8.57031e-06, 9.418284e-06, 1.005973e-05, 1.065313e-05,
  1.365596e-05, 1.203704e-05, 1.116285e-05, 9.207786e-06, 9.087644e-06, 
    6.904885e-06, 4.313001e-06, 9.165409e-06, 7.223346e-06, 4.96443e-06, 
    1.191711e-05, 1.366836e-05, 1.760404e-05, 2.069319e-05, 2.22523e-05,
  9.861689e-06, 8.005465e-06, 6.863038e-06, 8.413298e-06, 9.607954e-06, 
    5.384192e-06, 6.54395e-06, 8.237545e-06, 1.568175e-05, 2.247923e-05, 
    2.774575e-05, 2.831835e-05, 3.063422e-05, 3.474173e-05, 3.630744e-05,
  5.041693e-06, 7.277337e-06, 9.064072e-06, 6.424777e-06, 6.656059e-06, 
    5.963632e-06, 8.301714e-06, 1.861717e-05, 3.265906e-05, 3.125618e-05, 
    3.212578e-05, 3.524614e-05, 3.910042e-05, 4.064905e-05, 3.595277e-05,
  4.990898e-06, 6.863751e-06, 6.548036e-06, 2.419575e-06, 3.595575e-06, 
    5.325363e-06, 1.017482e-05, 2.039777e-05, 3.044615e-05, 3.622803e-05, 
    3.977385e-05, 4.140881e-05, 4.26409e-05, 4.232711e-05, 3.651512e-05,
  4.283218e-06, 4.290524e-06, 4.678221e-06, 4.790177e-06, 7.79253e-06, 
    1.101172e-05, 1.247264e-05, 1.896155e-05, 3.152972e-05, 3.466142e-05, 
    3.166043e-05, 3.326069e-05, 3.794338e-05, 4.174203e-05, 4.118079e-05,
  2.182552e-06, 4.169981e-06, 8.991585e-06, 1.801752e-05, 2.593175e-05, 
    2.593871e-05, 1.855103e-05, 2.17878e-05, 3.346959e-05, 3.779163e-05, 
    3.76522e-05, 4.085355e-05, 4.615076e-05, 4.913911e-05, 4.655766e-05,
  3.563034e-06, 3.974244e-06, 2.260103e-06, 4.259969e-07, 7.640682e-08, 
    1.222187e-07, 1.365549e-07, 4.636722e-07, 1.165042e-06, 2.805366e-06, 
    5.432577e-06, 1.279287e-05, 2.292187e-05, 2.847344e-05, 3.260748e-05,
  7.277794e-06, 3.852615e-06, 2.801604e-06, 4.368831e-07, 1.117547e-06, 
    1.493607e-07, 8.849337e-08, 2.063577e-07, 7.139902e-07, 2.548505e-06, 
    6.550359e-06, 1.659869e-05, 3.022136e-05, 4.3868e-05, 4.35654e-05,
  7.0109e-06, 6.042768e-06, 4.664692e-06, 1.72401e-06, 2.487013e-06, 
    1.165444e-06, 4.999892e-08, 5.081504e-07, 3.302091e-06, 1.184349e-05, 
    1.725673e-05, 2.173995e-05, 3.164302e-05, 4.004495e-05, 5.42499e-05,
  7.27919e-06, 6.008964e-06, 5.165936e-06, 3.810994e-06, 2.738492e-06, 
    8.317819e-07, 1.728456e-06, 8.911722e-07, 4.294864e-06, 1.51637e-05, 
    2.824302e-05, 2.521682e-05, 2.707565e-05, 3.250225e-05, 4.960516e-05,
  9.662532e-06, 5.882052e-06, 5.387394e-06, 3.930629e-06, 4.635594e-06, 
    3.749562e-06, 9.710576e-07, 8.956865e-06, 5.140247e-06, 7.279932e-06, 
    2.000816e-05, 1.981949e-05, 2.012622e-05, 2.156639e-05, 3.065107e-05,
  2.046303e-05, 9.940803e-06, 5.668974e-06, 3.75678e-06, 3.223375e-06, 
    2.727303e-06, 2.075514e-06, 4.32789e-06, 1.403911e-05, 1.966437e-05, 
    1.663313e-05, 1.298786e-05, 1.158603e-05, 1.249194e-05, 1.703436e-05,
  2.284935e-05, 1.694077e-05, 8.398665e-06, 5.007224e-06, 2.361965e-06, 
    1.786195e-06, 2.507406e-06, 8.233796e-06, 2.054578e-05, 1.239387e-05, 
    4.73454e-06, 3.719329e-06, 3.424817e-06, 4.56272e-06, 6.796795e-06,
  2.067193e-05, 1.537942e-05, 8.00352e-06, 4.590871e-06, 1.69864e-06, 
    1.925428e-06, 5.625437e-06, 1.489116e-05, 1.175363e-05, 5.219465e-06, 
    2.137026e-06, 1.444478e-06, 1.555089e-06, 1.932302e-06, 4.439916e-06,
  1.63178e-05, 1.218995e-05, 7.775515e-06, 4.84931e-06, 3.940135e-06, 
    5.598866e-06, 1.766371e-05, 1.599458e-05, 9.024575e-06, 3.685598e-06, 
    1.970203e-06, 6.753179e-07, 7.333138e-07, 1.502487e-06, 6.254442e-06,
  1.24938e-05, 7.632641e-06, 5.809557e-06, 5.050472e-06, 6.74684e-06, 
    1.659516e-05, 1.952463e-05, 1.184554e-05, 8.905676e-06, 3.159764e-06, 
    2.965948e-06, 3.775429e-07, 6.904727e-07, 3.669631e-06, 1.447341e-05,
  5.33387e-06, 3.71014e-06, 6.078503e-06, 6.3353e-06, 4.491275e-06, 
    3.411763e-06, 2.411645e-06, 8.322525e-07, 3.965886e-07, 3.592548e-07, 
    1.90834e-07, 1.054763e-06, 2.601449e-06, 1.705538e-06, 2.188187e-06,
  8.592951e-06, 6.591795e-06, 6.561503e-06, 6.378342e-06, 5.599831e-06, 
    3.963729e-06, 3.319368e-06, 1.435075e-06, 6.242867e-07, 3.717214e-07, 
    3.677501e-07, 1.402955e-06, 2.043462e-06, 2.624488e-06, 2.513468e-06,
  1.428433e-05, 1.106095e-05, 9.224145e-06, 9.361261e-06, 8.674685e-06, 
    6.363687e-06, 2.428886e-06, 2.439404e-06, 2.016972e-06, 1.344153e-06, 
    1.053694e-06, 2.410805e-06, 2.423831e-06, 2.492203e-06, 3.411199e-06,
  1.737762e-05, 2.127654e-05, 2.247908e-05, 1.895879e-05, 1.82999e-05, 
    8.576911e-06, 8.504107e-06, 2.356872e-06, 7.614999e-07, 5.558351e-07, 
    2.100157e-06, 2.736383e-06, 4.068543e-06, 5.50397e-06, 6.972972e-06,
  1.745599e-05, 2.241989e-05, 2.517188e-05, 2.838702e-05, 2.75827e-05, 
    1.871857e-05, 1.814261e-05, 1.374698e-05, 1.350368e-06, 2.411807e-06, 
    4.831918e-06, 5.032079e-06, 7.769529e-06, 1.049216e-05, 1.292547e-05,
  1.907644e-05, 2.115146e-05, 2.349561e-05, 2.569381e-05, 2.763707e-05, 
    2.579832e-05, 2.46279e-05, 1.248257e-05, 5.389917e-06, 6.909037e-06, 
    1.121319e-05, 1.22035e-05, 1.56414e-05, 1.72352e-05, 1.964158e-05,
  1.992592e-05, 2.638543e-05, 2.541506e-05, 2.153262e-05, 2.066399e-05, 
    1.976275e-05, 1.856636e-05, 1.106818e-05, 4.624759e-06, 5.38172e-06, 
    8.712937e-06, 1.399208e-05, 1.782045e-05, 1.755467e-05, 1.84101e-05,
  1.822978e-05, 2.264945e-05, 2.129475e-05, 1.985566e-05, 1.768897e-05, 
    1.721233e-05, 1.107094e-05, 6.389252e-06, 3.081909e-06, 6.538218e-06, 
    1.14944e-05, 1.705006e-05, 2.02614e-05, 2.116157e-05, 2.271824e-05,
  2.294974e-05, 2.46819e-05, 2.725845e-05, 1.887197e-05, 1.20918e-05, 
    9.106185e-06, 1.134745e-05, 4.318433e-06, 6.244141e-06, 1.356244e-05, 
    1.789402e-05, 2.268352e-05, 2.618843e-05, 2.999685e-05, 3.510633e-05,
  2.196498e-05, 1.726756e-05, 1.396841e-05, 7.395427e-06, 4.798083e-06, 
    2.458852e-06, 3.300554e-06, 5.916845e-06, 1.26568e-05, 2.242422e-05, 
    3.157185e-05, 3.535731e-05, 4.14553e-05, 4.685473e-05, 5.04373e-05,
  2.712642e-06, 2.504274e-06, 3.579719e-06, 5.346666e-06, 7.105124e-06, 
    8.576723e-06, 8.134809e-06, 8.759289e-06, 1.116917e-05, 1.331619e-05, 
    1.28581e-05, 1.48405e-05, 1.191335e-05, 6.145695e-06, 4.09722e-06,
  1.492207e-06, 1.96541e-06, 3.018567e-06, 4.52094e-06, 7.032009e-06, 
    7.037098e-06, 1.237309e-05, 1.021539e-05, 8.271759e-06, 1.272623e-05, 
    1.48874e-05, 1.401423e-05, 1.093774e-05, 6.750673e-06, 5.97998e-06,
  5.817978e-06, 2.025145e-06, 2.900636e-06, 5.839815e-06, 8.246787e-06, 
    1.454343e-05, 1.49512e-05, 2.199853e-05, 1.220297e-05, 7.744551e-06, 
    9.60533e-06, 1.224461e-05, 1.200896e-05, 1.193108e-05, 1.145783e-05,
  5.971286e-06, 1.261621e-05, 1.086802e-05, 9.126166e-06, 1.523385e-05, 
    1.552657e-05, 1.631287e-05, 1.512292e-05, 1.309674e-05, 1.283317e-05, 
    9.393785e-06, 8.222629e-06, 8.918064e-06, 7.838382e-06, 9.697856e-06,
  6.168431e-06, 8.68995e-06, 9.329316e-06, 1.034836e-05, 1.799174e-05, 
    2.010018e-05, 1.93857e-05, 1.924238e-05, 1.004189e-05, 1.829017e-05, 
    1.397069e-05, 6.604368e-06, 5.757168e-06, 4.191476e-06, 5.749197e-06,
  6.25074e-06, 8.111992e-06, 9.470894e-06, 1.213045e-05, 1.734173e-05, 
    1.87572e-05, 2.022345e-05, 1.423963e-05, 7.259486e-06, 9.900919e-06, 
    9.718047e-06, 5.925979e-06, 3.757532e-06, 2.640196e-06, 2.827012e-06,
  1.29298e-05, 1.490355e-05, 1.151165e-05, 1.249911e-05, 1.317221e-05, 
    1.148895e-05, 1.472467e-05, 1.32134e-05, 6.217043e-06, 5.747735e-06, 
    5.408411e-06, 5.409712e-06, 4.030728e-06, 2.490973e-06, 2.341857e-06,
  2.241913e-05, 1.951883e-05, 8.094334e-06, 6.377691e-06, 6.39e-06, 
    1.201066e-05, 1.038766e-05, 9.352418e-06, 4.328457e-06, 6.020576e-06, 
    4.823441e-06, 3.70417e-06, 3.371722e-06, 2.537541e-06, 2.280394e-06,
  2.711447e-05, 1.679235e-05, 1.417654e-05, 4.194528e-06, 5.175074e-06, 
    7.478294e-06, 9.207594e-06, 7.309583e-06, 5.207409e-06, 4.179194e-06, 
    4.411095e-06, 4.102176e-06, 3.678515e-06, 3.171141e-06, 3.401224e-06,
  1.077321e-05, 9.221157e-06, 6.229514e-06, 4.773986e-06, 2.208194e-06, 
    6.647461e-06, 6.14332e-06, 6.804597e-06, 5.360828e-06, 4.266468e-06, 
    8.117017e-06, 8.572208e-06, 8.42255e-06, 7.386209e-06, 5.828303e-06,
  3.840651e-07, 1.765217e-07, 5.016885e-07, 2.158577e-07, 2.755755e-07, 
    2.731399e-06, 5.635671e-06, 4.660318e-06, 4.853614e-06, 5.691588e-06, 
    6.83401e-06, 8.844111e-06, 1.266345e-05, 1.273384e-05, 1.350209e-05,
  2.686668e-07, 1.592988e-07, 4.955518e-07, 6.663742e-07, 7.976369e-07, 
    2.060684e-06, 3.31113e-06, 3.602022e-06, 3.698011e-06, 3.418512e-06, 
    4.942668e-06, 8.145415e-06, 8.706125e-06, 9.244292e-06, 1.189582e-05,
  2.894509e-07, 2.935364e-07, 1.895864e-06, 7.498243e-07, 1.865556e-06, 
    2.549988e-05, 3.410013e-06, 3.109001e-06, 3.578021e-06, 4.211789e-06, 
    3.23098e-06, 5.502576e-06, 7.715413e-06, 1.091668e-05, 1.323828e-05,
  3.591529e-07, 5.297837e-07, 1.743816e-06, 1.097864e-06, 4.781115e-06, 
    1.220283e-05, 3.6594e-05, 3.434049e-06, 2.397522e-06, 3.987534e-06, 
    3.476195e-06, 3.424311e-06, 7.758799e-06, 1.123136e-05, 1.59747e-05,
  3.451283e-08, 3.15816e-07, 1.8288e-06, 3.400241e-06, 8.33154e-06, 
    9.546772e-06, 1.442898e-05, 4.223632e-05, 2.302089e-05, 4.758042e-06, 
    5.617811e-06, 4.937669e-06, 7.627167e-06, 1.040086e-05, 1.329435e-05,
  8.107126e-08, 2.467277e-07, 1.548116e-06, 3.943253e-06, 5.827784e-06, 
    5.83744e-06, 6.236033e-06, 9.81627e-06, 1.037317e-05, 9.782036e-06, 
    9.607021e-06, 6.763169e-06, 8.364426e-06, 1.064783e-05, 1.130418e-05,
  6.320101e-07, 2.675765e-07, 7.242904e-07, 3.348845e-06, 3.138067e-06, 
    4.063263e-06, 7.781719e-06, 1.029891e-05, 1.007911e-05, 1.129834e-05, 
    1.150554e-05, 1.097657e-05, 1.138877e-05, 1.542771e-05, 1.1721e-05,
  6.514675e-07, 1.624939e-06, 1.407355e-06, 1.92435e-06, 2.69985e-06, 
    5.080071e-06, 3.771346e-06, 8.133315e-06, 9.333871e-06, 1.402643e-05, 
    1.742339e-05, 1.710889e-05, 1.516334e-05, 1.157016e-05, 1.104205e-05,
  1.984006e-07, 6.799395e-07, 1.425269e-06, 1.877181e-06, 2.202686e-06, 
    3.050543e-06, 2.840426e-06, 6.70761e-06, 1.315804e-05, 2.090417e-05, 
    2.523594e-05, 2.295158e-05, 1.413607e-05, 1.06767e-05, 1.146895e-05,
  2.967785e-07, 1.349351e-06, 2.500939e-06, 2.536453e-06, 3.580121e-06, 
    5.506372e-06, 6.415374e-06, 1.230625e-05, 2.327991e-05, 3.264334e-05, 
    3.476553e-05, 2.560448e-05, 1.3006e-05, 1.097292e-05, 9.279913e-06,
  5.022125e-07, 4.876343e-07, 1.062837e-06, 4.850242e-07, 3.267139e-07, 
    6.219394e-07, 1.885552e-06, 2.705644e-06, 3.019082e-06, 4.849731e-06, 
    2.75113e-06, 3.043571e-06, 6.725968e-06, 1.435761e-05, 2.517514e-05,
  4.016132e-07, 3.772312e-07, 4.621212e-07, 2.815753e-07, 9.123709e-07, 
    1.148074e-06, 6.598507e-07, 1.378646e-06, 1.961181e-06, 2.452124e-06, 
    2.492878e-06, 4.277445e-06, 1.051829e-05, 2.622551e-05, 4.020839e-05,
  2.264533e-07, 3.874864e-07, 1.598073e-06, 2.23153e-06, 3.297949e-06, 
    9.837577e-06, 1.008509e-06, 6.928692e-07, 1.18603e-06, 3.096911e-06, 
    4.164699e-06, 6.841676e-06, 1.56947e-05, 2.970239e-05, 4.861616e-05,
  1.843367e-07, 4.927851e-07, 2.524438e-07, 2.123757e-07, 1.392009e-06, 
    5.207421e-06, 1.648233e-05, 2.023581e-06, 5.036795e-07, 1.569087e-06, 
    4.786316e-06, 7.453794e-06, 1.568088e-05, 3.30658e-05, 4.551437e-05,
  1.573882e-07, 3.051139e-07, 2.451435e-07, 5.112502e-07, 2.106649e-06, 
    5.548179e-06, 1.140413e-05, 3.838804e-05, 1.852233e-05, 2.186193e-06, 
    5.655804e-06, 1.033994e-05, 2.016591e-05, 3.591408e-05, 3.777352e-05,
  6.613329e-07, 5.819042e-07, 1.482848e-06, 2.337759e-06, 3.771004e-06, 
    5.430515e-06, 1.017163e-05, 1.028141e-05, 7.66242e-06, 8.093003e-06, 
    1.347548e-05, 1.802318e-05, 3.031482e-05, 3.590551e-05, 3.865415e-05,
  2.487742e-06, 3.956594e-06, 6.075561e-06, 3.650489e-06, 4.406945e-06, 
    5.727687e-06, 7.746574e-06, 9.19652e-06, 8.902977e-06, 9.618183e-06, 
    1.315907e-05, 1.992603e-05, 3.243521e-05, 3.91902e-05, 4.234448e-05,
  6.481514e-06, 9.834132e-06, 4.447188e-06, 2.8288e-06, 3.838249e-06, 
    5.740615e-06, 6.856819e-06, 7.655614e-06, 7.824059e-06, 7.942662e-06, 
    1.030448e-05, 2.000276e-05, 3.929298e-05, 4.290049e-05, 3.689745e-05,
  8.48614e-06, 4.971517e-06, 5.817016e-06, 4.623883e-06, 3.728993e-06, 
    4.990351e-06, 6.634426e-06, 7.468645e-06, 9.18925e-06, 8.314199e-06, 
    1.070243e-05, 2.366803e-05, 4.164073e-05, 3.686777e-05, 2.134641e-05,
  2.574814e-06, 5.173451e-06, 5.039382e-06, 5.391473e-06, 4.323024e-06, 
    3.787897e-06, 4.361867e-06, 5.852812e-06, 8.783e-06, 1.084559e-05, 
    1.60847e-05, 3.2495e-05, 3.777056e-05, 2.067564e-05, 7.316914e-06,
  2.21388e-07, 2.541748e-07, 2.37368e-07, 2.059799e-07, 2.62354e-07, 
    4.811828e-07, 8.85836e-07, 2.31068e-06, 4.563209e-06, 7.720011e-06, 
    9.047901e-06, 8.855822e-06, 1.345618e-05, 1.299247e-05, 1.213876e-05,
  3.60802e-07, 3.790773e-07, 2.690031e-07, 2.421861e-07, 1.457086e-06, 
    3.034585e-06, 1.66721e-06, 3.539144e-06, 4.926539e-06, 5.479312e-06, 
    6.67131e-06, 6.41728e-06, 8.483119e-06, 1.988072e-05, 1.771877e-05,
  5.496339e-07, 9.799041e-07, 8.564597e-07, 2.066082e-06, 3.765361e-06, 
    1.065513e-05, 2.8121e-06, 2.829704e-06, 5.110999e-06, 5.725082e-06, 
    3.513081e-06, 2.257312e-06, 5.048377e-06, 1.319488e-05, 2.323947e-05,
  4.370918e-06, 5.893289e-06, 8.869832e-06, 9.257677e-06, 3.220494e-06, 
    3.778436e-06, 1.67778e-05, 4.611047e-06, 1.68679e-06, 1.959426e-06, 
    3.156106e-06, 3.547464e-06, 8.928056e-06, 1.465905e-05, 2.542795e-05,
  6.804135e-06, 1.052275e-05, 1.111852e-05, 1.327433e-05, 1.725229e-05, 
    1.280708e-05, 7.161326e-06, 3.596271e-05, 2.190336e-05, 3.14309e-06, 
    6.999227e-06, 9.306063e-06, 1.170886e-05, 1.513894e-05, 2.207549e-05,
  5.50231e-06, 1.045981e-05, 1.357653e-05, 1.495061e-05, 1.89088e-05, 
    1.605894e-05, 1.515364e-05, 9.228651e-06, 9.438689e-06, 1.184062e-05, 
    1.510001e-05, 1.238953e-05, 1.382647e-05, 1.658368e-05, 2.261197e-05,
  9.769252e-06, 1.51503e-05, 1.540138e-05, 1.187947e-05, 1.372791e-05, 
    1.190106e-05, 1.361532e-05, 1.216061e-05, 1.057867e-05, 1.051357e-05, 
    1.16565e-05, 1.21783e-05, 1.328576e-05, 1.71514e-05, 2.228936e-05,
  1.329461e-05, 1.516577e-05, 1.263922e-05, 6.788394e-06, 5.2654e-06, 
    8.044203e-06, 1.032769e-05, 9.858147e-06, 9.342401e-06, 1.164043e-05, 
    1.339007e-05, 1.193345e-05, 1.360508e-05, 2.016733e-05, 2.529125e-05,
  2.075547e-05, 1.368477e-05, 1.300195e-05, 8.597317e-06, 9.277812e-06, 
    1.029244e-05, 1.234626e-05, 1.277916e-05, 1.318694e-05, 1.43206e-05, 
    1.144037e-05, 1.204444e-05, 1.608627e-05, 2.284793e-05, 3.579233e-05,
  2.858484e-05, 2.508447e-05, 2.388624e-05, 1.989809e-05, 1.565431e-05, 
    1.30195e-05, 1.151986e-05, 1.083856e-05, 1.07139e-05, 9.165125e-06, 
    9.106899e-06, 9.815093e-06, 1.638264e-05, 3.135344e-05, 4.371831e-05,
  3.99376e-08, 6.108696e-08, 1.24767e-07, 1.756948e-07, 2.116063e-07, 
    2.778291e-07, 4.132345e-07, 7.247399e-07, 1.661385e-06, 3.685432e-06, 
    5.111272e-06, 5.59421e-06, 9.200289e-06, 1.142072e-05, 1.081102e-05,
  5.389086e-07, 7.139918e-07, 9.445865e-07, 1.105934e-06, 1.213961e-06, 
    1.33079e-06, 1.52204e-06, 1.964904e-06, 2.68348e-06, 4.100815e-06, 
    5.658878e-06, 8.469759e-06, 1.074279e-05, 1.724444e-05, 1.239649e-05,
  1.680995e-06, 1.786492e-06, 1.766143e-06, 1.922582e-06, 2.346866e-06, 
    4.482462e-06, 1.97239e-06, 2.518579e-06, 4.530018e-06, 4.662596e-06, 
    4.070663e-06, 4.585329e-06, 7.493186e-06, 9.390167e-06, 1.254977e-05,
  6.112529e-06, 3.962197e-06, 2.725314e-06, 2.928829e-06, 4.418564e-06, 
    5.742394e-06, 9.227163e-06, 3.337674e-06, 1.993071e-06, 5.089389e-06, 
    6.707646e-06, 4.41081e-06, 5.776598e-06, 8.42971e-06, 1.275858e-05,
  2.145859e-05, 1.987347e-05, 2.134094e-05, 2.621114e-05, 3.762413e-05, 
    2.840435e-05, 2.03073e-05, 2.183995e-05, 1.891009e-05, 8.452536e-06, 
    1.544321e-05, 6.134293e-06, 4.858897e-06, 7.783591e-06, 1.359895e-05,
  2.964655e-05, 3.541809e-05, 3.598825e-05, 3.848875e-05, 3.669945e-05, 
    2.969666e-05, 2.967243e-05, 1.557203e-05, 3.756122e-06, 8.021007e-06, 
    1.506153e-05, 9.244418e-06, 7.643915e-06, 8.359727e-06, 1.132218e-05,
  3.552568e-05, 3.247815e-05, 2.854158e-05, 2.766014e-05, 2.317514e-05, 
    1.736047e-05, 2.048677e-05, 2.125581e-05, 8.941094e-06, 7.351142e-06, 
    8.729132e-06, 1.060648e-05, 1.117123e-05, 9.978974e-06, 9.468687e-06,
  3.28032e-05, 2.763646e-05, 2.791094e-05, 1.973728e-05, 1.681809e-05, 
    1.697302e-05, 8.756057e-06, 6.221011e-06, 2.567554e-06, 3.755209e-06, 
    7.790414e-06, 9.515114e-06, 9.072823e-06, 9.437438e-06, 9.732744e-06,
  4.737316e-05, 4.430607e-05, 4.050917e-05, 3.308164e-05, 2.907871e-05, 
    2.438668e-05, 2.047354e-05, 1.573738e-05, 1.176487e-05, 8.524093e-06, 
    5.665393e-06, 6.783766e-06, 1.040341e-05, 1.264823e-05, 1.457223e-05,
  4.288847e-05, 4.057396e-05, 3.738966e-05, 3.376731e-05, 3.523496e-05, 
    3.98864e-05, 4.364654e-05, 4.364772e-05, 3.561191e-05, 2.446151e-05, 
    1.421363e-05, 1.345277e-05, 1.821972e-05, 1.938287e-05, 1.807407e-05,
  3.076706e-07, 2.613732e-06, 3.738907e-07, 5.518625e-07, 8.919779e-07, 
    8.532185e-07, 6.771242e-07, 3.589223e-07, 2.635633e-07, 3.283233e-07, 
    1.415088e-07, 1.625562e-07, 2.872985e-07, 4.43296e-07, 7.537236e-07,
  5.843681e-06, 2.202196e-06, 1.539816e-07, 4.317191e-07, 1.138872e-06, 
    7.595706e-07, 1.325699e-06, 4.447053e-07, 4.587274e-07, 3.14851e-07, 
    2.657289e-07, 2.095146e-07, 3.802615e-07, 1.012443e-06, 1.183865e-06,
  1.700381e-05, 7.431627e-06, 4.641727e-06, 1.699834e-06, 2.24362e-06, 
    1.292367e-06, 1.735072e-07, 2.752202e-07, 5.795746e-07, 3.394312e-07, 
    2.268833e-07, 2.750318e-07, 6.152689e-07, 1.916537e-06, 4.580392e-06,
  4.135493e-05, 2.763361e-05, 1.908494e-05, 1.50719e-05, 5.833544e-06, 
    4.843499e-06, 3.582637e-06, 7.285391e-07, 4.169605e-07, 2.424181e-07, 
    1.505892e-06, 2.143077e-06, 2.58146e-06, 5.447389e-06, 1.021302e-05,
  4.162294e-05, 4.122565e-05, 4.720215e-05, 5.318121e-05, 4.943652e-05, 
    2.736783e-05, 1.761099e-05, 1.661221e-05, 5.350209e-06, 1.069006e-06, 
    6.249666e-06, 3.207416e-06, 1.788335e-06, 4.528611e-06, 8.724636e-06,
  2.069525e-05, 2.141578e-05, 2.519459e-05, 2.918135e-05, 3.827305e-05, 
    4.901372e-05, 5.302395e-05, 3.04258e-05, 8.193886e-06, 1.175344e-05, 
    9.240052e-06, 4.096635e-06, 3.586321e-06, 6.115865e-06, 8.081334e-06,
  1.982664e-05, 1.484911e-05, 9.78657e-06, 7.012738e-06, 9.27594e-06, 
    1.122249e-05, 1.988496e-05, 2.365506e-05, 1.40003e-05, 4.531436e-06, 
    4.425793e-06, 5.581861e-06, 7.691438e-06, 1.002105e-05, 1.138633e-05,
  3.459427e-05, 2.651498e-05, 1.938177e-05, 1.472673e-05, 1.335445e-05, 
    1.638307e-05, 1.359567e-05, 8.856251e-06, 9.369944e-06, 2.293032e-06, 
    5.623784e-06, 6.515153e-06, 6.556168e-06, 8.134001e-06, 1.013577e-05,
  3.163177e-05, 3.230822e-05, 3.087076e-05, 2.633795e-05, 2.158091e-05, 
    1.886013e-05, 1.456324e-05, 9.130246e-06, 9.81886e-06, 7.003363e-06, 
    7.687046e-06, 6.725973e-06, 9.728024e-06, 1.139985e-05, 1.247789e-05,
  3.136e-05, 2.937903e-05, 3.246044e-05, 2.763657e-05, 1.926949e-05, 
    1.239243e-05, 6.120215e-06, 4.077523e-06, 1.190619e-05, 1.82357e-05, 
    2.476963e-05, 2.462787e-05, 2.735809e-05, 2.853524e-05, 3.22389e-05,
  5.580314e-06, 1.018319e-05, 7.312902e-06, 9.036933e-06, 4.877723e-06, 
    4.928887e-06, 4.444114e-06, 1.85424e-06, 2.919305e-06, 3.636683e-06, 
    2.567854e-06, 2.709181e-06, 4.30108e-06, 3.729281e-06, 3.125452e-06,
  1.172744e-05, 6.493171e-06, 1.845406e-06, 3.349855e-06, 5.955961e-06, 
    3.238957e-06, 1.359465e-05, 1.422912e-06, 2.194432e-06, 2.783975e-06, 
    2.589696e-06, 3.49795e-06, 5.111611e-06, 4.558991e-06, 2.089199e-06,
  1.337203e-05, 1.366415e-05, 2.262834e-05, 2.13572e-05, 1.852256e-05, 
    9.036547e-06, 4.951658e-06, 6.633722e-06, 4.057227e-06, 2.982903e-06, 
    2.450635e-06, 2.583969e-06, 3.818737e-06, 3.074518e-06, 3.332567e-06,
  2.837044e-05, 3.190703e-05, 2.907468e-05, 2.300585e-05, 2.262209e-05, 
    1.923715e-05, 1.467136e-05, 7.423662e-06, 6.4601e-06, 8.900789e-07, 
    2.895024e-06, 3.399142e-06, 4.14448e-06, 5.248791e-06, 7.409958e-06,
  1.634134e-05, 1.31304e-05, 1.716735e-05, 2.549909e-05, 3.586694e-05, 
    2.118099e-05, 3.100502e-05, 2.290093e-05, 4.95527e-06, 2.844263e-06, 
    4.959097e-06, 3.541711e-06, 3.290022e-06, 3.790158e-06, 4.477632e-06,
  2.036548e-05, 1.276506e-05, 1.223558e-05, 1.975603e-05, 2.012873e-05, 
    2.508864e-05, 4.426536e-05, 3.061244e-05, 1.559266e-05, 1.424377e-05, 
    6.149046e-06, 6.070788e-06, 1.021462e-05, 1.148559e-05, 1.497694e-05,
  2.495079e-05, 2.230756e-05, 1.560898e-05, 1.060681e-05, 9.505251e-06, 
    1.2751e-05, 1.806529e-05, 2.104975e-05, 1.848365e-05, 4.46252e-06, 
    1.972397e-06, 4.495121e-06, 4.959329e-06, 5.418674e-06, 7.151718e-06,
  2.329841e-05, 2.342032e-05, 1.956859e-05, 1.781234e-05, 1.406216e-05, 
    1.391065e-05, 1.1883e-05, 1.086926e-05, 6.435097e-06, 9.800109e-07, 
    8.820581e-07, 1.035522e-06, 4.378936e-07, 7.435826e-07, 8.217403e-07,
  2.186119e-05, 2.118791e-05, 2.111896e-05, 1.958266e-05, 1.90615e-05, 
    1.580654e-05, 1.096367e-05, 1.050553e-05, 8.701548e-06, 6.781045e-06, 
    1.143064e-05, 1.056245e-06, 5.512788e-07, 5.998613e-07, 1.311605e-06,
  1.676279e-05, 1.624359e-05, 1.581949e-05, 1.39396e-05, 1.46959e-05, 
    1.052609e-05, 5.941972e-06, 4.162531e-06, 3.865061e-06, 4.216454e-06, 
    8.568078e-06, 5.004872e-06, 3.07095e-06, 3.183286e-06, 6.583835e-06,
  3.568265e-06, 6.630577e-06, 6.300366e-06, 1.046613e-05, 5.064956e-06, 
    5.595305e-06, 8.997989e-06, 3.458402e-06, 7.031003e-06, 7.212685e-06, 
    4.814411e-06, 7.363697e-06, 1.17497e-05, 1.152628e-05, 6.951102e-06,
  7.751715e-06, 7.542379e-06, 4.008501e-06, 2.975512e-06, 4.202318e-06, 
    6.782427e-06, 1.334895e-05, 2.972282e-06, 4.543936e-06, 6.3944e-06, 
    7.244479e-06, 1.252587e-05, 1.421664e-05, 9.533675e-06, 5.433914e-06,
  2.802572e-05, 9.888328e-06, 1.273364e-05, 1.575854e-05, 1.793148e-05, 
    9.606872e-06, 7.524045e-06, 1.941877e-05, 1.104683e-05, 7.010698e-06, 
    5.704051e-06, 8.957979e-06, 1.244694e-05, 1.137125e-05, 1.367022e-05,
  4.383597e-05, 4.56715e-05, 3.561965e-05, 3.536737e-05, 1.39903e-05, 
    1.939846e-05, 1.141623e-05, 1.128625e-05, 9.847271e-06, 2.256627e-06, 
    7.15223e-06, 9.838568e-06, 1.198142e-05, 1.967145e-05, 2.462064e-05,
  3.260334e-05, 2.238513e-05, 2.429815e-05, 2.529522e-05, 3.270152e-05, 
    1.06272e-05, 2.862905e-05, 3.18705e-05, 1.157491e-05, 1.30079e-06, 
    5.283827e-06, 6.42504e-06, 9.594321e-06, 1.591751e-05, 2.066633e-05,
  3.043081e-05, 2.689e-05, 2.722449e-05, 2.167959e-05, 1.827173e-05, 
    2.559198e-05, 3.230468e-05, 1.313118e-05, 8.478103e-06, 8.221421e-06, 
    7.055124e-06, 5.727885e-06, 9.762592e-06, 1.2987e-05, 1.499764e-05,
  3.061816e-05, 3.234331e-05, 3.05859e-05, 2.230706e-05, 1.864404e-05, 
    1.771286e-05, 1.97111e-05, 2.270607e-05, 1.340603e-05, 3.839635e-06, 
    2.938917e-06, 6.152762e-06, 1.064091e-05, 1.00263e-05, 9.926863e-06,
  3.332934e-05, 3.403701e-05, 3.407001e-05, 2.516096e-05, 2.441115e-05, 
    2.238048e-05, 1.873613e-05, 1.417917e-05, 6.550285e-06, 1.649805e-06, 
    1.736823e-06, 3.536629e-06, 4.251148e-06, 5.783532e-06, 6.249614e-06,
  3.227837e-05, 3.725358e-05, 3.869264e-05, 2.79078e-05, 2.241462e-05, 
    1.829851e-05, 1.662803e-05, 1.204544e-05, 6.14469e-06, 4.231255e-06, 
    6.094985e-06, 8.955165e-07, 1.5159e-06, 2.833894e-06, 3.271397e-06,
  2.112007e-05, 2.359346e-05, 2.909814e-05, 2.067833e-05, 1.456658e-05, 
    1.105219e-05, 7.087957e-06, 6.149265e-06, 5.882649e-06, 2.731406e-06, 
    6.061031e-06, 1.459681e-06, 1.338535e-06, 1.762714e-06, 2.083945e-06,
  1.21951e-05, 9.970094e-06, 1.125878e-05, 1.184364e-05, 4.685462e-06, 
    3.788193e-06, 8.37284e-06, 4.16701e-06, 4.617024e-06, 4.84069e-06, 
    3.826625e-06, 4.614615e-06, 5.763905e-06, 5.605177e-06, 4.565331e-06,
  9.652812e-06, 8.546115e-06, 8.810194e-06, 5.950043e-06, 4.717644e-06, 
    1.251134e-05, 1.323813e-05, 4.309903e-06, 2.892195e-06, 4.270714e-06, 
    4.889191e-06, 7.435454e-06, 7.027097e-06, 4.727892e-06, 4.007893e-06,
  2.526126e-05, 1.585629e-05, 1.771357e-05, 1.827459e-05, 1.610512e-05, 
    1.187675e-05, 4.743673e-06, 4.355838e-06, 2.261469e-06, 1.921934e-06, 
    3.270646e-06, 4.148853e-06, 5.121152e-06, 5.260849e-06, 8.515711e-06,
  2.406459e-05, 2.65559e-05, 3.182537e-05, 3.792911e-05, 3.1349e-05, 
    2.333542e-05, 2.603485e-05, 1.314301e-05, 2.058494e-06, 1.123669e-06, 
    2.423764e-06, 2.962452e-06, 3.346505e-06, 7.968379e-06, 1.160736e-05,
  1.924642e-05, 1.70644e-05, 2.16656e-05, 2.835803e-05, 4.33171e-05, 
    4.941746e-05, 5.24043e-05, 3.963527e-05, 1.563851e-05, 1.239445e-06, 
    5.389544e-06, 6.048129e-06, 2.793023e-06, 6.203823e-06, 9.404684e-06,
  2.520214e-05, 2.006432e-05, 1.657294e-05, 1.860112e-05, 2.992947e-05, 
    4.383936e-05, 5.666413e-05, 3.670377e-05, 1.845244e-05, 1.767719e-05, 
    7.825043e-06, 1.83897e-06, 3.563865e-06, 6.652613e-06, 8.737001e-06,
  2.723043e-05, 2.222284e-05, 1.333214e-05, 1.654583e-05, 1.96775e-05, 
    2.516105e-05, 3.552268e-05, 3.812843e-05, 3.213017e-05, 2.3934e-05, 
    1.341293e-05, 7.783088e-06, 6.309546e-06, 6.573769e-06, 7.548867e-06,
  1.831582e-05, 1.740827e-05, 1.462403e-05, 1.749837e-05, 1.833015e-05, 
    2.109617e-05, 1.600808e-05, 1.264986e-05, 4.365928e-06, 6.331158e-06, 
    1.51338e-05, 1.996994e-05, 1.399775e-05, 9.099787e-06, 7.28193e-06,
  1.536406e-05, 1.52274e-05, 1.708686e-05, 1.760757e-05, 1.73991e-05, 
    1.565182e-05, 1.341209e-05, 9.53629e-06, 4.569225e-06, 5.008696e-06, 
    6.44103e-06, 1.069577e-05, 1.240378e-05, 1.080577e-05, 7.960326e-06,
  2.934844e-05, 1.214242e-05, 1.43362e-05, 1.38436e-05, 1.123007e-05, 
    7.831944e-06, 5.253338e-06, 4.262636e-06, 4.454429e-06, 2.51918e-06, 
    2.066276e-06, 2.05112e-06, 4.501399e-06, 4.78894e-06, 5.36687e-06,
  1.726794e-05, 1.361447e-05, 8.810215e-06, 1.044078e-05, 7.563349e-06, 
    7.10169e-06, 5.457326e-06, 1.890182e-06, 2.833369e-06, 3.794354e-06, 
    3.641313e-06, 4.715539e-06, 4.99275e-06, 3.987637e-06, 3.070571e-06,
  3.478982e-05, 2.470152e-05, 1.322908e-05, 1.389166e-05, 1.528264e-05, 
    1.173802e-05, 8.906609e-06, 2.960178e-06, 3.142663e-06, 2.926072e-06, 
    4.644201e-06, 8.433564e-06, 6.864108e-06, 4.554705e-06, 3.244765e-06,
  3.882687e-05, 4.185108e-05, 3.248525e-05, 1.947543e-05, 1.712518e-05, 
    1.559787e-05, 9.634991e-06, 1.044612e-05, 8.006269e-06, 4.555801e-06, 
    4.725719e-06, 7.906272e-06, 7.234786e-06, 6.985223e-06, 7.364358e-06,
  4.595118e-05, 3.361172e-05, 2.290675e-05, 1.436894e-05, 1.007407e-05, 
    1.014397e-05, 1.879811e-05, 1.985595e-05, 1.394851e-05, 6.580628e-06, 
    6.270385e-06, 5.936372e-06, 6.732026e-06, 9.949935e-06, 1.127233e-05,
  4.15718e-05, 2.311572e-05, 5.537352e-06, 9.5007e-06, 1.505661e-05, 
    1.82387e-05, 1.306498e-05, 2.096061e-05, 1.114009e-05, 1.202148e-05, 
    1.328105e-05, 6.163222e-06, 5.961147e-06, 8.617349e-06, 1.038881e-05,
  3.701841e-05, 1.1285e-05, 1.029344e-06, 4.521829e-06, 1.429976e-05, 
    2.738965e-05, 3.159625e-05, 8.215036e-06, 7.079916e-06, 1.019738e-05, 
    8.069128e-06, 6.814507e-06, 6.334636e-06, 6.777739e-06, 9.510956e-06,
  3.501832e-05, 1.387928e-05, 4.785323e-06, 5.265224e-06, 1.223272e-05, 
    2.206524e-05, 2.957881e-05, 1.999864e-05, 3.974304e-06, 2.425425e-06, 
    4.12338e-06, 7.019328e-06, 7.602669e-06, 5.751854e-06, 7.079163e-06,
  8.669456e-05, 4.286025e-05, 1.369377e-05, 1.771688e-05, 2.793329e-05, 
    3.184427e-05, 2.192597e-05, 1.022785e-05, 2.282846e-06, 8.393633e-07, 
    5.993393e-07, 5.779737e-06, 8.232157e-06, 7.628558e-06, 7.318808e-06,
  0.000113129, 4.351574e-05, 2.235454e-05, 2.63927e-05, 3.264225e-05, 
    3.303308e-05, 2.453807e-05, 1.307554e-05, 2.594948e-06, 3.948196e-06, 
    2.727197e-06, 3.420046e-06, 9.03857e-06, 1.035308e-05, 8.527365e-06,
  4.058194e-05, 2.552566e-05, 2.032095e-05, 1.891474e-05, 1.432643e-05, 
    7.280537e-06, 6.440712e-06, 3.937231e-06, 2.82073e-06, 1.370105e-06, 
    1.84626e-06, 1.998196e-06, 8.804999e-06, 1.473813e-05, 1.398986e-05,
  3.046773e-05, 2.912692e-05, 2.437296e-05, 1.756803e-05, 1.271595e-05, 
    8.504755e-06, 7.574607e-06, 2.325484e-06, 2.663611e-06, 4.124756e-06, 
    2.330102e-06, 1.876508e-06, 2.795973e-06, 3.623851e-06, 5.305765e-06,
  1.831821e-05, 2.629041e-05, 2.219061e-05, 1.92172e-05, 1.899452e-05, 
    1.667046e-05, 1.287764e-05, 4.232314e-06, 3.403675e-06, 4.141798e-06, 
    5.131345e-06, 5.53012e-06, 3.08906e-06, 2.642438e-06, 3.305082e-06,
  2.780463e-05, 2.895119e-05, 2.678732e-05, 1.521256e-05, 1.496814e-05, 
    1.177697e-05, 1.411966e-05, 1.511249e-05, 1.089622e-05, 5.540082e-06, 
    6.59057e-06, 5.936362e-06, 4.053482e-06, 2.197938e-06, 2.445336e-06,
  4.921764e-05, 4.463702e-05, 3.785638e-05, 2.750148e-05, 1.538866e-05, 
    8.75058e-06, 1.185755e-05, 1.656792e-05, 1.043704e-05, 7.144717e-06, 
    7.594652e-06, 5.704402e-06, 5.260397e-06, 4.420908e-06, 4.366958e-06,
  6.131966e-05, 4.369192e-05, 3.245121e-05, 3.229139e-05, 2.308422e-05, 
    2.09415e-05, 1.016442e-05, 1.212206e-05, 8.401584e-06, 3.101882e-06, 
    9.50899e-06, 7.485654e-06, 6.91255e-06, 5.277844e-06, 4.601406e-06,
  4.531816e-05, 2.441487e-05, 2.429748e-05, 2.103072e-05, 1.983637e-05, 
    1.738043e-05, 2.163481e-05, 6.235668e-06, 2.417768e-06, 5.346315e-06, 
    5.698912e-06, 6.134522e-06, 8.135667e-06, 7.142005e-06, 5.951656e-06,
  3.038153e-05, 2.341926e-05, 2.35487e-05, 2.248992e-05, 1.535363e-05, 
    1.313138e-05, 2.322866e-05, 1.965932e-05, 4.420694e-06, 3.128412e-06, 
    1.691039e-06, 2.61893e-06, 5.40754e-06, 6.747217e-06, 7.006117e-06,
  8.139233e-05, 5.205841e-05, 3.260065e-05, 2.100719e-05, 1.879807e-05, 
    1.970261e-05, 2.945697e-05, 2.606462e-05, 3.929483e-06, 2.485749e-06, 
    2.054518e-06, 2.024634e-06, 2.16405e-06, 2.200837e-06, 3.924537e-06,
  0.00011925, 6.398658e-05, 2.798241e-05, 1.287008e-05, 1.312123e-05, 
    1.170019e-05, 2.277989e-05, 4.029545e-05, 2.531429e-05, 1.124401e-05, 
    3.484107e-06, 1.340461e-06, 7.92075e-07, 6.104147e-07, 1.125018e-06,
  4.299207e-05, 2.44804e-05, 1.134082e-05, 1.055109e-05, 7.69019e-06, 
    6.664029e-06, 1.590584e-05, 3.742243e-05, 4.134321e-05, 3.078369e-05, 
    1.051989e-05, 1.872592e-06, 3.042517e-07, 1.550502e-07, 7.026804e-07,
  5.866977e-06, 1.277197e-05, 1.533523e-05, 2.13543e-05, 2.750404e-05, 
    2.723825e-05, 2.058691e-05, 9.562445e-06, 4.190881e-06, 3.258809e-06, 
    2.776021e-06, 2.167914e-06, 2.521228e-06, 3.483304e-06, 7.59003e-06,
  2.980862e-06, 8.574632e-06, 1.570768e-05, 2.011897e-05, 2.838331e-05, 
    2.641607e-05, 2.302622e-05, 1.752528e-05, 1.218343e-05, 7.843484e-06, 
    3.632969e-06, 3.0143e-06, 1.403333e-06, 1.969694e-06, 5.502703e-06,
  7.817965e-06, 1.622334e-05, 1.806938e-05, 1.8772e-05, 1.646416e-05, 
    2.174721e-05, 2.206231e-05, 2.685835e-05, 2.254885e-05, 1.492209e-05, 
    8.372655e-06, 4.984683e-06, 1.773048e-06, 1.241375e-06, 3.80689e-06,
  2.852659e-05, 4.591803e-05, 4.387434e-05, 3.106477e-05, 1.866039e-05, 
    1.072678e-05, 2.214375e-05, 2.619059e-05, 2.243646e-05, 1.561975e-05, 
    9.43168e-06, 4.469458e-06, 1.822034e-06, 1.971888e-06, 2.293457e-06,
  5.841381e-05, 5.591639e-05, 4.575165e-05, 4.012682e-05, 3.701903e-05, 
    2.429189e-05, 1.261101e-05, 1.218129e-05, 1.096423e-05, 5.699339e-06, 
    5.203757e-06, 2.036133e-06, 2.457349e-06, 2.480267e-06, 1.726099e-06,
  5.420929e-05, 3.486199e-05, 3.504971e-05, 3.706834e-05, 3.890053e-05, 
    4.002617e-05, 2.595053e-05, 1.308529e-05, 6.449236e-06, 6.458316e-06, 
    2.176598e-06, 6.405665e-07, 2.163675e-06, 2.712383e-06, 1.659625e-06,
  5.301091e-05, 4.639283e-05, 4.101628e-05, 3.592556e-05, 3.315708e-05, 
    3.041739e-05, 2.606589e-05, 2.501202e-05, 1.286612e-05, 6.751879e-06, 
    1.16366e-06, 1.825293e-06, 2.80293e-06, 2.301924e-06, 2.141325e-06,
  5.66676e-05, 5.240634e-05, 3.862749e-05, 3.077725e-05, 2.431395e-05, 
    2.113943e-05, 1.454954e-05, 1.161517e-05, 4.043912e-06, 5.459186e-06, 
    6.508935e-06, 5.612314e-06, 4.141719e-06, 2.646005e-06, 2.889871e-06,
  4.524839e-05, 4.334838e-05, 4.029241e-05, 2.503583e-05, 1.319617e-05, 
    9.985339e-06, 8.282725e-06, 6.596882e-06, 2.203941e-06, 1.461652e-06, 
    6.132853e-06, 6.399839e-06, 4.91572e-06, 3.161143e-06, 3.102548e-06,
  2.784846e-05, 3.037666e-05, 2.264767e-05, 9.578094e-06, 5.639591e-06, 
    5.065674e-06, 5.116042e-06, 5.307032e-06, 3.96382e-06, 1.708347e-06, 
    3.605384e-06, 5.667682e-06, 5.832377e-06, 4.63118e-06, 3.296218e-06,
  2.230954e-06, 1.983851e-06, 1.596967e-06, 2.740012e-06, 2.219149e-06, 
    3.148536e-06, 2.838648e-06, 1.95312e-06, 9.155815e-07, 1.142656e-06, 
    1.505601e-06, 2.254616e-06, 3.159747e-06, 3.933077e-06, 4.392729e-06,
  6.21698e-06, 4.596799e-06, 4.306203e-06, 5.32448e-06, 7.893709e-06, 
    9.228653e-06, 5.412831e-06, 3.363365e-06, 2.312606e-06, 2.565033e-06, 
    2.650913e-06, 4.188122e-06, 5.367323e-06, 3.009484e-06, 3.385014e-06,
  9.013596e-06, 1.101226e-05, 9.725253e-06, 5.79372e-06, 8.494966e-06, 
    8.905677e-06, 9.340602e-06, 1.333732e-05, 1.132949e-05, 7.664496e-06, 
    4.941177e-06, 3.800862e-06, 3.178838e-06, 3.380311e-06, 5.173967e-06,
  4.462645e-05, 3.132409e-05, 3.628789e-05, 1.916722e-05, 8.976848e-06, 
    7.819944e-06, 1.29105e-05, 1.654806e-05, 1.476682e-05, 1.065049e-05, 
    7.750008e-06, 5.698814e-06, 6.29551e-06, 6.359821e-06, 6.33533e-06,
  5.111007e-05, 4.415593e-05, 5.169122e-05, 3.965834e-05, 3.188848e-05, 
    2.62369e-05, 1.535698e-05, 1.957085e-05, 1.65549e-05, 5.247752e-06, 
    1.026705e-05, 6.570717e-06, 7.496072e-06, 5.937809e-06, 4.126695e-06,
  4.875611e-05, 4.45322e-05, 5.613244e-05, 5.976858e-05, 6.805267e-05, 
    5.648512e-05, 3.931066e-05, 1.485137e-05, 8.362393e-06, 1.198181e-05, 
    1.086596e-05, 7.009657e-06, 8.645434e-06, 6.092421e-06, 5.29909e-06,
  4.274205e-05, 4.292443e-05, 3.763827e-05, 4.30545e-05, 4.677424e-05, 
    4.495781e-05, 3.937364e-05, 3.565418e-05, 2.325311e-05, 1.891167e-05, 
    1.293882e-05, 1.099899e-05, 9.318615e-06, 6.023538e-06, 4.75241e-06,
  2.807795e-05, 4.152516e-05, 4.00004e-05, 2.845212e-05, 2.524388e-05, 
    2.270116e-05, 1.87504e-05, 2.018739e-05, 1.757079e-05, 1.553735e-05, 
    1.78159e-05, 1.699364e-05, 1.229666e-05, 7.573897e-06, 4.579656e-06,
  2.075901e-05, 3.869065e-05, 4.221686e-05, 3.098447e-05, 1.320565e-05, 
    8.497696e-06, 8.051783e-06, 1.197878e-05, 1.755895e-05, 2.044306e-05, 
    2.322222e-05, 2.033427e-05, 1.537949e-05, 9.877311e-06, 4.338161e-06,
  1.249722e-05, 2.019136e-05, 2.442008e-05, 1.107827e-05, 4.771007e-06, 
    4.632812e-06, 4.529563e-06, 5.523545e-06, 1.271892e-05, 1.610969e-05, 
    2.175384e-05, 2.222773e-05, 1.639341e-05, 9.063961e-06, 3.498764e-06,
  3.668737e-06, 2.530715e-06, 2.364348e-06, 2.329917e-06, 1.041667e-05, 
    1.315888e-05, 1.78967e-05, 1.757368e-05, 1.687441e-05, 1.429895e-05, 
    1.52618e-05, 1.815478e-05, 1.645375e-05, 1.223125e-05, 1.15655e-05,
  7.097921e-06, 1.248767e-06, 2.462885e-06, 1.234573e-06, 8.119626e-06, 
    1.181808e-05, 2.053951e-05, 1.677395e-05, 1.425449e-05, 1.849218e-05, 
    1.340823e-05, 1.650496e-05, 1.333907e-05, 7.825968e-06, 3.329933e-06,
  4.211209e-05, 1.257918e-05, 1.83991e-06, 5.708673e-07, 3.942881e-06, 
    5.273338e-06, 1.503314e-05, 2.293698e-05, 2.229204e-05, 2.116296e-05, 
    2.237862e-05, 1.804723e-05, 1.925104e-05, 1.092496e-05, 3.364416e-06,
  4.100969e-05, 6.011146e-05, 2.503239e-05, 1.154352e-05, 2.313172e-06, 
    5.562143e-06, 7.450498e-06, 1.475149e-05, 2.280428e-05, 2.724973e-05, 
    2.067518e-05, 1.768206e-05, 2.045225e-05, 1.449821e-05, 5.485299e-06,
  2.717459e-05, 5.165634e-05, 6.136546e-05, 2.732684e-05, 1.638057e-05, 
    9.1419e-06, 6.817955e-06, 1.794765e-06, 8.551877e-06, 1.901353e-05, 
    1.925894e-05, 1.441428e-05, 1.280955e-05, 8.750286e-06, 3.97168e-06,
  1.645563e-05, 4.377124e-05, 6.541172e-05, 4.869594e-05, 3.458444e-05, 
    2.518062e-05, 2.164878e-05, 9.649612e-06, 6.589878e-06, 1.350003e-05, 
    1.40746e-05, 1.319749e-05, 8.036625e-06, 3.357041e-06, 2.242428e-06,
  2.700808e-05, 3.65748e-05, 4.703565e-05, 5.303884e-05, 4.924081e-05, 
    3.712191e-05, 2.267826e-05, 2.029523e-05, 1.442872e-05, 1.339805e-05, 
    1.362252e-05, 1.105495e-05, 5.712034e-06, 2.791634e-06, 2.48068e-06,
  4.250103e-05, 4.41885e-05, 3.808317e-05, 3.98594e-05, 3.44157e-05, 
    3.407906e-05, 2.079693e-05, 1.242265e-05, 8.726824e-06, 9.749434e-06, 
    1.052638e-05, 1.024219e-05, 4.813386e-06, 3.45351e-06, 4.175528e-06,
  4.897351e-05, 4.943293e-05, 4.238148e-05, 2.255443e-05, 1.383106e-05, 
    1.257154e-05, 1.090441e-05, 7.778933e-06, 6.981464e-06, 8.010765e-06, 
    7.877193e-06, 6.886567e-06, 4.953535e-06, 6.03862e-06, 6.966564e-06,
  3.274261e-05, 3.534878e-05, 2.382463e-05, 8.920401e-06, 3.870369e-06, 
    3.469729e-06, 4.418179e-06, 6.301088e-06, 6.843102e-06, 6.618459e-06, 
    6.614979e-06, 5.976761e-06, 6.766949e-06, 9.750543e-06, 1.015241e-05,
  2.838422e-07, 2.339664e-06, 3.770786e-06, 1.211539e-05, 2.664841e-05, 
    3.936296e-05, 3.492589e-05, 2.132201e-05, 1.767775e-05, 1.040291e-05, 
    5.103002e-06, 3.3895e-06, 4.373248e-06, 4.592567e-06, 4.33749e-06,
  3.630637e-06, 1.099585e-06, 5.037138e-06, 1.363636e-05, 2.794571e-05, 
    3.492305e-05, 2.679159e-05, 1.664249e-05, 1.208505e-05, 9.479327e-06, 
    3.634144e-06, 5.759815e-06, 3.630088e-06, 2.71721e-06, 3.590481e-06,
  3.819317e-05, 1.56581e-05, 6.456773e-06, 1.297056e-05, 1.985779e-05, 
    1.205459e-05, 1.249748e-05, 1.506318e-05, 1.222107e-05, 8.713091e-06, 
    7.570491e-06, 2.548877e-06, 2.633127e-06, 4.164306e-06, 7.241117e-06,
  4.215604e-05, 5.867104e-05, 4.859871e-05, 2.111079e-05, 1.704838e-05, 
    1.013673e-05, 3.720763e-06, 7.595226e-06, 1.31221e-05, 1.08317e-05, 
    4.622508e-06, 2.653502e-06, 4.980557e-06, 9.705665e-06, 1.286862e-05,
  4.985067e-05, 5.874125e-05, 4.715277e-05, 2.915205e-05, 2.282018e-05, 
    1.78065e-05, 7.377109e-06, 1.013058e-06, 6.100913e-06, 6.53108e-06, 
    4.769706e-06, 5.742393e-06, 6.862619e-06, 7.464476e-06, 1.129112e-05,
  5.913063e-05, 5.685071e-05, 6.094461e-05, 4.285351e-05, 2.732052e-05, 
    2.45806e-05, 1.891126e-05, 5.910363e-06, 2.867641e-06, 9.109681e-06, 
    4.983144e-06, 5.621534e-06, 6.133954e-06, 5.259737e-06, 6.197562e-06,
  6.498343e-05, 6.375746e-05, 5.882223e-05, 4.882981e-05, 4.351318e-05, 
    3.460089e-05, 2.380343e-05, 2.173621e-05, 1.677662e-05, 1.611231e-05, 
    1.217132e-05, 6.104934e-06, 4.256038e-06, 3.864657e-06, 4.077563e-06,
  6.061849e-05, 5.83397e-05, 5.19253e-05, 3.96357e-05, 4.261967e-05, 
    3.593651e-05, 2.970032e-05, 2.215832e-05, 9.681215e-06, 7.725078e-06, 
    9.14928e-06, 6.974675e-06, 4.024774e-06, 2.623807e-06, 1.793547e-06,
  5.212054e-05, 4.839282e-05, 3.844353e-05, 2.842766e-05, 2.241937e-05, 
    2.347956e-05, 2.183919e-05, 1.756183e-05, 1.329128e-05, 1.257055e-05, 
    1.21063e-05, 7.659367e-06, 2.795538e-06, 1.365089e-06, 1.209071e-06,
  2.468251e-05, 1.552409e-05, 1.453626e-05, 1.145001e-05, 1.238339e-05, 
    1.144473e-05, 1.289017e-05, 1.655876e-05, 1.671345e-05, 1.161657e-05, 
    1.112834e-05, 6.342078e-06, 2.297309e-06, 8.388911e-07, 8.596539e-07,
  1.507717e-05, 2.21523e-05, 2.184138e-05, 1.617219e-05, 1.527377e-05, 
    2.615277e-05, 3.239099e-05, 9.393028e-06, 5.632238e-06, 4.47815e-06, 
    9.629677e-06, 1.460721e-05, 1.276595e-05, 1.06459e-05, 6.326707e-06,
  2.451115e-05, 1.10562e-05, 9.463226e-06, 4.538835e-06, 3.050313e-06, 
    2.220774e-05, 4.304878e-05, 1.602754e-05, 2.760082e-06, 7.98937e-06, 
    5.198445e-06, 9.113991e-06, 6.743033e-06, 3.701446e-06, 3.210432e-06,
  4.733371e-05, 1.742376e-05, 7.448386e-06, 3.2636e-06, 2.869447e-06, 
    1.620339e-05, 3.611185e-05, 2.580496e-05, 9.387883e-06, 8.36147e-06, 
    3.604346e-06, 2.418909e-06, 4.368642e-06, 2.312845e-06, 1.912495e-06,
  5.326469e-05, 5.056736e-05, 3.846442e-05, 2.265826e-05, 9.977407e-06, 
    6.248177e-06, 1.885965e-05, 2.168439e-05, 1.821114e-05, 7.73488e-06, 
    2.851864e-06, 6.620654e-07, 2.685503e-06, 2.984616e-06, 3.208592e-06,
  5.550749e-05, 5.289581e-05, 4.268056e-05, 3.637037e-05, 2.937465e-05, 
    1.530157e-05, 2.603641e-06, 4.923012e-06, 1.131974e-05, 4.516426e-06, 
    2.1913e-06, 1.901321e-06, 3.422036e-06, 4.369498e-06, 3.332323e-06,
  5.808794e-05, 5.151614e-05, 4.587306e-05, 4.175426e-05, 3.886547e-05, 
    2.921758e-05, 7.546519e-06, 4.827109e-07, 1.435964e-06, 5.344197e-06, 
    3.883355e-06, 5.548676e-06, 3.704225e-06, 3.37028e-06, 3.378772e-06,
  6.413024e-05, 5.80821e-05, 5.037379e-05, 4.213331e-05, 3.820646e-05, 
    3.44857e-05, 2.365046e-05, 1.115417e-05, 5.242963e-06, 9.307096e-06, 
    5.236863e-06, 4.746805e-06, 3.241744e-06, 2.128623e-06, 5.349939e-06,
  6.624966e-05, 5.632803e-05, 4.584897e-05, 3.632365e-05, 3.624291e-05, 
    2.793498e-05, 2.053448e-05, 1.389285e-05, 1.867077e-06, 1.920125e-06, 
    3.949694e-06, 2.118148e-06, 2.696506e-06, 5.447984e-06, 7.45973e-06,
  3.200039e-05, 3.980783e-05, 3.768355e-05, 2.587813e-05, 1.457905e-05, 
    1.50246e-05, 1.127121e-05, 5.598314e-06, 1.778315e-06, 7.897085e-07, 
    1.793589e-06, 3.383428e-06, 6.12664e-06, 6.188542e-06, 4.860869e-06,
  9.571145e-06, 1.595594e-05, 1.702411e-05, 9.682951e-06, 2.84143e-06, 
    1.869138e-06, 2.1484e-06, 5.929905e-06, 3.247972e-06, 1.232803e-06, 
    2.064168e-06, 3.155228e-06, 4.013461e-06, 2.266824e-06, 1.275988e-06,
  1.90656e-06, 2.003751e-06, 1.018725e-06, 2.239429e-06, 1.451484e-06, 
    3.360807e-06, 8.148457e-06, 1.06938e-05, 4.189583e-06, 4.392552e-07, 
    1.920342e-06, 9.405805e-06, 1.079723e-05, 1.440727e-05, 2.117596e-05,
  9.904272e-06, 2.990836e-06, 1.010896e-06, 1.758977e-06, 5.391896e-06, 
    1.22032e-05, 1.826765e-05, 6.96155e-06, 9.829089e-07, 4.515972e-06, 
    6.557453e-06, 1.792756e-05, 1.987769e-05, 1.571243e-05, 1.703798e-05,
  3.413814e-05, 2.227202e-05, 1.417289e-05, 9.903154e-06, 7.322018e-06, 
    1.020702e-05, 8.733945e-06, 5.772662e-06, 3.111963e-06, 6.050629e-06, 
    1.040681e-05, 1.544972e-05, 2.056474e-05, 1.873644e-05, 1.493008e-05,
  5.845852e-05, 5.14165e-05, 3.352e-05, 2.427579e-05, 1.225598e-05, 
    4.447661e-06, 1.68545e-06, 6.93972e-07, 2.359366e-06, 3.610582e-06, 
    4.617766e-06, 1.005777e-05, 1.699121e-05, 1.778356e-05, 1.655892e-05,
  4.330989e-05, 3.993617e-05, 3.237615e-05, 2.447751e-05, 1.525494e-05, 
    9.187738e-06, 1.218849e-06, 6.438558e-07, 5.909857e-06, 2.077677e-06, 
    3.465787e-06, 7.570029e-06, 1.323985e-05, 1.35977e-05, 1.540051e-05,
  3.179314e-05, 3.38469e-05, 2.824724e-05, 2.150578e-05, 1.868318e-05, 
    1.376341e-05, 7.531445e-06, 3.202227e-06, 1.600003e-06, 9.334111e-06, 
    5.585906e-06, 8.526404e-06, 1.181795e-05, 1.114888e-05, 1.044481e-05,
  2.592294e-05, 2.612079e-05, 2.824623e-05, 2.575485e-05, 2.740987e-05, 
    2.394927e-05, 1.58033e-05, 6.906374e-06, 8.779075e-06, 9.166852e-06, 
    5.299576e-06, 8.980387e-06, 1.132549e-05, 1.089766e-05, 8.183588e-06,
  2.110494e-05, 2.226965e-05, 2.039804e-05, 2.044957e-05, 2.485173e-05, 
    2.345119e-05, 1.78211e-05, 9.977897e-06, 3.889463e-06, 2.120466e-06, 
    1.837756e-06, 4.491058e-06, 6.702468e-06, 9.675072e-06, 9.637094e-06,
  1.723015e-05, 1.922536e-05, 1.782725e-05, 1.737745e-05, 1.128621e-05, 
    1.042554e-05, 1.109574e-05, 3.842024e-06, 8.45639e-07, 6.880022e-07, 
    9.732947e-07, 1.37004e-06, 2.772825e-06, 4.308197e-06, 5.946879e-06,
  1.37263e-05, 1.201134e-05, 8.593532e-06, 5.817982e-06, 3.61721e-06, 
    1.668001e-06, 1.942727e-06, 2.739657e-06, 7.245622e-07, 1.118227e-06, 
    1.433126e-06, 1.687574e-06, 1.922017e-06, 2.686681e-06, 3.417105e-06,
  3.665684e-06, 4.333014e-06, 2.300186e-06, 1.791015e-06, 3.071311e-06, 
    2.787089e-06, 4.904712e-06, 6.914939e-06, 8.894489e-06, 1.672865e-05, 
    3.212727e-05, 4.073312e-05, 3.531041e-05, 2.140876e-05, 8.780714e-06,
  1.103639e-05, 5.803375e-06, 3.823584e-06, 3.506689e-06, 3.525496e-06, 
    2.050121e-06, 2.339445e-06, 2.807609e-06, 5.558122e-06, 1.132388e-05, 
    2.022625e-05, 3.120803e-05, 2.300856e-05, 1.669272e-05, 1.008139e-05,
  1.790405e-05, 9.705592e-06, 8.270405e-06, 2.955152e-06, 2.378204e-06, 
    8.885028e-07, 1.355124e-06, 1.101332e-06, 1.157746e-06, 5.356306e-06, 
    1.060792e-05, 1.72096e-05, 1.731927e-05, 1.335079e-05, 9.006916e-06,
  3.668553e-05, 2.867011e-05, 2.103992e-05, 1.330965e-05, 6.356652e-06, 
    1.415214e-06, 1.289539e-06, 1.282677e-07, 2.474274e-07, 1.79604e-06, 
    4.852363e-06, 8.267999e-06, 1.058319e-05, 9.43846e-06, 6.454365e-06,
  2.199734e-05, 2.303494e-05, 2.114234e-05, 1.645375e-05, 8.761335e-06, 
    8.439891e-06, 4.617186e-06, 1.450117e-06, 3.851993e-06, 8.390465e-07, 
    2.993364e-06, 3.02965e-06, 6.423608e-06, 5.240972e-06, 5.229163e-06,
  1.498516e-05, 1.462722e-05, 1.517373e-05, 1.610392e-05, 1.409507e-05, 
    1.123191e-05, 6.637371e-06, 7.987488e-06, 2.81249e-06, 5.261258e-06, 
    1.232199e-06, 2.353818e-06, 2.817409e-06, 4.353649e-06, 3.768565e-06,
  1.265065e-05, 1.204526e-05, 1.131511e-05, 1.197692e-05, 1.50874e-05, 
    1.43468e-05, 1.191919e-05, 8.814197e-06, 5.475826e-06, 4.818284e-06, 
    2.417963e-06, 3.546363e-06, 3.049285e-06, 2.841323e-06, 3.632918e-06,
  1.040995e-05, 1.144951e-05, 9.238341e-06, 9.449583e-06, 1.179027e-05, 
    1.638896e-05, 1.064452e-05, 7.73827e-06, 1.705226e-06, 1.729792e-06, 
    1.982712e-06, 3.217423e-06, 4.030181e-06, 3.649394e-06, 3.968859e-06,
  9.206597e-06, 1.007361e-05, 1.28317e-05, 1.172311e-05, 6.649374e-06, 
    5.030916e-06, 5.661207e-06, 1.593846e-06, 1.311626e-06, 1.779431e-06, 
    1.404293e-06, 2.503524e-06, 4.846328e-06, 4.891397e-06, 5.668162e-06,
  8.762277e-06, 7.273047e-06, 2.962308e-06, 1.487943e-06, 1.596883e-06, 
    1.883632e-08, 5.962014e-08, 1.290789e-08, 1.64862e-06, 1.903686e-06, 
    1.088639e-06, 1.360305e-06, 3.179612e-06, 5.663256e-06, 6.405639e-06,
  1.151508e-06, 3.640921e-06, 2.037256e-06, 2.336164e-06, 4.992077e-06, 
    3.068752e-06, 5.945686e-06, 7.240499e-06, 2.080856e-05, 2.520629e-05, 
    2.372311e-05, 1.75379e-05, 1.287238e-05, 6.023639e-06, 2.847979e-06,
  2.90139e-06, 1.698479e-06, 2.11424e-06, 2.462057e-06, 1.245741e-06, 
    9.889171e-07, 3.616352e-06, 5.573621e-06, 1.500533e-05, 2.94589e-05, 
    2.423169e-05, 2.240959e-05, 1.515749e-05, 1.6252e-06, 1.654695e-06,
  1.482794e-05, 4.286951e-06, 3.304678e-06, 9.21513e-07, 6.763691e-08, 
    1.506791e-06, 1.237068e-06, 8.940148e-06, 1.852768e-05, 3.569293e-05, 
    2.567393e-05, 2.262839e-05, 1.436363e-05, 9.55047e-07, 5.441113e-07,
  1.601696e-05, 1.426253e-05, 1.236541e-05, 8.107813e-06, 3.733251e-07, 
    1.601662e-06, 1.841193e-06, 2.60516e-06, 7.607234e-06, 2.280499e-05, 
    2.559853e-05, 2.019985e-05, 1.089847e-05, 2.27083e-06, 8.426193e-07,
  1.151882e-05, 5.375689e-06, 6.773046e-06, 8.761472e-06, 5.302788e-06, 
    5.739016e-06, 3.198443e-06, 1.618633e-06, 1.156353e-05, 2.02772e-05, 
    2.370845e-05, 1.735132e-05, 8.649565e-06, 1.470302e-06, 2.71688e-06,
  1.941927e-05, 1.207827e-05, 1.233359e-05, 9.996123e-06, 1.096167e-05, 
    8.947633e-06, 7.215014e-06, 1.079195e-05, 1.920172e-05, 2.337904e-05, 
    1.72624e-05, 1.361703e-05, 6.800018e-06, 1.764848e-06, 1.207859e-06,
  2.692647e-05, 2.738044e-05, 2.344705e-05, 2.413862e-05, 1.917783e-05, 
    9.705392e-06, 9.431326e-06, 1.035796e-05, 1.412705e-05, 1.534571e-05, 
    1.369122e-05, 1.033256e-05, 6.48945e-06, 3.003239e-06, 1.082695e-06,
  2.069416e-05, 2.4089e-05, 2.533751e-05, 2.145389e-05, 1.393524e-05, 
    8.276269e-06, 4.972043e-06, 6.276777e-06, 6.874454e-06, 9.724362e-06, 
    1.008496e-05, 8.258463e-06, 5.874098e-06, 3.851778e-06, 2.461019e-06,
  1.744002e-05, 2.204204e-05, 1.94373e-05, 7.925743e-06, 6.076847e-06, 
    9.228289e-07, 1.007529e-06, 1.333074e-06, 3.913332e-06, 6.861683e-06, 
    6.557375e-06, 5.664885e-06, 4.668766e-06, 3.177769e-06, 3.14949e-06,
  2.043505e-05, 1.995807e-05, 1.685773e-05, 2.874379e-06, 5.098785e-07, 
    6.486128e-08, 2.535454e-08, 4.489933e-07, 1.407638e-06, 2.973362e-06, 
    2.917719e-06, 3.186633e-06, 2.579466e-06, 2.26088e-06, 2.200894e-06,
  3.467455e-06, 2.335257e-06, 3.378676e-06, 2.084284e-06, 3.852399e-06, 
    3.094285e-06, 7.881607e-06, 1.17976e-05, 1.436697e-05, 6.674846e-06, 
    1.379967e-06, 1.699604e-06, 6.531374e-06, 7.166725e-06, 6.274015e-06,
  6.744394e-06, 3.126057e-06, 1.931918e-06, 1.970646e-06, 6.970665e-07, 
    6.772717e-06, 1.866693e-05, 1.87696e-05, 1.26186e-05, 7.815188e-06, 
    4.155255e-06, 3.380988e-06, 4.955246e-06, 5.034762e-06, 5.588744e-06,
  2.000204e-05, 4.789829e-06, 1.61335e-06, 8.871928e-07, 1.08216e-05, 
    3.220479e-05, 2.679425e-05, 2.442425e-05, 1.187514e-05, 8.739311e-06, 
    7.052502e-06, 5.61387e-06, 4.724897e-06, 5.062506e-06, 5.866867e-06,
  3.033933e-05, 1.884449e-05, 1.348785e-05, 1.931524e-05, 3.798205e-05, 
    3.239881e-05, 1.361536e-05, 1.176557e-05, 1.052202e-05, 7.16431e-06, 
    7.52138e-06, 3.125202e-06, 3.472075e-06, 4.382749e-06, 7.49537e-06,
  1.651476e-05, 8.767088e-06, 2.293867e-05, 3.704724e-05, 3.816115e-05, 
    1.557928e-05, 6.46728e-06, 1.001512e-06, 5.18665e-06, 7.001535e-06, 
    4.011131e-06, 2.087812e-06, 2.207265e-06, 2.727512e-06, 7.054235e-06,
  1.87999e-05, 1.637729e-05, 2.223204e-05, 4.913741e-05, 3.88448e-05, 
    1.373545e-05, 9.647176e-06, 8.662489e-06, 8.004344e-06, 4.899833e-06, 
    3.260084e-06, 1.84632e-06, 2.614888e-06, 3.740084e-06, 4.007768e-06,
  2.436882e-05, 1.897019e-05, 3.674007e-05, 4.847477e-05, 3.361295e-05, 
    2.353213e-05, 2.218938e-05, 1.664195e-05, 1.010837e-05, 3.376206e-06, 
    2.29119e-06, 1.748214e-06, 2.387848e-06, 3.692248e-06, 2.406113e-06,
  2.453719e-05, 2.940593e-05, 4.350132e-05, 3.274206e-05, 2.665585e-05, 
    2.530854e-05, 2.210118e-05, 1.355742e-05, 4.567381e-06, 2.59913e-06, 
    2.109627e-06, 2.443178e-06, 2.67146e-06, 3.8536e-06, 3.447851e-06,
  2.433486e-05, 3.350383e-05, 3.195435e-05, 1.179191e-05, 1.083527e-05, 
    1.245766e-05, 1.210979e-05, 5.194849e-06, 3.815383e-06, 2.222991e-06, 
    2.357536e-06, 2.579578e-06, 3.427128e-06, 3.342354e-06, 4.688454e-06,
  2.047907e-05, 2.239933e-05, 1.026245e-05, 4.615849e-06, 5.130528e-06, 
    1.948617e-06, 2.113593e-06, 3.802673e-06, 2.716995e-06, 2.046297e-06, 
    2.315752e-06, 2.082608e-06, 2.111224e-06, 2.423505e-06, 2.400981e-06,
  4.691558e-05, 4.307595e-05, 3.081175e-05, 1.751258e-05, 7.125682e-06, 
    3.614528e-06, 2.651105e-06, 1.267748e-06, 4.228614e-06, 8.231788e-06, 
    8.506322e-06, 8.277048e-06, 1.025133e-05, 1.154524e-05, 1.282026e-05,
  1.756733e-05, 2.033837e-05, 2.599692e-05, 1.999283e-05, 1.23518e-05, 
    5.655928e-06, 2.894732e-06, 4.560548e-06, 8.947231e-06, 1.425795e-05, 
    1.362041e-05, 1.09703e-05, 1.11978e-05, 8.014487e-06, 8.817999e-06,
  1.664507e-05, 9.970067e-06, 1.516947e-05, 1.5178e-05, 1.066515e-05, 
    9.602027e-06, 4.606859e-06, 9.43961e-06, 1.040925e-05, 1.097501e-05, 
    8.69361e-06, 4.461168e-06, 6.306677e-06, 7.254322e-06, 6.584558e-06,
  1.132625e-05, 1.406776e-05, 1.898201e-05, 2.138339e-05, 2.093038e-05, 
    1.098832e-05, 8.977063e-06, 1.114078e-05, 9.647515e-06, 7.294685e-06, 
    2.235081e-06, 1.020009e-06, 4.88368e-06, 5.622652e-06, 5.927773e-06,
  3.1199e-05, 2.809352e-05, 3.063928e-05, 3.093912e-05, 1.756831e-05, 
    8.284223e-06, 5.262346e-06, 4.060782e-06, 7.514525e-06, 2.93576e-06, 
    1.478275e-06, 2.568445e-06, 6.161961e-06, 5.664024e-06, 5.521984e-06,
  4.855455e-05, 4.085842e-05, 3.669698e-05, 3.499665e-05, 2.243068e-05, 
    1.434656e-05, 8.527553e-06, 1.740008e-06, 1.21626e-06, 1.729256e-06, 
    1.697496e-06, 4.724089e-06, 6.091983e-06, 5.356354e-06, 3.906921e-06,
  5.22822e-05, 5.410182e-05, 4.765428e-05, 4.384309e-05, 4.146797e-05, 
    3.434117e-05, 2.30982e-05, 1.24186e-05, 2.982549e-06, 1.330453e-06, 
    4.005004e-06, 4.973072e-06, 4.065983e-06, 3.219603e-06, 1.695328e-06,
  6.350696e-05, 6.299395e-05, 5.824623e-05, 4.982144e-05, 4.912876e-05, 
    4.564021e-05, 1.582497e-05, 1.151509e-05, 1.281836e-06, 2.036919e-06, 
    3.297089e-06, 2.840163e-06, 1.508986e-06, 1.030022e-06, 1.113692e-06,
  7.275477e-05, 6.347682e-05, 5.02268e-05, 3.430249e-05, 2.208066e-05, 
    1.976398e-05, 1.360307e-05, 6.934708e-06, 9.263194e-07, 3.024388e-06, 
    1.918586e-06, 3.165858e-06, 1.7024e-06, 1.51851e-06, 1.586679e-06,
  3.752568e-05, 2.574893e-05, 1.140874e-05, 1.023914e-05, 7.441503e-06, 
    2.663153e-07, 4.028789e-07, 8.191711e-06, 1.192964e-06, 3.268748e-06, 
    2.450213e-06, 1.993654e-06, 2.23649e-06, 2.004477e-06, 1.686122e-06,
  8.933483e-06, 2.509235e-05, 2.781023e-05, 1.689653e-05, 4.706574e-06, 
    1.168286e-06, 1.136177e-06, 8.12252e-07, 6.836239e-07, 4.842211e-07, 
    2.078872e-07, 1.108474e-07, 3.93784e-07, 8.211426e-07, 1.788685e-06,
  7.860543e-06, 1.070956e-05, 2.368824e-05, 2.387819e-05, 1.281845e-05, 
    5.35522e-06, 2.521991e-06, 1.908965e-06, 1.521961e-06, 1.023817e-06, 
    7.325286e-07, 1.211554e-06, 2.386985e-06, 3.339147e-06, 3.838054e-06,
  1.651113e-05, 1.290652e-05, 1.564565e-05, 2.392114e-05, 1.636488e-05, 
    7.290098e-06, 3.879988e-06, 3.294011e-06, 2.375798e-06, 1.513146e-06, 
    1.431852e-06, 2.191663e-06, 5.237232e-06, 7.285252e-06, 8.930862e-06,
  2.317319e-05, 2.500118e-05, 3.11281e-05, 3.300421e-05, 2.330489e-05, 
    6.751255e-06, 5.011928e-06, 3.495034e-06, 2.066569e-06, 1.348494e-06, 
    1.274789e-06, 1.147899e-06, 4.845491e-06, 8.987171e-06, 1.05092e-05,
  3.412975e-05, 3.821254e-05, 5.123162e-05, 3.243583e-05, 2.187504e-05, 
    9.549216e-06, 2.609435e-06, 1.841557e-06, 1.347821e-06, 5.94664e-07, 
    1.05779e-06, 1.072344e-06, 4.364434e-06, 6.331518e-06, 5.757581e-06,
  4.544576e-05, 4.792206e-05, 4.84852e-05, 3.693768e-05, 2.238588e-05, 
    1.303645e-05, 2.925339e-06, 2.108539e-07, 5.27258e-08, 1.922233e-06, 
    8.238027e-07, 1.919228e-06, 3.308294e-06, 3.150513e-06, 3.661055e-06,
  4.896145e-05, 5.367171e-05, 4.274222e-05, 3.600477e-05, 2.98923e-05, 
    1.711189e-05, 8.79493e-06, 4.745412e-06, 2.085059e-06, 1.015055e-06, 
    1.284331e-06, 1.578117e-06, 1.820827e-06, 1.907049e-06, 2.053116e-06,
  5.825617e-05, 5.113159e-05, 4.482604e-05, 4.08915e-05, 3.783337e-05, 
    2.538212e-05, 1.18247e-05, 4.845545e-06, 1.383314e-06, 9.874818e-07, 
    6.476076e-07, 7.417222e-07, 7.252219e-07, 7.542839e-07, 1.157977e-06,
  5.157898e-05, 5.910188e-05, 4.393524e-05, 2.612343e-05, 1.926116e-05, 
    1.601563e-05, 7.362559e-06, 2.967481e-06, 9.800765e-07, 2.920236e-07, 
    5.515444e-07, 6.130683e-07, 5.605029e-07, 5.447444e-07, 3.016456e-07,
  2.719991e-05, 2.185773e-05, 9.702884e-06, 3.410054e-06, 5.963408e-07, 
    1.493662e-06, 1.733193e-07, 1.840566e-06, 7.575222e-07, 4.089921e-07, 
    9.855005e-07, 9.685486e-07, 7.348568e-07, 6.633277e-07, 3.277092e-07,
  2.278139e-06, 6.299737e-06, 1.029713e-05, 1.324107e-05, 1.357707e-05, 
    1.306913e-05, 1.263794e-05, 7.307987e-06, 1.931318e-06, 6.401115e-07, 
    3.295868e-07, 2.213435e-07, 4.396371e-07, 4.731679e-07, 1.07344e-06,
  2.489017e-06, 3.275365e-06, 9.148525e-06, 1.467306e-05, 1.561249e-05, 
    1.172481e-05, 1.245315e-05, 5.897631e-06, 7.50609e-07, 3.335174e-07, 
    4.458052e-07, 7.213084e-07, 5.935049e-07, 1.324982e-06, 2.669978e-06,
  1.317355e-05, 7.975004e-06, 9.71626e-06, 1.694802e-05, 1.235794e-05, 
    4.868827e-06, 7.007438e-06, 3.301629e-06, 7.390067e-07, 3.470305e-07, 
    6.817282e-07, 6.739552e-07, 1.120015e-06, 2.620539e-06, 5.209028e-06,
  3.542606e-05, 2.295579e-05, 2.566222e-05, 2.078235e-05, 1.401216e-05, 
    2.051448e-06, 1.162161e-06, 1.194289e-06, 7.766965e-07, 8.312508e-07, 
    4.575514e-07, 7.439182e-07, 1.153846e-06, 5.505855e-06, 7.104932e-06,
  3.264797e-05, 2.687586e-05, 3.28753e-05, 2.44926e-05, 1.031471e-05, 
    2.859747e-06, 9.670538e-07, 6.632132e-07, 4.195998e-07, 2.789502e-07, 
    4.132827e-07, 4.092286e-07, 2.191326e-06, 2.356798e-06, 4.26302e-06,
  4.050886e-05, 3.61394e-05, 3.264516e-05, 2.638178e-05, 1.411294e-05, 
    5.66096e-06, 8.866497e-07, 1.015861e-07, 4.489445e-08, 1.477463e-07, 
    9.596129e-07, 4.647247e-07, 1.455092e-06, 1.277547e-06, 1.129626e-06,
  4.27583e-05, 4.184149e-05, 3.5837e-05, 2.891089e-05, 1.796569e-05, 
    7.125836e-06, 4.506878e-06, 2.362076e-07, 2.815538e-07, 1.288382e-07, 
    2.578793e-07, 7.105639e-07, 9.035077e-07, 9.787129e-07, 1.25366e-06,
  4.39901e-05, 3.983081e-05, 3.377431e-05, 2.71229e-05, 2.74175e-05, 
    1.809932e-05, 8.397777e-06, 5.287057e-06, 1.370149e-06, 3.292182e-07, 
    7.177838e-07, 7.715793e-07, 8.527622e-07, 8.640694e-07, 1.078835e-06,
  3.639225e-05, 3.835045e-05, 3.297274e-05, 2.48581e-05, 1.927826e-05, 
    1.363823e-05, 5.836133e-06, 8.66894e-07, 8.206516e-07, 8.107176e-07, 
    7.940715e-07, 9.873671e-07, 8.64297e-07, 5.994629e-07, 6.955583e-07,
  2.374634e-05, 1.795555e-05, 4.559719e-06, 5.470313e-07, 7.190997e-07, 
    9.854582e-07, 1.888632e-06, 2.330868e-07, 7.559794e-07, 7.921176e-07, 
    9.610749e-07, 9.794575e-07, 9.216565e-07, 6.287814e-07, 2.139869e-07,
  3.414702e-06, 4.253316e-06, 4.968169e-06, 2.485471e-06, 2.593448e-06, 
    3.652501e-06, 9.497204e-06, 2.141896e-05, 2.088893e-05, 1.507372e-05, 
    9.829269e-06, 7.450378e-06, 3.844262e-06, 1.33201e-06, 7.983639e-07,
  4.228306e-06, 6.424157e-07, 2.049045e-06, 1.960248e-06, 2.148161e-06, 
    3.539635e-06, 2.095309e-05, 2.086486e-05, 1.411998e-05, 9.952053e-06, 
    3.071206e-06, 1.507307e-06, 5.117121e-07, 3.115979e-07, 5.222121e-07,
  1.028885e-05, 5.076567e-06, 3.955885e-06, 1.787723e-06, 2.401529e-06, 
    2.626703e-06, 1.269648e-05, 1.571622e-05, 7.588694e-06, 2.506649e-06, 
    2.748141e-07, 1.461297e-07, 3.629722e-08, 4.760994e-07, 1.831054e-06,
  1.927155e-05, 2.137852e-05, 1.740783e-05, 1.040741e-05, 6.511628e-06, 
    4.359419e-06, 1.794339e-06, 2.476348e-06, 1.684982e-06, 9.212746e-07, 
    4.127372e-07, 1.691219e-07, 4.566498e-07, 1.470242e-06, 2.875555e-06,
  2.269331e-05, 2.283902e-05, 2.232342e-05, 1.633655e-05, 3.803068e-06, 
    5.470489e-06, 5.348087e-07, 5.13353e-08, 2.427896e-07, 4.690617e-07, 
    9.07686e-07, 7.496168e-07, 3.784905e-07, 1.424032e-06, 3.100979e-06,
  2.321537e-05, 2.57975e-05, 2.488574e-05, 1.374734e-05, 6.894581e-06, 
    1.255e-06, 1.893534e-07, 3.297451e-09, 2.608452e-08, 8.623273e-07, 
    7.593064e-07, 5.268296e-07, 8.501927e-07, 3.089616e-07, 2.4658e-06,
  2.283913e-05, 2.508023e-05, 2.443865e-05, 1.969748e-05, 1.116366e-05, 
    4.30336e-06, 1.073895e-06, 1.393383e-06, 8.314694e-07, 4.283274e-07, 
    8.506993e-08, 3.509772e-07, 3.052202e-07, 8.064145e-07, 4.774596e-07,
  2.209625e-05, 2.691289e-05, 2.436774e-05, 2.12846e-05, 2.042689e-05, 
    1.177073e-05, 8.773084e-06, 3.055498e-06, 1.084705e-06, 3.381583e-07, 
    3.253494e-07, 3.554684e-07, 4.209214e-07, 5.49119e-07, 3.412595e-07,
  3.097482e-05, 3.096693e-05, 2.77431e-05, 2.510835e-05, 1.742223e-05, 
    1.013482e-05, 6.33829e-06, 2.190515e-06, 1.423391e-06, 8.91169e-07, 
    6.535089e-07, 7.220158e-07, 7.711855e-07, 5.584062e-07, 6.369968e-07,
  3.810339e-05, 3.637878e-05, 1.338626e-05, 1.146227e-06, 5.698261e-07, 
    8.214113e-07, 2.259204e-06, 1.501404e-06, 6.813667e-07, 6.505707e-07, 
    9.564334e-07, 7.144233e-07, 6.165907e-07, 4.62242e-07, 3.309516e-07,
  2.229688e-06, 4.099081e-06, 2.895998e-06, 1.994349e-06, 7.308973e-07, 
    1.218212e-06, 3.159109e-06, 4.894784e-06, 5.373329e-06, 3.346826e-06, 
    1.664645e-06, 1.627435e-06, 2.075956e-06, 8.716909e-07, 1.159128e-06,
  4.707055e-06, 1.250511e-06, 1.893235e-06, 1.046368e-06, 5.370115e-07, 
    8.706325e-07, 3.506557e-06, 4.445576e-06, 4.296523e-06, 4.798381e-06, 
    1.426178e-06, 8.358986e-07, 4.657297e-07, 1.953667e-07, 2.488336e-07,
  1.076287e-05, 4.015008e-06, 2.543728e-06, 7.744647e-07, 4.706827e-07, 
    1.501431e-07, 8.337095e-07, 2.566989e-06, 2.184829e-06, 1.232051e-06, 
    1.403627e-06, 3.675111e-07, 2.569194e-07, 1.855808e-07, 8.592108e-07,
  1.7491e-05, 1.405089e-05, 9.990049e-06, 3.990743e-06, 4.921109e-07, 
    1.58562e-07, 3.108452e-07, 5.197024e-07, 3.19141e-07, 1.399898e-06, 
    1.315075e-06, 1.09347e-06, 1.671676e-06, 2.347505e-06, 4.099407e-07,
  2.337597e-05, 1.931214e-05, 1.639929e-05, 5.677717e-06, 3.446192e-08, 
    1.17116e-07, 4.594254e-08, 8.878649e-08, 1.321249e-06, 1.781677e-06, 
    1.542589e-06, 1.072241e-06, 1.373e-06, 1.504574e-06, 1.990978e-06,
  3.09816e-05, 1.950466e-05, 1.686775e-05, 1.028955e-05, 4.048681e-06, 
    2.61841e-06, 2.045805e-06, 2.438496e-06, 1.745914e-06, 2.084689e-06, 
    1.010736e-06, 6.533656e-07, 9.539676e-07, 4.489558e-07, 1.400674e-06,
  3.389299e-05, 2.406127e-05, 1.979958e-05, 1.807578e-05, 1.408929e-05, 
    1.27768e-05, 4.012485e-06, 2.416852e-06, 1.956221e-06, 1.799412e-06, 
    1.117455e-06, 9.632171e-07, 8.324523e-07, 4.95639e-07, 4.12246e-07,
  3.380329e-05, 3.166603e-05, 2.423289e-05, 1.964312e-05, 2.469109e-05, 
    1.73292e-05, 1.007946e-05, 2.753512e-06, 1.813749e-06, 8.266804e-07, 
    8.981982e-07, 1.162662e-06, 1.121155e-06, 8.525396e-07, 1.148381e-06,
  2.959201e-05, 3.332751e-05, 3.091682e-05, 2.337055e-05, 1.795414e-05, 
    1.075573e-05, 3.894243e-06, 1.882529e-06, 1.960933e-06, 6.494491e-07, 
    6.764088e-07, 9.790483e-07, 1.253062e-06, 1.187013e-06, 1.949341e-06,
  2.845599e-05, 2.672494e-05, 4.397818e-06, 3.922944e-06, 1.801196e-06, 
    1.585691e-06, 9.717656e-07, 1.758854e-06, 6.717023e-07, 5.103592e-07, 
    7.375048e-07, 6.563591e-07, 7.299367e-07, 8.086366e-07, 9.090737e-07,
  5.809568e-06, 4.087439e-06, 2.774716e-06, 2.119651e-06, 1.317067e-06, 
    6.140615e-07, 6.466643e-07, 5.361229e-07, 3.52975e-07, 1.721379e-07, 
    2.948648e-07, 1.964983e-07, 5.846107e-07, 4.498428e-07, 6.555498e-07,
  3.933382e-06, 1.334871e-06, 1.154554e-06, 1.826267e-06, 3.348599e-07, 
    1.722632e-07, 1.42491e-07, 3.283332e-07, 3.141062e-07, 9.264447e-07, 
    1.700607e-07, 9.190904e-08, 3.958489e-07, 2.480575e-07, 2.108914e-07,
  6.905189e-06, 2.827781e-06, 1.645036e-06, 1.122858e-06, 5.927272e-07, 
    2.438546e-07, 1.78902e-07, 4.503198e-07, 4.678782e-07, 6.199394e-07, 
    5.409112e-07, 5.653649e-07, 8.302437e-07, 6.872815e-07, 2.549461e-07,
  1.52603e-05, 1.164257e-05, 8.854139e-06, 6.370071e-06, 3.575092e-06, 
    2.792135e-07, 4.830258e-07, 5.20588e-07, 5.032426e-07, 1.061719e-07, 
    4.855278e-07, 5.330878e-07, 1.061891e-06, 8.577397e-07, 6.468526e-07,
  1.959613e-05, 1.712739e-05, 1.577334e-05, 1.15842e-05, 1.277221e-07, 
    3.450918e-06, 1.037262e-06, 4.351475e-07, 6.124787e-07, 8.772062e-07, 
    5.227411e-07, 2.840709e-07, 1.111696e-06, 1.290544e-06, 2.202974e-06,
  2.314723e-05, 1.812664e-05, 1.618189e-05, 1.24041e-05, 7.872067e-06, 
    3.499266e-06, 2.422338e-06, 2.70616e-06, 1.412963e-06, 2.66292e-06, 
    1.04402e-06, 7.373698e-07, 6.488388e-07, 1.008601e-06, 1.090938e-06,
  3.024438e-05, 1.824765e-05, 2.015715e-05, 1.969e-05, 1.807663e-05, 
    1.196534e-05, 3.714676e-06, 2.651365e-06, 2.778905e-06, 2.361074e-06, 
    1.669692e-06, 1.031361e-06, 4.454437e-07, 4.6057e-07, 1.679271e-07,
  3.428408e-05, 2.354149e-05, 2.319416e-05, 2.078432e-05, 2.019322e-05, 
    1.514352e-05, 8.483341e-06, 2.662222e-06, 2.231855e-06, 1.720883e-06, 
    1.752183e-06, 1.453893e-06, 6.731636e-07, 4.37937e-07, 2.127566e-07,
  3.248472e-05, 2.735995e-05, 2.971741e-05, 1.979996e-05, 1.31354e-05, 
    9.044379e-06, 3.58424e-06, 2.661619e-06, 2.550254e-06, 1.756897e-06, 
    1.328713e-06, 1.147801e-06, 1.074435e-06, 4.707385e-07, 6.734886e-08,
  3.033988e-05, 1.313729e-05, 5.996134e-06, 3.119784e-06, 2.199662e-06, 
    2.35879e-06, 2.841597e-06, 2.675009e-06, 1.444954e-06, 9.266566e-07, 
    8.399709e-07, 5.681823e-07, 5.203959e-07, 2.830384e-07, 8.893672e-08,
  1.198659e-05, 1.98838e-05, 2.394551e-05, 2.525161e-05, 2.313836e-05, 
    1.930085e-05, 1.603508e-05, 1.109463e-05, 6.074131e-06, 2.27829e-06, 
    7.707893e-07, 2.751254e-07, 2.833386e-07, 1.570762e-07, 2.979888e-07,
  5.007153e-06, 5.266357e-06, 6.75067e-06, 8.34589e-06, 5.259332e-06, 
    4.144538e-06, 4.179273e-06, 2.420898e-06, 8.920208e-07, 7.550473e-07, 
    2.783318e-07, 8.846528e-08, 6.578352e-09, 3.911628e-07, 5.277763e-07,
  9.252285e-06, 3.141567e-06, 2.722941e-06, 3.283577e-06, 1.835873e-06, 
    5.964416e-07, 1.030166e-06, 9.955653e-07, 5.080336e-07, 4.105086e-08, 
    2.475572e-07, 3.197083e-07, 4.512859e-07, 3.60369e-08, 4.531787e-07,
  2.086224e-05, 1.795343e-05, 1.104268e-05, 4.377793e-06, 2.001781e-06, 
    2.600204e-06, 5.446585e-07, 4.743996e-07, 5.484594e-07, 3.456824e-07, 
    6.474711e-08, 3.39053e-07, 1.645353e-08, 2.427249e-07, 8.183169e-07,
  2.358494e-05, 2.127078e-05, 1.856041e-05, 1.299608e-05, 3.869291e-08, 
    3.048865e-06, 2.596223e-06, 7.335164e-07, 3.872864e-07, 2.410918e-07, 
    3.683124e-07, 2.221854e-07, 1.606563e-07, 5.959909e-07, 7.414725e-07,
  1.963389e-05, 1.617664e-05, 1.637152e-05, 1.094039e-05, 7.164296e-06, 
    1.10812e-06, 3.16994e-06, 1.074135e-06, 4.665639e-09, 1.207409e-07, 
    3.508936e-07, 2.57543e-07, 2.900785e-07, 8.183646e-08, 2.258773e-08,
  2.304129e-05, 1.505641e-05, 1.544996e-05, 1.250042e-05, 1.384463e-05, 
    1.107842e-05, 4.041509e-06, 1.828053e-06, 1.10304e-06, 4.072631e-07, 
    1.014642e-07, 1.20191e-07, 2.441663e-07, 4.906233e-07, 8.885134e-08,
  2.863199e-05, 2.504204e-05, 2.440547e-05, 1.733676e-05, 1.915041e-05, 
    1.581932e-05, 8.459705e-06, 1.740535e-06, 7.63945e-07, 1.938883e-07, 
    1.403715e-07, 1.501356e-07, 2.600847e-07, 4.542035e-07, 6.536509e-07,
  1.910925e-05, 2.003335e-05, 2.392938e-05, 1.789904e-05, 1.537679e-05, 
    9.70657e-06, 3.306081e-06, 1.376015e-06, 3.600571e-07, 2.70637e-07, 
    1.787649e-07, 3.308938e-07, 7.725192e-07, 1.177078e-06, 1.001646e-06,
  2.018858e-05, 2.038868e-05, 9.464126e-06, 3.956206e-06, 3.187581e-06, 
    1.883678e-06, 7.847332e-07, 4.043358e-07, 2.794567e-07, 3.407937e-07, 
    8.426778e-07, 2.470072e-06, 5.963811e-06, 1.058871e-05, 1.278093e-05,
  2.247338e-05, 5.497442e-05, 6.487512e-05, 7.69682e-05, 8.256343e-05, 
    7.477737e-05, 6.342655e-05, 5.135422e-05, 3.873288e-05, 2.527641e-05, 
    1.710361e-05, 1.519041e-05, 1.542377e-05, 1.408392e-05, 1.108349e-05,
  9.481085e-06, 2.200011e-05, 3.813907e-05, 5.656371e-05, 4.951813e-05, 
    4.482274e-05, 5.206445e-05, 3.889872e-05, 2.717896e-05, 1.795305e-05, 
    9.519747e-06, 9.343456e-06, 9.176719e-06, 7.903537e-06, 5.73744e-06,
  7.394661e-06, 4.39625e-06, 7.5491e-06, 1.060352e-05, 9.747168e-06, 
    1.025674e-05, 1.297766e-05, 1.475848e-05, 1.169604e-05, 6.820172e-06, 
    3.730247e-06, 2.455343e-06, 2.949311e-06, 3.422921e-06, 1.908014e-06,
  2.520586e-05, 1.878973e-05, 8.879405e-06, 3.700886e-06, 2.858244e-06, 
    2.055236e-06, 1.744975e-06, 1.909014e-06, 1.527687e-06, 1.802853e-06, 
    4.403115e-07, 2.051673e-07, 2.914799e-07, 6.226022e-07, 4.439495e-07,
  1.898505e-05, 2.216171e-05, 1.80613e-05, 8.048169e-06, 1.369201e-06, 
    1.599058e-06, 7.491616e-07, 2.314609e-07, 3.650434e-07, 6.357157e-07, 
    5.888836e-07, 7.834977e-07, 4.875553e-08, 5.657664e-09, 9.695563e-09,
  1.072721e-05, 1.386127e-05, 1.679449e-05, 1.042802e-05, 7.003775e-06, 
    1.049008e-06, 2.503493e-06, 4.17013e-07, 3.342607e-09, 3.530589e-07, 
    4.349263e-07, 5.111453e-07, 1.071795e-07, 2.872376e-08, 2.465306e-08,
  9.419412e-06, 4.052482e-06, 8.765036e-06, 1.160826e-05, 1.461285e-05, 
    8.948038e-06, 2.996527e-06, 9.173634e-07, 3.962265e-07, 3.642869e-07, 
    2.724397e-07, 1.020833e-07, 2.60515e-07, 7.341396e-07, 2.290924e-07,
  4.530495e-05, 1.59008e-05, 1.415644e-05, 1.573885e-05, 1.253798e-05, 
    1.221583e-05, 3.821303e-06, 6.295296e-07, 1.361731e-07, 3.761324e-07, 
    3.160394e-07, 3.713703e-07, 5.458016e-07, 5.199722e-07, 2.418919e-07,
  6.979654e-05, 5.408105e-05, 4.486703e-05, 3.237692e-05, 8.748232e-06, 
    5.132181e-06, 1.53119e-06, 1.433282e-06, 2.131558e-06, 3.131672e-06, 
    3.593023e-06, 4.065197e-06, 4.4706e-06, 3.692668e-06, 1.482655e-06,
  1.86878e-05, 2.828561e-05, 1.496186e-05, 1.251759e-06, 9.543738e-07, 
    4.161297e-06, 8.768383e-06, 1.226116e-05, 1.319164e-05, 1.749725e-05, 
    2.570595e-05, 3.276149e-05, 3.288817e-05, 2.477531e-05, 1.11593e-05,
  2.084849e-06, 1.713065e-05, 4.200431e-05, 7.705107e-05, 9.335952e-05, 
    7.666548e-05, 6.117464e-05, 5.001589e-05, 3.914263e-05, 2.600627e-05, 
    2.519197e-05, 3.721104e-05, 4.363648e-05, 3.65191e-05, 2.795077e-05,
  6.899076e-07, 4.683283e-06, 1.743525e-05, 5.876632e-05, 8.204049e-05, 
    6.83589e-05, 7.762278e-05, 5.677858e-05, 4.182164e-05, 3.146217e-05, 
    2.414873e-05, 3.524589e-05, 4.080439e-05, 3.544439e-05, 3.318064e-05,
  7.414491e-06, 1.879704e-06, 5.034423e-06, 1.118701e-05, 1.527519e-05, 
    1.626297e-05, 1.957157e-05, 3.794494e-05, 3.546348e-05, 2.695273e-05, 
    2.136301e-05, 2.85413e-05, 3.992558e-05, 4.421669e-05, 3.575453e-05,
  1.807606e-05, 1.947175e-05, 8.966237e-06, 3.396979e-06, 3.666546e-06, 
    2.877337e-06, 9.36874e-07, 1.392501e-06, 3.865251e-06, 1.307741e-05, 
    1.169614e-05, 1.417179e-05, 2.093745e-05, 2.615259e-05, 2.291756e-05,
  1.794967e-05, 1.560407e-05, 1.489286e-05, 2.660413e-06, 6.389815e-07, 
    5.870043e-07, 1.258894e-07, 1.792656e-08, 3.345789e-07, 1.248027e-06, 
    2.685251e-06, 3.957063e-06, 5.737561e-06, 7.505084e-06, 1.050662e-05,
  2.325135e-05, 1.570479e-05, 9.888739e-06, 6.826252e-06, 1.134057e-06, 
    3.516849e-07, 1.920114e-07, 1.131516e-08, 1.112802e-07, 6.783527e-08, 
    6.424603e-07, 7.72041e-07, 1.426232e-06, 2.261329e-06, 3.774397e-06,
  6.708279e-05, 2.538239e-05, 5.237781e-06, 1.028744e-05, 1.170444e-05, 
    6.63607e-06, 1.957796e-07, 9.655134e-09, 7.109553e-08, 4.26839e-07, 
    2.15741e-07, 3.535022e-07, 8.95669e-07, 1.277151e-06, 1.180052e-06,
  7.299881e-05, 3.473553e-05, 2.504417e-05, 1.519707e-05, 7.840908e-06, 
    6.418344e-06, 4.713171e-06, 8.214049e-07, 3.246736e-06, 2.761902e-06, 
    1.13395e-06, 3.340384e-07, 5.39261e-07, 6.717866e-07, 9.250273e-07,
  3.027802e-05, 2.613423e-05, 2.084891e-05, 8.61244e-06, 5.619894e-06, 
    7.22531e-06, 5.875721e-06, 5.63458e-06, 7.545102e-06, 1.264743e-05, 
    1.551386e-05, 1.106167e-05, 3.558099e-06, 9.614512e-07, 7.888593e-07,
  1.371416e-05, 8.144068e-06, 3.897225e-06, 3.098846e-06, 4.167006e-06, 
    7.992925e-06, 9.559688e-06, 7.896024e-06, 7.845911e-06, 1.043459e-05, 
    1.651973e-05, 2.220478e-05, 1.904536e-05, 9.423285e-06, 3.337988e-06,
  3.704431e-07, 4.745986e-07, 1.317223e-06, 7.916789e-06, 2.035666e-05, 
    2.179884e-05, 1.691894e-05, 7.042021e-06, 5.420142e-06, 9.143184e-06, 
    1.215574e-05, 1.140678e-05, 7.168139e-06, 4.33764e-06, 4.028371e-06,
  6.840273e-07, 5.98123e-07, 5.953858e-07, 3.650065e-06, 9.324032e-06, 
    1.166197e-05, 1.715612e-05, 1.942563e-05, 1.613294e-05, 1.712916e-05, 
    1.913247e-05, 1.909018e-05, 1.490773e-05, 7.361266e-06, 6.403727e-06,
  1.610424e-06, 1.360959e-06, 8.334713e-07, 1.411829e-06, 1.889955e-06, 
    1.818362e-06, 5.473657e-06, 1.924984e-05, 2.553122e-05, 2.345994e-05, 
    2.095543e-05, 2.172812e-05, 2.185604e-05, 1.942151e-05, 1.711482e-05,
  2.657823e-06, 1.163094e-05, 1.106097e-05, 1.180364e-06, 1.339177e-06, 
    1.161123e-06, 6.607388e-07, 2.140319e-06, 4.202658e-06, 1.072971e-05, 
    1.428911e-05, 1.588159e-05, 2.068638e-05, 2.593094e-05, 2.30701e-05,
  1.463285e-06, 7.435142e-06, 1.028162e-05, 2.781951e-06, 1.697861e-06, 
    1.849492e-06, 4.553574e-07, 2.628965e-08, 8.446047e-08, 5.514052e-07, 
    2.276698e-06, 3.949911e-06, 1.035331e-05, 1.654339e-05, 2.468448e-05,
  4.537449e-06, 1.475776e-05, 3.355188e-06, 5.237712e-06, 3.28806e-06, 
    2.463152e-06, 2.164488e-06, 1.962705e-07, 4.130217e-08, 1.167604e-07, 
    2.247622e-07, 2.86492e-07, 8.793272e-07, 4.681766e-06, 1.590597e-05,
  1.628279e-05, 1.520209e-05, 7.974718e-06, 3.069415e-06, 7.452529e-06, 
    3.984482e-06, 2.885123e-06, 1.277442e-06, 2.732253e-06, 8.536127e-07, 
    6.245489e-08, 9.433543e-08, 3.540201e-07, 1.152044e-06, 3.422219e-06,
  1.596676e-05, 1.990455e-05, 1.422348e-05, 7.092973e-06, 9.88748e-06, 
    9.243703e-06, 3.638552e-06, 2.219278e-06, 2.465634e-06, 2.974081e-06, 
    8.812981e-07, 9.321166e-08, 2.152305e-07, 6.0433e-07, 1.266203e-06,
  1.63579e-05, 2.274414e-05, 1.877287e-05, 4.629973e-06, 4.101745e-06, 
    2.192974e-06, 9.597397e-07, 8.791233e-09, 1.28773e-06, 1.745118e-06, 
    6.535606e-07, 7.478744e-07, 1.061108e-06, 4.86961e-07, 6.49579e-07,
  1.640768e-05, 1.599999e-05, 6.777202e-06, 2.612357e-06, 1.126879e-06, 
    7.716174e-07, 5.424218e-07, 9.212624e-09, 8.073079e-07, 1.296904e-06, 
    8.764292e-07, 7.961344e-07, 1.5584e-06, 1.588168e-06, 1.045431e-06,
  3.738094e-06, 1.743475e-06, 1.042703e-06, 1.043415e-06, 2.828069e-07, 
    2.373975e-07, 6.905639e-07, 2.683772e-06, 3.301845e-06, 4.560316e-06, 
    4.164035e-06, 3.677985e-06, 3.432438e-06, 1.341483e-06, 1.420442e-06,
  5.080967e-06, 2.454479e-06, 1.739459e-06, 1.17977e-06, 1.343112e-06, 
    6.679763e-07, 4.782628e-07, 1.866478e-07, 1.936055e-06, 3.974634e-06, 
    4.991648e-06, 5.164352e-06, 4.971861e-06, 5.041555e-06, 3.550169e-06,
  5.735102e-06, 3.245739e-06, 2.443895e-06, 1.704405e-06, 1.171373e-06, 
    2.930367e-06, 8.104163e-07, 5.370582e-07, 5.949875e-07, 1.430944e-06, 
    1.819624e-06, 3.924525e-06, 4.507045e-06, 5.287633e-06, 4.351044e-06,
  1.694653e-05, 8.987953e-06, 3.809652e-06, 2.025714e-06, 1.068555e-06, 
    7.67241e-07, 2.682374e-06, 7.363229e-07, 1.734278e-07, 3.500582e-07, 
    8.930646e-07, 2.510007e-07, 1.255146e-06, 2.573346e-06, 4.726818e-06,
  2.656949e-05, 1.870987e-05, 1.225796e-05, 3.214316e-06, 1.615452e-06, 
    1.451653e-06, 1.526284e-06, 3.154029e-06, 4.373047e-07, 2.639032e-07, 
    2.244248e-07, 3.24726e-07, 3.411205e-07, 2.503605e-07, 2.405729e-06,
  4.325556e-05, 3.100582e-05, 1.942591e-05, 9.368125e-06, 1.448506e-06, 
    2.325952e-06, 2.561251e-06, 1.654121e-06, 7.066637e-07, 3.104794e-07, 
    1.272527e-07, 3.308991e-08, 2.009311e-07, 2.104369e-07, 7.750074e-07,
  4.645477e-05, 4.379969e-05, 2.831888e-05, 1.118861e-05, 5.660671e-06, 
    4.310426e-06, 3.789582e-06, 2.006663e-06, 1.65986e-06, 1.502262e-06, 
    1.634783e-07, 9.395175e-09, 9.084583e-08, 1.703691e-07, 4.076244e-07,
  4.470369e-05, 4.100278e-05, 3.02665e-05, 1.437437e-05, 1.345012e-05, 
    1.494728e-05, 4.416102e-06, 2.119628e-06, 1.713269e-06, 2.368293e-06, 
    1.032276e-06, 2.282564e-08, 6.386973e-08, 7.896102e-08, 2.208626e-08,
  4.248709e-05, 3.833165e-05, 2.842392e-05, 1.166927e-05, 6.550031e-06, 
    2.537269e-06, 2.158926e-06, 2.095207e-06, 2.135181e-06, 1.357547e-06, 
    1.077097e-06, 2.94852e-07, 5.689801e-08, 7.476635e-08, 4.239399e-08,
  3.878346e-05, 3.295146e-05, 1.082113e-05, 3.138174e-06, 2.218989e-06, 
    2.335668e-06, 3.120203e-06, 3.124299e-06, 1.790188e-06, 1.686173e-06, 
    1.486743e-06, 5.510808e-07, 7.737781e-08, 1.003662e-07, 7.487069e-08,
  1.002261e-05, 1.300508e-05, 2.123673e-05, 2.415569e-05, 1.54745e-05, 
    6.550293e-06, 2.761349e-06, 1.942022e-06, 3.137825e-06, 5.349551e-06, 
    6.510968e-06, 6.274766e-06, 4.432273e-06, 2.20082e-06, 2.459282e-06,
  7.809961e-06, 7.152735e-06, 1.258237e-05, 1.781876e-05, 1.386598e-05, 
    4.991332e-06, 2.108462e-06, 1.511657e-06, 1.234424e-06, 2.690159e-06, 
    3.328312e-06, 6.128702e-06, 3.912153e-06, 3.254523e-06, 3.453968e-06,
  5.763479e-06, 6.282279e-06, 8.341337e-06, 1.417084e-05, 1.026841e-05, 
    4.502827e-06, 1.904857e-06, 1.394821e-06, 7.519715e-07, 6.138328e-07, 
    8.53786e-07, 1.053163e-06, 1.933304e-06, 4.08877e-06, 2.012356e-06,
  1.691516e-05, 1.123402e-05, 1.014305e-05, 1.219704e-05, 1.039716e-05, 
    4.706012e-06, 3.910392e-06, 1.535459e-06, 8.194655e-07, 2.993788e-07, 
    2.456751e-07, 2.466351e-07, 4.577115e-07, 7.192464e-07, 4.716583e-07,
  2.213007e-05, 1.886514e-05, 1.731329e-05, 1.36614e-05, 1.020585e-05, 
    7.483199e-06, 4.296412e-06, 5.258951e-06, 3.344277e-06, 9.270949e-07, 
    2.851637e-07, 8.894482e-08, 1.595475e-07, 3.239537e-07, 6.779746e-07,
  3.355317e-05, 2.749858e-05, 1.550251e-05, 1.542412e-05, 1.05349e-05, 
    6.560779e-06, 5.324903e-06, 5.658895e-06, 2.961576e-06, 4.083936e-07, 
    3.699186e-07, 1.112359e-07, 1.207115e-07, 3.015309e-07, 5.515066e-07,
  5.636282e-05, 4.732815e-05, 3.24291e-05, 1.37804e-05, 1.46927e-05, 
    9.929533e-06, 4.060797e-06, 4.736636e-06, 2.885778e-06, 1.957268e-06, 
    7.909385e-07, 1.058534e-07, 3.232547e-08, 9.238666e-08, 2.767914e-07,
  5.332501e-05, 5.166496e-05, 3.715577e-05, 1.888223e-05, 1.871002e-05, 
    1.891944e-05, 3.759762e-06, 4.143548e-06, 2.545458e-06, 2.43444e-06, 
    1.335827e-06, 7.035648e-07, 1.798498e-07, 1.270514e-07, 1.465116e-08,
  2.853686e-05, 3.322267e-05, 3.33967e-05, 1.998371e-05, 1.636182e-05, 
    6.128267e-06, 4.548167e-06, 3.666117e-06, 2.183562e-06, 2.676299e-06, 
    1.509904e-06, 1.102972e-06, 1.519856e-07, 1.951129e-07, 5.717125e-08,
  2.032275e-05, 1.794341e-05, 9.37396e-06, 5.72431e-06, 5.376611e-06, 
    5.018314e-06, 5.249626e-06, 4.95162e-06, 2.188923e-06, 2.344216e-06, 
    2.241896e-06, 5.431074e-07, 1.972284e-07, 2.454506e-07, 1.991233e-07,
  3.918236e-06, 1.630734e-06, 3.278267e-06, 4.753313e-06, 8.10136e-06, 
    1.138696e-05, 1.750577e-05, 2.758828e-05, 3.171087e-05, 2.547738e-05, 
    1.640234e-05, 9.914282e-06, 4.78198e-06, 4.815191e-06, 3.059838e-06,
  2.262394e-06, 1.810061e-06, 2.392478e-06, 4.806646e-06, 7.15236e-06, 
    7.795821e-06, 1.587894e-05, 2.156379e-05, 2.236606e-05, 2.144505e-05, 
    1.38785e-05, 1.129622e-05, 5.472916e-06, 1.188586e-06, 3.473401e-06,
  2.597837e-06, 1.629152e-06, 3.686995e-06, 7.268598e-06, 5.699285e-06, 
    5.544183e-06, 1.057216e-05, 2.014336e-05, 2.144018e-05, 1.782343e-05, 
    1.286005e-05, 7.17363e-06, 4.262272e-06, 2.161533e-06, 5.391542e-07,
  1.145168e-05, 1.063569e-05, 6.393755e-06, 7.335982e-06, 7.550377e-06, 
    8.438966e-06, 6.657797e-06, 1.210788e-05, 1.51401e-05, 1.573932e-05, 
    9.370006e-06, 3.639532e-06, 1.632167e-06, 6.097247e-07, 5.247261e-08,
  1.447172e-05, 1.63811e-05, 1.436229e-05, 9.578325e-06, 5.726391e-06, 
    9.332061e-06, 8.870295e-06, 2.113522e-06, 1.974792e-06, 6.726129e-06, 
    4.410128e-06, 1.299115e-06, 5.946002e-07, 9.163808e-08, 1.517707e-08,
  1.899771e-05, 2.01811e-05, 1.631627e-05, 1.375128e-05, 7.469602e-06, 
    5.668726e-06, 1.04996e-05, 9.880395e-06, 6.402741e-06, 4.209071e-06, 
    1.695805e-06, 9.293067e-07, 2.6313e-07, 2.436168e-08, 1.430506e-08,
  1.751487e-05, 2.947107e-05, 1.515043e-05, 1.36219e-05, 1.495119e-05, 
    1.136922e-05, 7.382664e-06, 9.621207e-06, 7.170947e-06, 4.246391e-06, 
    1.752399e-06, 5.644319e-07, 2.056386e-07, 2.396253e-07, 1.094312e-08,
  1.305878e-05, 2.340616e-05, 1.357658e-05, 1.341585e-05, 2.000244e-05, 
    1.952168e-05, 7.884069e-06, 5.205297e-06, 3.8424e-06, 2.802563e-06, 
    1.833672e-06, 8.567601e-07, 2.909796e-07, 2.200761e-07, 4.179592e-09,
  1.400284e-05, 2.279945e-05, 1.218394e-05, 8.782249e-06, 1.591799e-05, 
    9.480282e-06, 5.026709e-06, 4.552455e-06, 3.565377e-06, 2.726267e-06, 
    1.745247e-06, 5.0515e-07, 3.18843e-07, 2.148452e-07, 2.60554e-08,
  1.475727e-05, 1.99706e-05, 9.587568e-06, 3.626408e-06, 1.825503e-06, 
    2.536648e-06, 4.931187e-06, 4.499249e-06, 3.080037e-06, 2.656844e-06, 
    1.408623e-06, 3.379045e-07, 3.383187e-07, 4.319981e-07, 4.886247e-07,
  1.02661e-05, 6.481072e-06, 7.314729e-06, 7.715804e-06, 4.447549e-06, 
    3.010789e-06, 2.596185e-06, 4.690359e-06, 9.778532e-06, 1.640989e-05, 
    2.182371e-05, 1.999979e-05, 1.276732e-05, 3.911226e-06, 1.735047e-06,
  1.203702e-05, 8.32177e-06, 1.079413e-05, 1.049386e-05, 6.387526e-06, 
    3.556489e-06, 1.439387e-06, 4.313099e-06, 1.002005e-05, 1.885415e-05, 
    2.634994e-05, 2.437782e-05, 1.538023e-05, 3.192836e-06, 1.548861e-06,
  1.712569e-05, 1.451124e-05, 1.673554e-05, 1.55166e-05, 8.164289e-06, 
    2.025733e-06, 1.11976e-06, 5.122464e-06, 1.078169e-05, 2.036364e-05, 
    2.916608e-05, 2.677645e-05, 1.787345e-05, 7.05408e-06, 2.687206e-06,
  2.906211e-05, 3.023279e-05, 2.21431e-05, 1.786725e-05, 6.653544e-06, 
    1.647868e-06, 2.60052e-06, 3.581652e-06, 9.76525e-06, 1.926818e-05, 
    2.412031e-05, 2.394354e-05, 1.603064e-05, 7.906152e-06, 2.618192e-06,
  4.599498e-05, 4.539936e-05, 3.648326e-05, 1.536203e-05, 1.853719e-06, 
    1.26651e-06, 4.652468e-06, 1.56686e-06, 4.368445e-06, 1.211893e-05, 
    1.519855e-05, 1.550053e-05, 1.105418e-05, 5.199694e-06, 1.991128e-06,
  6.184679e-05, 5.268906e-05, 2.20933e-05, 1.208598e-05, 1.421496e-06, 
    7.004965e-07, 4.486201e-06, 8.772382e-06, 1.08612e-05, 1.087341e-05, 
    9.592977e-06, 9.278818e-06, 6.524303e-06, 3.544512e-06, 4.08107e-07,
  7.456303e-05, 4.08968e-05, 2.301297e-05, 1.405381e-05, 8.979438e-06, 
    8.456907e-06, 5.286231e-06, 1.103277e-05, 1.224828e-05, 9.106844e-06, 
    8.801632e-06, 7.330701e-06, 3.176512e-06, 1.149125e-06, 1.029395e-07,
  5.088366e-05, 3.066545e-05, 2.286633e-05, 1.642029e-05, 1.710276e-05, 
    1.303432e-05, 7.478015e-06, 6.280446e-06, 7.005077e-06, 6.671843e-06, 
    5.950906e-06, 4.109958e-06, 1.502585e-06, 5.101936e-07, 3.757414e-08,
  2.932997e-05, 2.128541e-05, 2.021781e-05, 2.136692e-05, 1.659944e-05, 
    8.382111e-06, 5.255194e-06, 5.91722e-06, 5.453644e-06, 4.114646e-06, 
    3.513745e-06, 1.752811e-06, 7.16507e-07, 2.993449e-07, 2.100603e-08,
  1.555406e-05, 7.394597e-06, 7.806731e-06, 3.764953e-07, 1.024057e-07, 
    2.053942e-06, 3.130464e-06, 3.990162e-06, 3.494605e-06, 2.537706e-06, 
    1.815186e-06, 9.404219e-07, 5.935387e-07, 5.057615e-07, 1.302866e-07,
  7.500432e-06, 6.276397e-06, 9.686873e-06, 1.186457e-05, 1.621335e-05, 
    2.316682e-05, 2.54918e-05, 3.009324e-05, 3.071205e-05, 2.684601e-05, 
    2.264406e-05, 1.807772e-05, 1.512922e-05, 9.408494e-06, 7.041894e-06,
  2.029599e-06, 2.277784e-06, 4.419565e-06, 1.109387e-05, 1.910815e-05, 
    3.313061e-05, 3.479791e-05, 2.913418e-05, 2.396856e-05, 1.831239e-05, 
    1.363726e-05, 1.17603e-05, 1.164785e-05, 6.111868e-06, 7.885887e-06,
  2.882682e-06, 2.465515e-06, 6.392329e-06, 1.783007e-05, 3.221219e-05, 
    3.974924e-05, 3.027392e-05, 2.109661e-05, 1.327985e-05, 7.667522e-06, 
    5.886417e-06, 6.849648e-06, 1.316818e-05, 1.457786e-05, 1.484811e-05,
  1.25783e-05, 1.407898e-05, 1.650421e-05, 2.679464e-05, 3.436295e-05, 
    1.896481e-05, 1.207677e-05, 1.141167e-05, 5.786248e-06, 3.376701e-06, 
    3.246004e-06, 8.364134e-06, 1.796407e-05, 2.052852e-05, 1.596666e-05,
  1.910347e-05, 2.437037e-05, 2.798059e-05, 2.208933e-05, 1.550651e-05, 
    1.12715e-05, 5.963661e-06, 3.891077e-06, 1.721341e-06, 2.235362e-06, 
    4.491907e-06, 1.327103e-05, 2.162529e-05, 1.883666e-05, 1.624404e-05,
  2.662209e-05, 2.801894e-05, 2.386016e-05, 1.43765e-05, 1.137532e-05, 
    6.638287e-06, 6.226e-06, 5.163729e-06, 2.68192e-06, 3.914221e-06, 
    7.749346e-06, 1.633876e-05, 2.297385e-05, 2.238568e-05, 1.614264e-05,
  2.79868e-05, 2.824463e-05, 2.838491e-05, 2.374069e-05, 1.990947e-05, 
    1.397134e-05, 6.524056e-06, 5.485941e-06, 5.52637e-06, 7.298049e-06, 
    1.264435e-05, 1.876028e-05, 2.128714e-05, 2.054624e-05, 1.348991e-05,
  2.54805e-05, 2.846113e-05, 3.169584e-05, 2.104206e-05, 2.270032e-05, 
    1.623183e-05, 6.725594e-06, 5.435504e-06, 7.118705e-06, 1.000851e-05, 
    1.519139e-05, 1.748473e-05, 1.70643e-05, 1.373863e-05, 9.106657e-06,
  1.661746e-05, 2.298328e-05, 1.923476e-05, 1.634393e-05, 1.573469e-05, 
    1.044251e-05, 5.838257e-06, 8.045972e-06, 9.66631e-06, 1.08556e-05, 
    1.182265e-05, 1.23911e-05, 1.036308e-05, 7.420772e-06, 3.56383e-06,
  9.793564e-06, 8.977941e-06, 4.01507e-06, 2.199294e-06, 3.876281e-07, 
    4.261337e-06, 5.697485e-06, 6.894397e-06, 7.44917e-06, 7.440951e-06, 
    7.10952e-06, 6.583027e-06, 4.887634e-06, 2.814894e-06, 1.314346e-06,
  1.465965e-06, 6.21954e-07, 4.488605e-07, 1.069178e-06, 3.988895e-06, 
    3.216951e-06, 3.614449e-06, 2.982127e-06, 6.103458e-06, 7.964066e-06, 
    8.877403e-06, 1.128938e-05, 1.869366e-05, 2.509514e-05, 2.709818e-05,
  3.915974e-06, 5.423079e-07, 6.744094e-08, 5.318657e-06, 4.194224e-06, 
    1.833396e-06, 3.009242e-06, 2.194523e-06, 1.776645e-06, 4.314571e-06, 
    4.800116e-06, 8.828812e-06, 1.285068e-05, 1.876489e-05, 2.553723e-05,
  7.672255e-06, 8.889693e-07, 3.837896e-07, 2.599234e-06, 4.230523e-06, 
    1.996916e-06, 1.666152e-06, 7.054029e-06, 4.628785e-06, 1.629025e-06, 
    2.810186e-06, 5.835046e-06, 1.012714e-05, 1.810517e-05, 1.918484e-05,
  1.922769e-05, 1.895546e-05, 8.435586e-06, 4.433317e-06, 7.520426e-06, 
    7.195339e-06, 2.012606e-06, 1.852155e-06, 2.047414e-06, 1.383837e-06, 
    2.061012e-06, 4.420805e-06, 8.050122e-06, 1.456048e-05, 1.276262e-05,
  2.032015e-05, 1.459773e-05, 1.961146e-05, 1.158763e-05, 3.0559e-06, 
    1.037855e-05, 9.227243e-06, 1.687829e-06, 2.14584e-06, 2.784339e-06, 
    3.951252e-06, 3.972805e-06, 7.599303e-06, 9.828771e-06, 1.118859e-05,
  2.270099e-05, 1.60068e-05, 1.969465e-05, 1.791925e-05, 8.992979e-06, 
    8.115885e-06, 1.089874e-05, 1.143769e-05, 9.196466e-06, 7.01063e-06, 
    4.782364e-06, 4.499675e-06, 5.585126e-06, 6.244267e-06, 5.262765e-06,
  2.385942e-05, 1.801114e-05, 2.093212e-05, 1.966529e-05, 2.32998e-05, 
    1.509428e-05, 7.39292e-06, 8.526657e-06, 7.351793e-06, 5.66489e-06, 
    5.6875e-06, 6.262261e-06, 5.703084e-06, 5.861928e-06, 5.146781e-06,
  2.263777e-05, 1.941481e-05, 1.788681e-05, 1.791216e-05, 2.386957e-05, 
    1.626531e-05, 6.009393e-06, 5.62708e-06, 7.106192e-06, 7.624613e-06, 
    7.396301e-06, 7.571454e-06, 7.23396e-06, 9.764952e-06, 1.109576e-05,
  2.322378e-05, 1.85846e-05, 1.33608e-05, 7.698451e-06, 1.077314e-05, 
    7.651593e-06, 4.695394e-06, 5.340069e-06, 6.693395e-06, 7.437671e-06, 
    8.270659e-06, 1.041144e-05, 1.106889e-05, 1.059733e-05, 7.102509e-06,
  2.184197e-05, 1.218207e-05, 8.711478e-06, 2.514586e-06, 9.863611e-07, 
    1.471378e-06, 2.148703e-06, 2.588908e-06, 2.781677e-06, 3.609101e-06, 
    5.94764e-06, 8.659257e-06, 8.570541e-06, 6.2402e-06, 3.603171e-06,
  2.330482e-05, 7.670861e-06, 1.541746e-06, 6.880825e-07, 1.531325e-06, 
    2.524191e-06, 1.52616e-06, 1.401784e-06, 2.802648e-06, 3.430477e-06, 
    5.912229e-06, 9.117658e-06, 1.256891e-05, 1.139843e-05, 9.187956e-06,
  2.777975e-05, 8.493864e-06, 1.682397e-06, 1.788343e-07, 1.71558e-06, 
    7.085832e-07, 1.200717e-06, 1.199454e-06, 1.763713e-06, 2.736565e-06, 
    5.651933e-06, 8.248034e-06, 1.154465e-05, 1.000433e-05, 9.524196e-06,
  3.943063e-05, 1.532194e-05, 3.905258e-06, 2.836666e-07, 2.518962e-06, 
    4.798524e-07, 2.562938e-07, 5.586401e-06, 5.850955e-06, 5.211981e-06, 
    5.960464e-06, 7.868308e-06, 8.342846e-06, 8.592656e-06, 1.034784e-05,
  5.460326e-05, 3.471784e-05, 1.523437e-05, 1.181574e-06, 5.016772e-06, 
    2.568703e-06, 5.209785e-07, 2.386732e-06, 2.635081e-06, 5.269239e-06, 
    8.850811e-06, 8.653848e-06, 7.790601e-06, 7.220422e-06, 9.30483e-06,
  6.643739e-05, 4.894125e-05, 2.605669e-05, 7.2119e-06, 1.626073e-06, 
    4.280874e-06, 3.606587e-06, 6.233872e-07, 4.755762e-06, 7.303273e-06, 
    9.744679e-06, 9.053348e-06, 8.886236e-06, 5.464107e-06, 8.208337e-06,
  7.618195e-05, 6.569538e-05, 4.167958e-05, 9.576251e-06, 3.911701e-06, 
    4.599705e-06, 5.661767e-06, 4.467712e-06, 5.390471e-06, 9.695054e-06, 
    6.3471e-06, 6.869147e-06, 7.189444e-06, 3.853641e-06, 3.205971e-06,
  8.460083e-05, 8.360187e-05, 5.935109e-05, 1.60484e-05, 7.250846e-06, 
    6.065704e-06, 3.457653e-06, 2.43328e-06, 3.087699e-06, 3.913538e-06, 
    3.019168e-06, 3.904529e-06, 4.225626e-06, 2.759758e-06, 1.672761e-06,
  8.837183e-05, 9.56881e-05, 7.528481e-05, 3.114056e-05, 6.760357e-06, 
    5.914074e-06, 2.065501e-06, 1.597724e-06, 1.429879e-06, 1.26408e-06, 
    1.863349e-06, 1.957597e-06, 2.506782e-06, 2.375029e-06, 1.647495e-06,
  9.854021e-05, 0.0001034592, 9.047279e-05, 5.684164e-05, 7.260568e-06, 
    1.574511e-06, 1.776064e-06, 8.20609e-07, 7.000588e-07, 6.198237e-07, 
    9.389245e-07, 1.450374e-06, 1.669475e-06, 1.127634e-06, 5.565163e-07,
  0.0001002569, 0.0001031726, 8.961857e-05, 7.790478e-05, 2.472395e-05, 
    7.863225e-07, 3.751956e-07, 5.695377e-07, 4.113091e-07, 2.378432e-07, 
    4.913866e-07, 8.277875e-07, 9.324611e-07, 6.032565e-07, 3.010057e-07,
  8.346894e-05, 8.520084e-05, 4.378451e-05, 1.69686e-06, 7.531766e-07, 
    1.271977e-06, 1.197663e-06, 2.941062e-06, 6.552918e-06, 7.871186e-06, 
    7.843612e-06, 7.849076e-06, 6.99077e-06, 4.552373e-06, 2.422817e-06,
  8.342534e-05, 7.842143e-05, 3.653023e-05, 1.789353e-06, 7.080303e-07, 
    1.28401e-06, 1.136621e-06, 1.394136e-06, 3.212193e-06, 6.221606e-06, 
    6.919135e-06, 7.683828e-06, 7.31979e-06, 3.290456e-06, 1.201776e-06,
  7.617329e-05, 7.68613e-05, 3.959262e-05, 1.728615e-06, 6.233783e-07, 
    1.334967e-06, 7.065544e-07, 2.94286e-06, 7.724323e-06, 6.739822e-06, 
    4.917105e-06, 4.615119e-06, 3.130067e-06, 1.290331e-06, 1.185098e-06,
  6.216995e-05, 7.6207e-05, 5.206746e-05, 2.768907e-06, 1.81455e-06, 
    1.985059e-07, 1.022425e-06, 2.339721e-06, 3.137269e-06, 8.762342e-06, 
    5.831669e-06, 2.672703e-06, 2.311768e-06, 2.096993e-06, 4.076026e-06,
  4.584041e-05, 7.747547e-05, 7.415206e-05, 7.589092e-06, 3.019535e-06, 
    3.192879e-06, 4.958005e-07, 8.672862e-07, 4.262285e-06, 8.737335e-06, 
    7.856104e-06, 5.295424e-06, 7.920959e-06, 9.927136e-06, 1.378568e-05,
  3.295397e-05, 5.700791e-05, 8.271032e-05, 1.784947e-05, 4.789771e-06, 
    5.150137e-06, 4.551979e-06, 2.875574e-06, 2.767773e-06, 7.972891e-06, 
    5.019493e-06, 4.74468e-06, 8.663947e-06, 1.011144e-05, 1.109858e-05,
  2.549784e-05, 3.523669e-05, 7.207553e-05, 2.842172e-05, 8.114507e-06, 
    7.233625e-06, 4.477253e-06, 2.566751e-06, 1.890506e-06, 2.396163e-06, 
    2.342544e-06, 3.800514e-06, 6.932552e-06, 9.961757e-06, 1.272095e-05,
  2.122107e-05, 2.236886e-05, 5.391936e-05, 3.469976e-05, 1.215068e-05, 
    8.966001e-06, 4.071103e-06, 1.738159e-06, 7.747362e-07, 1.025233e-06, 
    1.783627e-06, 3.286376e-06, 6.120503e-06, 9.79573e-06, 1.394318e-05,
  2.122872e-05, 2.214413e-05, 3.817843e-05, 3.803272e-05, 8.776588e-06, 
    6.448665e-06, 3.084116e-06, 1.522437e-06, 7.618314e-07, 7.716606e-07, 
    1.530714e-06, 3.049075e-06, 5.607119e-06, 9.315502e-06, 1.510954e-05,
  1.896386e-05, 2.232265e-05, 2.774505e-05, 3.864215e-05, 6.677767e-06, 
    3.02125e-06, 1.086349e-06, 1.568551e-06, 1.117854e-06, 1.202373e-06, 
    1.907597e-06, 2.830702e-06, 4.441009e-06, 7.927294e-06, 1.408851e-05,
  1.037417e-05, 5.223651e-06, 1.089607e-06, 1.840369e-06, 1.871359e-06, 
    3.1431e-06, 3.306606e-06, 1.790352e-06, 1.655179e-06, 1.244997e-06, 
    1.637978e-06, 2.002346e-06, 2.057684e-06, 1.515947e-06, 1.329775e-06,
  4.966552e-06, 2.419493e-06, 9.848313e-07, 1.197218e-06, 1.810503e-06, 
    2.730501e-06, 3.155516e-06, 2.280835e-06, 1.340712e-06, 6.121189e-07, 
    7.562411e-07, 1.174018e-06, 1.358728e-06, 6.756191e-07, 6.077585e-07,
  9.869738e-06, 2.563723e-06, 1.752074e-06, 1.734649e-06, 6.261181e-07, 
    2.110878e-06, 2.951625e-06, 8.628619e-06, 9.479334e-06, 2.594601e-06, 
    9.041263e-07, 1.404319e-06, 6.910819e-07, 3.300496e-07, 5.741829e-07,
  1.836387e-05, 1.464449e-05, 1.084703e-05, 3.725003e-06, 6.697519e-06, 
    5.532411e-06, 4.401249e-06, 8.19414e-06, 8.960184e-06, 9.577771e-06, 
    7.197315e-06, 3.178608e-06, 2.018705e-06, 2.881469e-06, 1.943898e-06,
  2.335363e-05, 1.74718e-05, 1.432307e-05, 9.898404e-06, 6.59879e-06, 
    1.034265e-05, 5.831996e-06, 2.422272e-06, 6.431058e-06, 1.650575e-05, 
    1.673008e-05, 1.149776e-05, 8.559875e-06, 5.90938e-06, 5.006256e-06,
  2.587642e-05, 1.951905e-05, 1.601471e-05, 1.336233e-05, 8.883638e-06, 
    8.191531e-06, 1.200315e-05, 1.975838e-05, 2.924082e-05, 2.813866e-05, 
    2.016764e-05, 1.65841e-05, 1.408708e-05, 1.084733e-05, 8.287136e-06,
  2.806521e-05, 2.64901e-05, 2.181145e-05, 2.044863e-05, 1.516905e-05, 
    9.457375e-06, 1.001383e-05, 1.761366e-05, 2.451482e-05, 2.436516e-05, 
    2.316776e-05, 2.150528e-05, 1.801324e-05, 1.436975e-05, 1.06376e-05,
  3.415694e-05, 2.887066e-05, 1.878901e-05, 1.972972e-05, 1.689345e-05, 
    1.069989e-05, 9.166148e-06, 1.03574e-05, 1.464694e-05, 1.736564e-05, 
    2.208761e-05, 2.330075e-05, 2.118765e-05, 1.759571e-05, 1.335048e-05,
  3.657789e-05, 2.274739e-05, 2.299594e-05, 1.669717e-05, 1.436694e-05, 
    1.022549e-05, 7.240347e-06, 3.328927e-06, 6.573459e-06, 1.143655e-05, 
    1.784145e-05, 2.347145e-05, 2.259819e-05, 2.088569e-05, 1.839794e-05,
  2.549213e-05, 1.834999e-05, 1.372072e-05, 1.132664e-05, 9.381365e-06, 
    6.635712e-06, 9.179916e-07, 3.938805e-06, 3.641198e-06, 4.107123e-06, 
    1.030321e-05, 1.834849e-05, 2.320004e-05, 2.269155e-05, 2.296344e-05,
  3.031824e-06, 2.933662e-06, 5.595495e-06, 4.657883e-06, 6.380658e-07, 
    2.451401e-06, 1.764407e-06, 1.549201e-06, 1.189145e-06, 1.020952e-06, 
    6.553028e-07, 1.209138e-06, 2.293415e-06, 3.576677e-06, 1.212976e-05,
  5.19617e-07, 3.414178e-07, 3.718049e-06, 2.828177e-06, 1.379741e-06, 
    1.877263e-06, 2.315551e-06, 1.121912e-06, 1.134381e-06, 7.070686e-07, 
    5.315616e-07, 7.185871e-07, 1.598149e-06, 2.534093e-06, 7.964442e-06,
  8.513694e-06, 1.50441e-06, 1.321666e-06, 5.773779e-06, 2.790356e-06, 
    6.519353e-07, 1.427638e-06, 4.693366e-06, 5.122143e-06, 1.897854e-06, 
    9.723968e-07, 7.580389e-07, 9.246012e-07, 3.674612e-06, 6.890335e-06,
  2.354956e-05, 2.429684e-05, 1.231774e-05, 7.273635e-06, 8.68393e-06, 
    5.216858e-06, 2.542226e-06, 3.384e-06, 4.54139e-06, 3.237654e-06, 
    2.994757e-06, 1.637432e-06, 9.371807e-07, 2.955646e-06, 4.940441e-06,
  2.634454e-05, 2.731902e-05, 2.193062e-05, 1.036776e-05, 8.757954e-06, 
    8.9788e-06, 6.236626e-06, 1.576643e-06, 4.485081e-06, 3.656542e-06, 
    2.949774e-06, 1.822088e-06, 1.808173e-06, 1.693477e-06, 3.439902e-06,
  3.158868e-05, 2.081706e-05, 2.149045e-05, 1.829165e-05, 1.424295e-05, 
    8.105604e-06, 9.77303e-06, 1.095963e-05, 1.302269e-05, 9.554073e-06, 
    1.982322e-06, 6.990244e-07, 2.200479e-06, 1.337688e-06, 2.139734e-06,
  2.57734e-05, 3.086436e-05, 1.934433e-05, 2.308184e-05, 2.140263e-05, 
    9.95026e-06, 7.782482e-06, 1.04761e-05, 1.47868e-05, 1.094759e-05, 
    3.59576e-06, 1.753938e-06, 2.995803e-07, 2.984402e-07, 1.333208e-06,
  2.819819e-05, 1.91967e-05, 2.356379e-05, 1.724796e-05, 1.549885e-05, 
    1.134525e-05, 7.611474e-06, 5.204551e-06, 6.580946e-06, 1.017314e-05, 
    8.887755e-06, 3.374944e-06, 1.699321e-06, 1.49128e-06, 5.742854e-07,
  2.409309e-05, 1.893252e-05, 1.237677e-05, 1.022907e-05, 1.100531e-05, 
    9.130623e-06, 8.341334e-06, 4.155506e-06, 6.438552e-06, 1.118064e-05, 
    1.187264e-05, 9.324905e-06, 4.979966e-06, 2.779455e-06, 2.247607e-06,
  1.624958e-05, 1.251341e-05, 1.176749e-05, 6.665174e-06, 4.967611e-06, 
    5.519866e-06, 6.29837e-06, 7.938393e-06, 8.115549e-06, 7.680006e-06, 
    9.873776e-06, 1.232066e-05, 9.883292e-06, 6.932671e-06, 5.175779e-06,
  2.127666e-06, 1.491698e-06, 2.210309e-06, 2.843156e-06, 6.470639e-07, 
    9.822237e-07, 1.016336e-06, 1.757282e-06, 1.75382e-06, 1.382677e-06, 
    1.654525e-06, 1.67525e-06, 1.407593e-06, 7.831504e-07, 1.222631e-06,
  2.642817e-07, 2.761549e-07, 2.826359e-06, 2.979736e-06, 1.33406e-06, 
    8.772185e-07, 4.699261e-07, 8.060669e-07, 9.248104e-07, 1.886758e-06, 
    2.00992e-06, 1.734768e-06, 1.885357e-06, 1.218886e-06, 1.357243e-06,
  4.73204e-06, 8.657358e-07, 5.139525e-07, 3.677617e-06, 3.289098e-06, 
    1.44594e-06, 2.820031e-07, 1.39488e-06, 1.631928e-06, 6.523464e-07, 
    9.726308e-07, 1.670331e-06, 2.001053e-06, 2.386467e-06, 2.102225e-06,
  2.12238e-05, 1.67713e-05, 1.022043e-05, 1.742943e-06, 6.915172e-06, 
    2.788783e-06, 6.314569e-07, 1.110657e-06, 2.766114e-06, 2.522109e-06, 
    1.727508e-06, 2.080569e-06, 2.069154e-06, 3.433987e-06, 3.37548e-06,
  2.402893e-05, 2.163293e-05, 1.920456e-05, 6.801034e-06, 5.57798e-06, 
    6.638588e-06, 5.302069e-06, 5.452933e-07, 3.248362e-07, 2.980783e-06, 
    2.728302e-06, 1.268828e-06, 1.875953e-06, 3.0271e-06, 4.594582e-06,
  2.652872e-05, 2.33165e-05, 2.283241e-05, 1.591398e-05, 1.449091e-05, 
    8.025558e-06, 8.986673e-06, 6.084706e-06, 5.256754e-06, 5.92576e-06, 
    2.9678e-06, 2.102873e-06, 1.012753e-06, 3.13785e-06, 5.594371e-06,
  2.974565e-05, 3.02163e-05, 2.779469e-05, 2.72184e-05, 2.318653e-05, 
    9.192082e-06, 8.604084e-06, 7.365986e-06, 7.034303e-06, 5.747999e-06, 
    3.169106e-06, 2.034967e-06, 1.021119e-06, 1.557656e-06, 6.302173e-06,
  3.209148e-05, 3.002474e-05, 2.987702e-05, 1.652072e-05, 1.598648e-05, 
    8.869193e-06, 8.450893e-06, 8.149206e-06, 7.734687e-06, 6.052152e-06, 
    4.9507e-06, 2.234332e-06, 1.995417e-06, 2.478942e-06, 6.015149e-06,
  2.918527e-05, 1.956466e-05, 1.07687e-05, 8.26741e-06, 6.998775e-06, 
    4.829887e-06, 5.968186e-06, 9.448709e-06, 9.775013e-06, 8.909926e-06, 
    6.791229e-06, 3.836899e-06, 1.871363e-06, 2.005161e-06, 4.848538e-06,
  1.984759e-05, 1.009382e-05, 4.556801e-06, 3.176567e-06, 2.211771e-06, 
    2.806811e-06, 3.845162e-06, 9.283475e-06, 8.329998e-06, 7.369511e-06, 
    6.215758e-06, 5.852249e-06, 3.965003e-06, 2.454553e-06, 2.897894e-06,
  2.213573e-06, 2.067568e-06, 7.204149e-07, 7.515467e-07, 1.173558e-06, 
    9.697495e-07, 8.014809e-07, 6.343073e-07, 8.986715e-07, 1.980124e-06, 
    2.580897e-06, 2.951725e-06, 2.730782e-06, 2.23495e-06, 1.295311e-06,
  6.789421e-07, 1.329427e-07, 8.17214e-07, 5.32371e-07, 7.086199e-07, 
    5.220808e-07, 4.453571e-07, 7.62159e-07, 5.99008e-07, 1.599047e-06, 
    2.36845e-06, 3.546369e-06, 3.4845e-06, 3.116416e-06, 1.511272e-06,
  3.332791e-06, 1.626436e-07, 1.920225e-06, 9.924978e-07, 1.073941e-06, 
    7.729652e-07, 2.111399e-07, 4.21218e-07, 4.010832e-07, 4.722034e-07, 
    1.235279e-06, 2.494958e-06, 2.830952e-06, 2.768413e-06, 2.315957e-06,
  1.37533e-05, 1.118841e-05, 4.426928e-06, 1.472192e-06, 5.606419e-06, 
    1.63128e-06, 1.718231e-07, 1.969219e-07, 2.68458e-07, 5.878442e-07, 
    1.45589e-06, 2.093212e-06, 2.410064e-06, 3.249468e-06, 3.168449e-06,
  1.790215e-05, 1.811551e-05, 1.406684e-05, 3.597919e-06, 2.426129e-06, 
    3.823049e-06, 2.79311e-06, 4.384274e-07, 3.251406e-07, 1.802535e-06, 
    2.903221e-06, 2.076898e-06, 1.985946e-06, 2.429749e-06, 3.879693e-06,
  1.528511e-05, 1.714566e-05, 1.131189e-05, 8.431703e-06, 6.019888e-06, 
    4.07928e-06, 5.078743e-06, 4.129086e-06, 2.852899e-06, 2.631132e-06, 
    1.730742e-06, 1.348245e-06, 8.213319e-07, 3.404058e-06, 3.49776e-06,
  1.308645e-05, 1.797787e-05, 1.691305e-05, 1.673264e-05, 1.575873e-05, 
    3.96159e-06, 3.626669e-06, 3.798298e-06, 3.539248e-06, 2.144847e-06, 
    8.586729e-07, 7.002837e-07, 6.573763e-07, 1.93639e-06, 3.182102e-06,
  1.573968e-05, 1.744213e-05, 1.98479e-05, 1.58414e-05, 1.053238e-05, 
    3.313136e-06, 2.623521e-06, 2.710925e-06, 2.702079e-06, 2.049739e-06, 
    1.172872e-06, 8.330847e-07, 7.907828e-07, 1.900642e-06, 3.283298e-06,
  1.296856e-05, 1.427695e-05, 1.187815e-05, 6.565706e-06, 2.129818e-06, 
    2.312142e-06, 3.551499e-06, 3.738761e-06, 3.007281e-06, 2.431161e-06, 
    1.841431e-06, 1.444264e-06, 1.264558e-06, 2.276696e-06, 3.675862e-06,
  9.192044e-06, 4.430045e-06, 1.561775e-06, 2.0613e-06, 4.168063e-06, 
    5.483426e-06, 7.551071e-06, 1.148819e-05, 6.720082e-06, 2.517126e-06, 
    1.491383e-06, 1.547162e-06, 1.688042e-06, 2.483654e-06, 3.787181e-06,
  1.208575e-07, 4.032256e-07, 7.988679e-07, 7.013358e-07, 3.990068e-07, 
    6.522548e-07, 6.60233e-07, 6.213457e-07, 3.188078e-07, 7.275413e-07, 
    3.616136e-06, 9.714195e-06, 1.820508e-05, 2.371835e-05, 2.849306e-05,
  1.008418e-09, 1.172534e-07, 6.482917e-08, 4.239405e-08, 1.445942e-07, 
    4.539877e-07, 6.013208e-07, 7.883549e-07, 8.201721e-07, 7.01423e-07, 
    7.20745e-07, 1.607078e-06, 3.38047e-06, 6.528724e-06, 1.310444e-05,
  7.822359e-07, 2.028556e-08, 2.686908e-07, 3.338853e-07, 3.159661e-07, 
    1.602955e-06, 7.586546e-07, 5.285083e-07, 6.543796e-07, 3.439291e-07, 
    5.315486e-07, 1.314691e-06, 2.232676e-06, 2.08331e-06, 3.556703e-06,
  7.393344e-06, 3.963489e-06, 2.401912e-06, 2.614953e-06, 4.498228e-06, 
    6.488928e-06, 9.601748e-06, 6.521206e-06, 4.61145e-06, 5.51766e-06, 
    5.036363e-06, 2.174571e-06, 1.087148e-06, 9.844539e-07, 1.472091e-06,
  7.949875e-06, 8.473869e-06, 1.601866e-05, 5.116159e-06, 8.759104e-06, 
    1.681481e-05, 2.223554e-05, 2.111947e-05, 1.031482e-05, 8.357851e-06, 
    1.660607e-05, 1.134877e-05, 4.227488e-06, 2.689186e-06, 2.737804e-06,
  1.573487e-05, 1.877009e-05, 2.032089e-05, 9.8597e-06, 1.294573e-05, 
    2.060454e-05, 3.405183e-05, 3.814528e-05, 2.69999e-05, 1.977953e-05, 
    1.644714e-05, 1.188854e-05, 7.94899e-06, 7.221995e-06, 5.336737e-06,
  3.760064e-05, 4.836873e-05, 2.696183e-05, 1.507105e-05, 2.364936e-05, 
    2.169555e-05, 2.951597e-05, 3.147883e-05, 2.681516e-05, 1.881533e-05, 
    1.478008e-05, 1.203901e-05, 1.205224e-05, 1.166489e-05, 8.845827e-06,
  6.268493e-05, 4.086014e-05, 2.924143e-05, 2.845631e-05, 3.054038e-05, 
    2.655625e-05, 2.481787e-05, 2.2607e-05, 1.916257e-05, 1.638137e-05, 
    1.514842e-05, 1.395273e-05, 1.336436e-05, 1.217759e-05, 9.338996e-06,
  5.115058e-05, 3.200006e-05, 3.089594e-05, 2.783715e-05, 2.20804e-05, 
    2.242987e-05, 2.325457e-05, 2.084364e-05, 1.810271e-05, 1.438095e-05, 
    1.253625e-05, 1.144619e-05, 1.268719e-05, 1.139237e-05, 8.40762e-06,
  2.467376e-05, 1.522089e-05, 1.551134e-05, 2.060487e-05, 2.097989e-05, 
    1.629154e-05, 1.594637e-05, 2.182606e-05, 1.980596e-05, 1.347328e-05, 
    1.289846e-05, 1.218126e-05, 1.075808e-05, 1.037779e-05, 8.041709e-06,
  1.248813e-07, 6.986331e-07, 1.692257e-06, 1.856714e-06, 9.959947e-07, 
    1.812949e-06, 8.020675e-07, 3.15631e-07, 2.486522e-07, 2.19038e-07, 
    1.402101e-07, 1.694663e-07, 2.945862e-07, 4.498586e-07, 4.236643e-07,
  1.217088e-08, 3.572632e-08, 7.24375e-07, 2.108116e-06, 1.010094e-06, 
    2.688542e-06, 1.135773e-06, 1.654247e-06, 1.367513e-06, 1.000646e-06, 
    8.906674e-07, 7.19136e-07, 3.997027e-07, 6.179675e-07, 4.564822e-07,
  5.187848e-07, 9.933014e-08, 1.346566e-06, 6.27906e-06, 8.008457e-06, 
    1.548221e-05, 4.106656e-06, 8.898815e-06, 1.320396e-05, 1.079847e-05, 
    8.503763e-06, 8.469654e-06, 7.710201e-06, 4.752413e-06, 4.251252e-06,
  1.599092e-07, 3.643712e-06, 4.133853e-06, 1.047465e-05, 1.179667e-05, 
    1.013913e-05, 1.166701e-05, 3.800349e-06, 5.795989e-06, 1.710112e-05, 
    1.798751e-05, 1.303011e-05, 1.171578e-05, 1.177518e-05, 1.106349e-05,
  1.50438e-06, 6.541744e-06, 3.775845e-05, 1.3656e-05, 6.511764e-06, 
    8.112595e-06, 1.075828e-05, 1.178481e-05, 5.601099e-06, 6.88696e-06, 
    9.326823e-06, 7.877062e-06, 9.849963e-06, 1.145472e-05, 1.279621e-05,
  8.580659e-06, 4.491996e-05, 2.003376e-05, 9.868859e-06, 3.484829e-06, 
    9.302657e-06, 2.521649e-05, 2.222795e-05, 1.375169e-05, 7.003605e-06, 
    2.549688e-06, 2.969858e-06, 3.450701e-06, 6.062195e-06, 1.160766e-05,
  7.296288e-05, 3.776253e-05, 1.945438e-05, 1.089955e-05, 1.742854e-05, 
    2.070434e-05, 2.082797e-05, 1.047325e-05, 4.663524e-06, 2.073678e-06, 
    5.822682e-07, 3.403713e-07, 1.03722e-06, 1.627765e-06, 4.55058e-06,
  5.147436e-05, 2.927658e-05, 2.130247e-05, 2.180288e-05, 2.458381e-05, 
    1.291947e-05, 2.483252e-06, 1.389254e-06, 2.148701e-06, 1.059223e-06, 
    1.049898e-06, 1.050521e-06, 2.185791e-06, 2.923127e-06, 4.235852e-06,
  3.031698e-05, 2.585314e-05, 2.930941e-05, 2.015456e-05, 1.285967e-05, 
    3.325459e-06, 1.372301e-06, 2.821933e-06, 2.971228e-06, 7.793284e-06, 
    2.385233e-06, 2.557913e-06, 3.799994e-06, 4.813322e-06, 4.612807e-06,
  2.023492e-05, 1.486777e-05, 1.601154e-05, 1.351638e-05, 2.520957e-06, 
    1.47461e-06, 4.007647e-06, 8.057581e-06, 8.667391e-06, 4.417219e-06, 
    4.317028e-06, 3.600794e-06, 2.937313e-06, 3.52487e-06, 4.701229e-06,
  1.80594e-07, 2.053463e-08, 7.284962e-10, 4.767139e-09, 1.271713e-06, 
    2.539312e-06, 3.866496e-06, 1.496927e-06, 2.540087e-06, 3.001475e-06, 
    1.942126e-06, 1.512177e-06, 1.524177e-06, 1.021611e-06, 9.43807e-07,
  7.177132e-08, 8.087165e-09, 9.271001e-09, 1.958687e-07, 1.22026e-06, 
    5.311316e-06, 4.343138e-06, 7.183871e-07, 1.259661e-06, 3.147119e-06, 
    2.999526e-06, 2.955589e-06, 2.688704e-06, 2.565107e-06, 1.731896e-06,
  2.195624e-09, 3.776736e-10, 6.065251e-08, 3.340673e-06, 1.079772e-05, 
    1.829059e-05, 2.368498e-06, 2.452187e-06, 3.269849e-06, 4.479722e-06, 
    5.131011e-06, 4.133414e-06, 5.233893e-06, 4.422926e-06, 3.229686e-06,
  2.224176e-10, 4.058815e-08, 4.009165e-06, 2.514197e-05, 2.546623e-05, 
    5.360716e-06, 4.366052e-06, 2.111572e-06, 7.597134e-06, 1.263041e-05, 
    1.047231e-05, 8.043347e-06, 7.755868e-06, 6.98678e-06, 7.067491e-06,
  2.916179e-08, 3.06054e-06, 3.147623e-05, 3.76061e-05, 1.08273e-05, 
    1.386404e-06, 1.275843e-06, 3.332001e-06, 3.606139e-06, 1.089086e-05, 
    1.43848e-05, 1.056448e-05, 1.008902e-05, 9.828463e-06, 1.031196e-05,
  2.240929e-06, 3.250428e-05, 3.524979e-05, 1.044008e-05, 1.08546e-06, 
    2.867964e-07, 2.967988e-07, 1.781188e-06, 2.601633e-06, 2.396661e-06, 
    3.780905e-06, 5.51287e-06, 5.937238e-06, 6.988422e-06, 1.013903e-05,
  5.070297e-05, 3.409633e-05, 1.588854e-05, 6.08382e-06, 9.946469e-06, 
    1.033721e-06, 5.075067e-07, 7.183899e-07, 5.487612e-07, 5.8805e-07, 
    6.427246e-07, 9.961443e-07, 9.964291e-07, 1.176553e-06, 1.412371e-06,
  3.713957e-05, 1.522254e-05, 6.739696e-06, 7.936998e-06, 9.245709e-06, 
    1.639172e-06, 9.058567e-07, 9.174428e-07, 9.435637e-07, 7.468592e-07, 
    6.563514e-07, 1.688224e-06, 1.064976e-06, 8.488569e-07, 1.834775e-06,
  2.202958e-05, 4.749607e-06, 9.295182e-06, 8.023248e-06, 4.478879e-06, 
    2.510673e-06, 2.332137e-06, 3.122876e-06, 4.269317e-06, 4.026739e-06, 
    3.46501e-07, 2.640098e-07, 2.896388e-06, 2.000829e-06, 1.905298e-06,
  1.056164e-05, 3.300258e-06, 7.077395e-06, 2.58608e-06, 1.599519e-06, 
    3.376234e-06, 4.31516e-06, 1.176594e-05, 9.217517e-06, 1.908047e-06, 
    2.820715e-06, 4.198562e-07, 7.956857e-07, 3.433741e-06, 1.989288e-06,
  2.685793e-06, 1.782934e-06, 1.078179e-06, 6.899973e-07, 5.420082e-07, 
    5.610473e-07, 8.058383e-07, 1.262516e-06, 8.478331e-07, 4.407702e-07, 
    7.256671e-07, 4.991812e-07, 5.21202e-07, 5.71717e-07, 9.812269e-07,
  3.411124e-06, 2.515136e-06, 1.770924e-06, 1.361233e-06, 1.092209e-06, 
    1.865516e-06, 2.916063e-06, 1.966137e-06, 8.563865e-07, 9.515333e-07, 
    7.026792e-07, 1.677631e-07, 3.573781e-07, 1.767726e-06, 1.667915e-06,
  3.313019e-06, 3.458553e-06, 2.688375e-06, 2.397775e-06, 2.818067e-06, 
    8.825654e-06, 4.124186e-06, 5.498396e-06, 2.498391e-06, 8.409432e-07, 
    2.823847e-07, 2.297231e-07, 7.480983e-07, 8.776882e-07, 1.438055e-06,
  1.02271e-05, 5.855537e-06, 4.348386e-06, 4.612282e-06, 8.828351e-06, 
    8.601313e-06, 6.580472e-06, 3.114558e-06, 2.093347e-06, 6.829973e-07, 
    4.170571e-07, 7.542821e-07, 7.925127e-07, 9.28395e-07, 1.547487e-06,
  1.261516e-05, 1.089884e-05, 1.291016e-05, 7.624131e-06, 1.125504e-05, 
    7.960832e-06, 2.874835e-06, 5.708402e-06, 1.1887e-06, 6.8548e-08, 
    1.590269e-06, 1.064126e-06, 7.63423e-07, 1.40419e-06, 2.883637e-06,
  8.940412e-06, 1.006738e-05, 1.039383e-05, 1.066602e-05, 7.987232e-06, 
    5.183768e-06, 3.795188e-06, 2.118858e-06, 6.893283e-07, 8.769333e-07, 
    1.058742e-06, 1.463893e-06, 1.80645e-06, 1.798488e-06, 1.906361e-06,
  4.057249e-06, 1.437272e-05, 2.005262e-05, 1.357086e-05, 7.203781e-06, 
    3.144851e-06, 3.947948e-06, 2.846255e-06, 1.710971e-06, 1.347973e-06, 
    1.324574e-06, 2.554018e-06, 2.406281e-06, 2.1652e-06, 1.909075e-06,
  1.785454e-05, 1.978271e-05, 1.615496e-05, 7.606292e-06, 8.691098e-06, 
    6.630974e-06, 4.232588e-06, 1.807252e-06, 1.78078e-06, 1.536439e-06, 
    1.452721e-06, 2.655294e-06, 1.950684e-06, 1.533247e-06, 1.798178e-06,
  3.098622e-05, 1.986832e-05, 9.374673e-06, 1.446184e-05, 1.685255e-05, 
    8.859904e-06, 2.721404e-06, 1.929062e-06, 3.288076e-06, 2.062718e-06, 
    1.045978e-06, 1.026179e-06, 1.371295e-06, 1.888801e-06, 1.182879e-06,
  1.78484e-05, 1.95914e-05, 3.10087e-05, 3.282864e-05, 1.745862e-05, 
    4.266079e-06, 1.980388e-06, 5.861489e-06, 7.066651e-06, 1.78932e-06, 
    2.016384e-06, 3.802206e-07, 8.17496e-07, 1.578522e-06, 1.577511e-06,
  2.229675e-05, 1.806293e-05, 1.238953e-05, 6.271703e-06, 2.414155e-06, 
    1.215607e-06, 1.07038e-06, 1.070831e-06, 9.894637e-07, 1.023375e-06, 
    8.722344e-07, 1.203922e-06, 1.573736e-06, 1.937693e-06, 1.784025e-06,
  1.593504e-05, 1.700456e-05, 1.183503e-05, 6.989644e-06, 3.564628e-06, 
    1.964827e-06, 1.578303e-06, 1.618991e-06, 1.58744e-06, 1.903233e-06, 
    2.667989e-06, 2.890205e-06, 2.679538e-06, 3.329167e-06, 2.602107e-06,
  1.229424e-05, 1.404041e-05, 1.097461e-05, 6.601852e-06, 3.607694e-06, 
    4.043823e-06, 2.57701e-06, 2.768309e-06, 3.152019e-06, 2.873457e-06, 
    2.98838e-06, 3.498994e-06, 3.080626e-06, 3.06775e-06, 4.393512e-06,
  1.454092e-05, 1.557934e-05, 1.416321e-05, 7.648295e-06, 3.940404e-06, 
    3.176742e-06, 4.730146e-06, 3.845633e-06, 4.263049e-06, 4.211444e-06, 
    4.472868e-06, 4.094562e-06, 4.190538e-06, 5.311122e-06, 8.777375e-06,
  1.631286e-05, 1.554409e-05, 1.518412e-05, 1.009629e-05, 5.518741e-06, 
    4.44222e-06, 4.045267e-06, 5.116954e-06, 4.377687e-06, 3.86019e-06, 
    6.011271e-06, 5.442946e-06, 4.904917e-06, 7.779627e-06, 1.116968e-05,
  1.189253e-05, 1.726224e-05, 1.808169e-05, 1.101739e-05, 8.386477e-06, 
    5.500256e-06, 5.701416e-06, 6.010598e-06, 4.035692e-06, 6.808547e-06, 
    8.33687e-06, 6.133911e-06, 6.921141e-06, 9.720386e-06, 9.776637e-06,
  1.046815e-05, 1.610478e-05, 1.827963e-05, 1.440013e-05, 1.301857e-05, 
    6.243121e-06, 6.887706e-06, 1.25474e-05, 1.614517e-05, 1.296065e-05, 
    9.048308e-06, 8.558403e-06, 9.478555e-06, 7.499088e-06, 3.911407e-06,
  1.423629e-05, 1.59529e-05, 1.4574e-05, 1.444978e-05, 1.587191e-05, 
    7.178458e-06, 1.222021e-05, 1.81579e-05, 1.884957e-05, 1.622518e-05, 
    1.403671e-05, 1.13627e-05, 5.666949e-06, 2.358719e-06, 1.707372e-06,
  1.430404e-05, 1.765369e-05, 1.775783e-05, 1.362731e-05, 7.727194e-06, 
    1.729421e-05, 2.664163e-05, 2.827206e-05, 2.213174e-05, 1.44398e-05, 
    7.155728e-06, 2.706602e-06, 1.742475e-06, 1.05106e-06, 9.786324e-07,
  1.563852e-05, 2.78672e-05, 1.482931e-05, 1.749023e-05, 2.996789e-05, 
    3.873275e-05, 3.277592e-05, 1.837437e-05, 8.47854e-06, 2.089538e-06, 
    7.046715e-07, 6.89121e-07, 4.383204e-07, 1.254055e-06, 2.499214e-06,
  2.357137e-06, 6.770687e-06, 1.370914e-05, 1.506099e-05, 1.296124e-05, 
    8.541745e-06, 6.485814e-06, 5.455179e-06, 5.57744e-06, 7.547234e-06, 
    7.594253e-06, 5.960915e-06, 4.120192e-06, 3.366984e-06, 3.070883e-06,
  4.835043e-06, 9.88687e-06, 1.887682e-05, 2.458689e-05, 2.43693e-05, 
    1.597134e-05, 1.089123e-05, 1.069841e-05, 9.57825e-06, 9.929677e-06, 
    8.408115e-06, 7.088377e-06, 4.733559e-06, 3.640385e-06, 2.942863e-06,
  1.066835e-05, 8.026489e-06, 1.969154e-05, 3.043207e-05, 3.190414e-05, 
    2.066354e-05, 1.748518e-05, 2.054906e-05, 1.741733e-05, 1.137003e-05, 
    7.815408e-06, 7.122303e-06, 5.950579e-06, 4.365609e-06, 3.560063e-06,
  1.931941e-05, 1.432774e-05, 2.687361e-05, 3.280207e-05, 3.607689e-05, 
    2.777914e-05, 2.170529e-05, 2.081443e-05, 1.706914e-05, 1.321958e-05, 
    1.002122e-05, 8.190933e-06, 7.639231e-06, 6.779766e-06, 5.593988e-06,
  1.693828e-05, 1.380663e-05, 2.400543e-05, 3.744852e-05, 3.632809e-05, 
    3.144824e-05, 2.190977e-05, 9.262796e-06, 7.929289e-06, 1.090261e-05, 
    1.35968e-05, 1.004323e-05, 8.728556e-06, 7.288558e-06, 6.666672e-06,
  1.911411e-05, 1.592975e-05, 1.958639e-05, 3.68096e-05, 3.65427e-05, 
    2.368558e-05, 1.69529e-05, 1.098328e-05, 8.438401e-06, 8.302274e-06, 
    7.861698e-06, 7.053489e-06, 6.733959e-06, 6.53976e-06, 7.843531e-06,
  2.694474e-05, 2.310234e-05, 2.768668e-05, 3.771338e-05, 3.644886e-05, 
    1.850991e-05, 8.997544e-06, 7.106433e-06, 5.698098e-06, 4.241961e-06, 
    4.022028e-06, 4.367607e-06, 4.871067e-06, 6.193531e-06, 9.545039e-06,
  4.272882e-05, 3.513519e-05, 3.481135e-05, 3.698807e-05, 3.168832e-05, 
    1.637493e-05, 7.011251e-06, 5.007201e-06, 3.77187e-06, 4.068133e-06, 
    4.554726e-06, 7.649685e-06, 1.042263e-05, 9.823353e-06, 7.897075e-06,
  4.091962e-05, 4.613561e-05, 3.594806e-05, 2.629157e-05, 1.842831e-05, 
    1.398514e-05, 1.124266e-05, 1.043277e-05, 9.877552e-06, 8.944126e-06, 
    5.487955e-06, 2.916468e-06, 1.955952e-06, 8.250584e-07, 5.364593e-07,
  2.980238e-05, 1.842049e-05, 1.249301e-05, 7.852163e-06, 9.556576e-06, 
    9.546022e-06, 5.661635e-06, 5.988201e-06, 4.011185e-06, 8.52552e-07, 
    4.43657e-07, 3.815752e-07, 2.537111e-07, 2.168471e-07, 4.061581e-07,
  4.909546e-06, 3.405466e-06, 6.015767e-06, 8.085258e-06, 8.685886e-06, 
    9.358845e-06, 8.947199e-06, 9.63804e-06, 1.445951e-05, 1.523138e-05, 
    7.9204e-06, 9.325228e-06, 1.209241e-05, 1.264227e-05, 1.66668e-05,
  2.380655e-06, 3.104394e-06, 5.204581e-06, 6.503514e-06, 9.207677e-06, 
    7.787364e-06, 8.654167e-06, 1.247453e-05, 1.569669e-05, 1.879325e-05, 
    1.550862e-05, 1.513965e-05, 1.35654e-05, 1.262273e-05, 1.35675e-05,
  9.179865e-06, 4.660564e-06, 5.891153e-06, 6.675009e-06, 9.398344e-06, 
    1.423284e-05, 7.58787e-06, 1.493324e-05, 1.395308e-05, 1.431522e-05, 
    1.421766e-05, 1.414393e-05, 1.451593e-05, 1.470729e-05, 1.598787e-05,
  2.016406e-05, 2.620385e-05, 2.245969e-05, 1.377953e-05, 1.329553e-05, 
    1.348808e-05, 1.250149e-05, 1.586084e-05, 1.556388e-05, 1.257019e-05, 
    1.229451e-05, 1.317211e-05, 1.423787e-05, 1.742431e-05, 1.666613e-05,
  2.934751e-05, 3.030226e-05, 3.026717e-05, 2.112452e-05, 1.472341e-05, 
    1.397412e-05, 1.09987e-05, 9.497604e-06, 9.903657e-06, 1.565081e-05, 
    1.690704e-05, 1.450632e-05, 1.499709e-05, 1.747352e-05, 1.827471e-05,
  3.515164e-05, 3.081218e-05, 2.85897e-05, 2.203028e-05, 1.357792e-05, 
    1.121986e-05, 1.175549e-05, 1.634201e-05, 2.465887e-05, 2.72171e-05, 
    2.526472e-05, 2.553394e-05, 2.464514e-05, 2.42728e-05, 2.552467e-05,
  3.461646e-05, 3.463996e-05, 3.246075e-05, 2.528125e-05, 1.483736e-05, 
    7.166952e-06, 6.97308e-06, 1.155051e-05, 1.882808e-05, 2.215541e-05, 
    2.526158e-05, 2.80041e-05, 2.667534e-05, 2.511445e-05, 2.501554e-05,
  3.051609e-05, 3.091655e-05, 2.685323e-05, 2.154522e-05, 1.481579e-05, 
    5.774513e-06, 4.531724e-06, 4.274327e-06, 5.097461e-06, 7.861648e-06, 
    1.061615e-05, 1.251236e-05, 1.230348e-05, 1.116292e-05, 1.051271e-05,
  3.174938e-05, 2.451474e-05, 1.765125e-05, 8.807538e-06, 3.215458e-06, 
    1.916248e-06, 2.410724e-06, 2.403719e-06, 2.077795e-06, 9.681193e-07, 
    4.131875e-07, 3.570376e-07, 4.725566e-07, 3.665193e-07, 3.696804e-07,
  2.688095e-05, 2.120903e-05, 1.416987e-05, 3.944517e-06, 1.418146e-06, 
    1.36502e-06, 1.287233e-06, 2.22265e-06, 1.750496e-06, 3.242727e-07, 
    4.325672e-07, 4.526933e-07, 3.60305e-07, 2.323158e-07, 2.141756e-07,
  3.998788e-07, 6.963038e-08, 3.674177e-08, 7.157196e-08, 4.111437e-07, 
    1.791936e-06, 4.139951e-06, 3.452632e-06, 4.090749e-06, 9.055969e-06, 
    9.816889e-06, 1.329898e-05, 1.777081e-05, 1.977997e-05, 1.711927e-05,
  9.722713e-08, 1.821511e-08, 7.167203e-09, 2.234615e-07, 1.993144e-07, 
    5.916309e-07, 1.316063e-06, 1.675597e-06, 8.682349e-07, 2.979599e-06, 
    8.977568e-06, 1.508627e-05, 1.906269e-05, 1.896363e-05, 1.432491e-05,
  6.114923e-06, 1.836594e-07, 1.005445e-07, 6.059562e-07, 7.142229e-07, 
    5.10889e-06, 1.484119e-06, 1.962736e-06, 3.465372e-06, 4.066663e-06, 
    6.659467e-06, 1.0625e-05, 1.328531e-05, 1.585407e-05, 1.839682e-05,
  1.459387e-05, 1.282071e-05, 1.021314e-05, 3.222748e-06, 3.795857e-06, 
    5.530244e-06, 4.571159e-06, 7.343016e-07, 1.820295e-06, 5.026159e-06, 
    4.634129e-06, 5.917308e-06, 7.830048e-06, 1.227274e-05, 1.60426e-05,
  1.752058e-05, 1.32018e-05, 1.569916e-05, 8.468629e-06, 1.298882e-05, 
    1.157688e-05, 7.281296e-06, 1.599018e-06, 3.484447e-06, 4.400486e-06, 
    4.839403e-06, 4.535521e-06, 5.033768e-06, 5.849617e-06, 8.930686e-06,
  2.543651e-05, 1.094763e-05, 1.285109e-05, 2.312789e-05, 2.763908e-05, 
    2.11858e-05, 7.515304e-06, 3.346433e-06, 4.466824e-06, 5.241063e-06, 
    3.899541e-06, 5.153176e-06, 7.060192e-06, 8.93894e-06, 1.092814e-05,
  4.561491e-05, 3.148537e-05, 3.468828e-05, 5.678512e-05, 5.499419e-05, 
    1.088827e-05, 2.169524e-06, 2.352457e-06, 2.571505e-06, 2.325852e-06, 
    2.514665e-06, 3.240747e-06, 4.603381e-06, 7.19585e-06, 1.133592e-05,
  5.905917e-05, 5.666031e-05, 7.610414e-05, 7.586123e-05, 1.467651e-05, 
    1.475074e-06, 7.118794e-07, 1.280352e-06, 1.743521e-06, 2.211792e-06, 
    2.095132e-06, 1.358917e-06, 1.19686e-06, 2.145927e-06, 4.392459e-06,
  5.352266e-05, 5.870904e-05, 6.717681e-05, 2.595508e-05, 2.798153e-06, 
    7.971179e-07, 1.185024e-06, 1.456019e-06, 2.444524e-06, 3.407905e-06, 
    2.549235e-06, 1.081782e-06, 3.476506e-07, 4.107979e-07, 6.976858e-07,
  4.646806e-05, 4.094244e-05, 3.413262e-05, 1.002089e-05, 7.991576e-07, 
    1.056546e-06, 1.642215e-06, 3.710451e-06, 3.53861e-06, 2.593778e-06, 
    2.390609e-06, 1.435535e-06, 5.153219e-07, 2.551616e-07, 2.958951e-07,
  4.115419e-06, 4.509863e-06, 5.264014e-06, 5.220728e-06, 4.370555e-06, 
    3.741314e-06, 4.624622e-06, 5.649318e-06, 5.107532e-06, 4.649345e-06, 
    3.665195e-06, 2.497364e-06, 2.286863e-06, 2.294823e-06, 4.340702e-06,
  1.779456e-06, 2.074192e-06, 2.971874e-06, 4.15516e-06, 3.461752e-06, 
    2.542168e-06, 3.589937e-06, 4.109815e-06, 4.082977e-06, 2.974092e-06, 
    2.968075e-06, 4.538788e-06, 5.462869e-06, 6.976812e-06, 7.425596e-06,
  9.410035e-07, 3.365367e-06, 2.053925e-06, 2.723077e-06, 9.002674e-07, 
    2.091205e-06, 1.628823e-06, 3.662745e-06, 3.114402e-06, 3.74337e-06, 
    5.782893e-06, 9.8747e-06, 1.369723e-05, 1.595266e-05, 1.631466e-05,
  4.985486e-06, 6.191286e-06, 5.860712e-06, 4.477513e-06, 6.626279e-07, 
    4.197716e-07, 5.465154e-06, 8.646e-06, 1.277626e-05, 1.720442e-05, 
    1.581655e-05, 1.260884e-05, 1.139258e-05, 1.108014e-05, 1.048636e-05,
  1.689815e-05, 1.693712e-05, 1.956372e-05, 5.099536e-06, 3.755324e-06, 
    8.820569e-06, 1.58333e-05, 2.923606e-05, 1.734128e-05, 1.243366e-05, 
    9.956118e-06, 5.895695e-06, 4.377902e-06, 4.007692e-06, 4.497198e-06,
  3.335627e-05, 3.202609e-05, 3.536393e-05, 2.90359e-05, 2.905321e-05, 
    3.839867e-05, 3.528488e-05, 1.291379e-05, 3.982007e-06, 2.198185e-06, 
    1.692195e-06, 2.212261e-06, 2.609171e-06, 2.868915e-06, 2.497096e-06,
  5.323295e-05, 4.951038e-05, 3.673269e-05, 3.272396e-05, 2.269534e-05, 
    1.293157e-05, 3.7264e-06, 2.217595e-06, 1.251857e-06, 1.283711e-06, 
    2.253322e-06, 2.652329e-06, 2.07234e-06, 2.14846e-06, 2.045121e-06,
  4.054676e-05, 3.503322e-05, 2.178072e-05, 9.740887e-06, 3.900291e-06, 
    1.539585e-06, 9.043328e-07, 4.236316e-07, 1.045431e-06, 1.413401e-06, 
    1.536086e-06, 1.379464e-06, 8.331945e-07, 1.07897e-06, 1.35625e-06,
  2.156424e-05, 2.009707e-05, 9.755225e-06, 6.817098e-06, 2.721866e-06, 
    1.024218e-06, 5.31224e-07, 5.287101e-07, 1.027831e-06, 9.018125e-07, 
    9.735803e-07, 1.466101e-06, 2.482745e-06, 2.850761e-06, 2.17753e-06,
  1.087821e-05, 8.922071e-06, 7.001562e-06, 1.6411e-06, 7.212939e-07, 
    5.097515e-07, 4.171369e-07, 1.525672e-06, 1.761364e-06, 1.292811e-06, 
    2.694502e-06, 4.727234e-06, 6.446136e-06, 5.088122e-06, 2.702967e-06,
  1.382932e-05, 2.62202e-05, 8.028926e-05, 0.0001393281, 0.0001429296, 
    0.0001290288, 0.0001057481, 7.795159e-05, 5.522622e-05, 4.731688e-05, 
    4.716304e-05, 4.923122e-05, 5.002783e-05, 4.408939e-05, 3.861147e-05,
  9.162965e-06, 1.124388e-05, 3.320499e-05, 0.0001045496, 0.0001427837, 
    0.0001336592, 0.0001171391, 8.987501e-05, 6.469672e-05, 5.146631e-05, 
    4.928187e-05, 5.14723e-05, 4.563592e-05, 4.023583e-05, 4.01132e-05,
  6.69046e-06, 4.52662e-06, 7.513324e-06, 2.211895e-05, 5.766088e-05, 
    9.645944e-05, 0.0001038359, 0.0001065164, 9.5966e-05, 7.804141e-05, 
    6.135907e-05, 5.086347e-05, 4.161417e-05, 3.185804e-05, 2.687448e-05,
  2.123619e-05, 1.495856e-05, 1.026701e-05, 4.30716e-06, 1.027787e-05, 
    2.891645e-05, 5.757955e-05, 6.262466e-05, 6.803749e-05, 6.847796e-05, 
    5.319432e-05, 3.927577e-05, 2.853585e-05, 1.957708e-05, 1.097696e-05,
  2.800252e-05, 2.124255e-05, 1.791507e-05, 2.855123e-06, 1.83136e-06, 
    6.509983e-06, 9.803878e-06, 1.843315e-05, 3.432885e-05, 3.256711e-05, 
    2.38208e-05, 1.663034e-05, 9.516535e-06, 4.738639e-06, 2.519299e-06,
  2.598838e-05, 2.255016e-05, 1.320579e-05, 3.813932e-06, 1.681987e-06, 
    2.653044e-06, 3.070676e-06, 4.636831e-06, 6.297482e-06, 5.770738e-06, 
    4.215714e-06, 2.479135e-06, 1.305673e-06, 5.92279e-07, 3.506735e-07,
  1.718816e-05, 9.16703e-06, 3.897636e-06, 1.276852e-08, 3.400267e-09, 
    2.225003e-07, 4.341221e-07, 2.029621e-06, 1.346267e-06, 9.380963e-07, 
    7.134956e-07, 4.75037e-07, 2.782302e-07, 1.407254e-07, 9.236664e-08,
  1.071745e-05, 1.247921e-05, 8.366643e-06, 3.850108e-06, 1.759572e-07, 
    8.101851e-08, 4.000256e-08, 6.097103e-08, 3.486591e-07, 3.660222e-07, 
    1.73065e-07, 2.330981e-07, 4.898197e-07, 9.50513e-07, 2.157175e-06,
  1.153235e-05, 9.988294e-06, 9.647932e-06, 6.287079e-06, 1.955942e-07, 
    6.950057e-08, 2.010743e-07, 4.93089e-07, 4.949882e-07, 5.585829e-07, 
    4.415905e-07, 4.723441e-07, 2.200445e-06, 6.007785e-06, 9.146805e-06,
  2.194183e-05, 1.5827e-05, 1.398104e-05, 3.401965e-06, 4.207266e-07, 
    5.498288e-08, 2.150613e-07, 8.987222e-07, 3.290286e-07, 6.604113e-07, 
    1.217465e-06, 1.942988e-06, 5.841284e-06, 1.151689e-05, 1.581442e-05,
  1.27105e-06, 6.418084e-06, 4.543457e-05, 9.93421e-05, 8.997634e-05, 
    6.460482e-05, 4.522901e-05, 2.847009e-05, 1.961976e-05, 9.082013e-06, 
    3.958487e-06, 4.069648e-06, 2.314717e-06, 5.998032e-06, 5.260761e-06,
  9.539234e-07, 1.528715e-06, 1.621191e-05, 8.46378e-05, 0.0001126973, 
    9.356533e-05, 7.920782e-05, 3.483188e-05, 1.806266e-05, 8.057896e-06, 
    2.619543e-06, 2.585358e-06, 1.202804e-06, 4.911942e-06, 3.23577e-06,
  6.658607e-06, 1.770935e-06, 4.092759e-06, 4.512348e-05, 0.0001046662, 
    0.0001017736, 8.26652e-05, 6.217987e-05, 2.190505e-05, 8.427603e-06, 
    3.487214e-06, 2.424922e-06, 2.326795e-06, 4.104957e-06, 6.88745e-06,
  9.169349e-06, 3.772298e-06, 2.476328e-06, 1.325308e-05, 7.146217e-05, 
    9.567245e-05, 8.426827e-05, 6.622593e-05, 4.025456e-05, 1.88659e-05, 
    1.274446e-05, 9.335682e-06, 1.170693e-05, 1.558151e-05, 1.930249e-05,
  9.803961e-06, 2.456559e-06, 3.738681e-07, 2.951748e-06, 2.647152e-05, 
    9.520617e-05, 8.060009e-05, 5.876657e-05, 7.822653e-05, 4.892761e-05, 
    3.440371e-05, 2.615372e-05, 2.616225e-05, 2.560151e-05, 2.813205e-05,
  3.909835e-06, 8.191795e-07, 2.884808e-09, 4.03501e-07, 4.182345e-06, 
    3.316128e-05, 0.0001071334, 9.217676e-05, 6.053752e-05, 4.83284e-05, 
    3.544313e-05, 2.956725e-05, 2.683557e-05, 2.471603e-05, 2.590719e-05,
  1.741254e-06, 5.193853e-07, 2.222914e-09, 8.366613e-08, 1.020116e-06, 
    3.777513e-06, 2.988616e-05, 7.797305e-05, 6.398784e-05, 3.50898e-05, 
    2.735727e-05, 2.632581e-05, 2.502395e-05, 2.257059e-05, 2.11457e-05,
  1.123855e-06, 1.52073e-06, 6.360384e-07, 5.596669e-07, 8.311298e-07, 
    4.394382e-07, 2.921525e-06, 1.637577e-05, 2.913807e-05, 3.182172e-05, 
    3.230324e-05, 3.074719e-05, 2.816907e-05, 2.726118e-05, 2.581952e-05,
  2.097509e-05, 1.695331e-05, 1.418526e-05, 1.135159e-05, 5.228318e-06, 
    8.849697e-07, 4.091885e-07, 2.094044e-06, 1.147909e-05, 2.019986e-05, 
    2.509717e-05, 2.817512e-05, 3.106585e-05, 3.463577e-05, 3.101984e-05,
  8.424965e-05, 9.195059e-05, 6.750884e-05, 4.836814e-05, 3.534351e-05, 
    1.494673e-05, 1.236816e-06, 1.849693e-07, 1.066521e-06, 5.516538e-06, 
    1.200099e-05, 2.2991e-05, 2.90035e-05, 3.017067e-05, 2.168488e-05,
  3.642578e-08, 5.593555e-09, 2.206906e-08, 2.239176e-06, 1.079628e-05, 
    2.581876e-05, 1.688167e-05, 3.123885e-06, 3.690692e-07, 3.541106e-06, 
    4.448807e-06, 4.836881e-06, 6.018652e-06, 1.021168e-05, 1.214272e-05,
  1.576469e-06, 1.563465e-07, 1.334255e-07, 4.902794e-06, 1.272386e-05, 
    2.229711e-05, 1.765728e-05, 5.156907e-06, 3.945821e-06, 3.615541e-06, 
    2.885761e-06, 3.649986e-06, 8.62764e-06, 1.62642e-05, 1.224378e-05,
  9.672151e-06, 3.191669e-06, 6.009247e-07, 6.632486e-06, 1.923448e-05, 
    2.748349e-05, 2.291134e-05, 1.696496e-05, 1.21012e-05, 6.053163e-06, 
    2.669027e-06, 6.081967e-06, 1.325308e-05, 1.600583e-05, 1.112037e-05,
  2.035674e-05, 1.27442e-05, 6.523913e-06, 5.500369e-06, 2.155213e-05, 
    3.032636e-05, 2.704067e-05, 2.346879e-05, 1.567385e-05, 8.154543e-06, 
    7.233792e-06, 1.321387e-05, 1.719178e-05, 1.267106e-05, 9.842167e-06,
  2.797102e-05, 2.177122e-05, 1.157515e-05, 3.3051e-06, 1.52937e-05, 
    3.54704e-05, 2.169382e-05, 2.738391e-05, 2.603352e-05, 8.507252e-06, 
    1.63359e-05, 2.212358e-05, 1.339393e-05, 7.230904e-06, 6.868157e-06,
  2.487049e-05, 2.374646e-05, 1.141959e-05, 2.822598e-06, 6.237781e-06, 
    2.002859e-05, 3.356009e-05, 9.175748e-06, 4.057615e-06, 7.936133e-06, 
    1.868164e-05, 1.615506e-05, 8.796331e-06, 5.612947e-06, 7.30815e-06,
  2.929017e-05, 2.394767e-05, 1.71588e-05, 4.264676e-06, 2.05871e-06, 
    9.905368e-06, 2.145599e-05, 1.607743e-05, 5.774696e-06, 8.744107e-06, 
    1.688987e-05, 1.141123e-05, 7.750362e-06, 6.710735e-06, 5.619077e-06,
  4.313924e-05, 3.035152e-05, 1.999962e-05, 9.383009e-06, 1.079418e-06, 
    4.647899e-06, 1.336936e-05, 2.046905e-05, 9.417749e-06, 8.883308e-06, 
    1.256715e-05, 1.026764e-05, 7.068888e-06, 6.47792e-06, 6.409043e-06,
  5.26428e-05, 3.810195e-05, 2.585025e-05, 1.443809e-05, 4.000138e-06, 
    2.14208e-06, 7.262773e-06, 1.268062e-05, 1.760943e-05, 1.037576e-05, 
    9.256534e-06, 8.796308e-06, 7.085468e-06, 9.493761e-06, 1.114797e-05,
  2.089038e-05, 2.081962e-05, 3.243902e-05, 2.66497e-05, 1.322971e-05, 
    5.491115e-06, 4.80583e-06, 6.843585e-06, 9.554927e-06, 1.034041e-05, 
    9.256945e-06, 9.017022e-06, 1.012425e-05, 1.659999e-05, 1.7259e-05,
  8.481023e-06, 6.53405e-06, 5.400012e-06, 7.007673e-06, 4.656521e-06, 
    2.01286e-06, 3.636959e-06, 3.722636e-06, 2.864392e-06, 5.077317e-06, 
    3.951695e-06, 3.776035e-06, 4.277756e-06, 4.780653e-06, 7.457878e-06,
  1.013628e-05, 9.264144e-06, 8.082746e-06, 7.761374e-06, 6.675528e-06, 
    3.878734e-06, 3.505148e-06, 3.397304e-06, 3.927722e-06, 1.479694e-06, 
    5.75172e-06, 5.597981e-06, 6.040478e-06, 6.242711e-06, 7.095908e-06,
  1.893335e-05, 1.309389e-05, 1.341858e-05, 1.198077e-05, 9.415575e-06, 
    9.447467e-06, 4.875717e-06, 3.385524e-06, 3.46035e-06, 3.995917e-06, 
    5.951469e-06, 5.195654e-06, 6.15457e-06, 5.419266e-06, 7.476406e-06,
  2.331684e-05, 3.800853e-05, 4.324695e-05, 1.575238e-05, 1.291972e-05, 
    1.368389e-05, 1.172765e-05, 5.943537e-06, 3.459609e-06, 7.962256e-06, 
    4.900692e-06, 6.288496e-06, 7.871667e-06, 6.723245e-06, 6.04847e-06,
  2.967002e-05, 3.017539e-05, 4.040391e-05, 1.511947e-05, 1.113899e-05, 
    1.123224e-05, 1.427566e-05, 1.764728e-05, 6.470272e-06, 3.354538e-06, 
    7.903473e-06, 9.856101e-06, 5.48155e-06, 4.346108e-06, 6.12227e-06,
  3.751572e-05, 3.572556e-05, 3.689205e-05, 1.3198e-05, 6.760674e-06, 
    3.060755e-06, 1.012052e-05, 5.972306e-06, 2.960349e-06, 6.008652e-06, 
    4.430103e-06, 5.27165e-06, 5.905492e-06, 8.341573e-06, 1.829272e-05,
  4.305034e-05, 4.725371e-05, 4.470745e-05, 2.509654e-05, 1.36527e-05, 
    3.307246e-06, 8.20689e-06, 3.146501e-06, 4.916117e-06, 9.283932e-06, 
    4.237649e-06, 5.103183e-06, 8.552883e-06, 1.65871e-05, 2.148382e-05,
  4.983707e-05, 5.708155e-05, 4.891448e-05, 3.134017e-05, 1.989397e-05, 
    4.721412e-06, 6.198904e-06, 6.116865e-06, 7.261492e-06, 1.148576e-05, 
    4.482326e-06, 5.697063e-06, 1.34636e-05, 1.799986e-05, 4.663428e-06,
  4.510094e-05, 4.597657e-05, 2.312474e-05, 2.219962e-05, 1.57358e-05, 
    6.86397e-06, 6.507978e-06, 7.596538e-06, 1.428982e-05, 1.207051e-05, 
    5.400243e-06, 9.764682e-06, 1.498271e-05, 5.202085e-06, 1.255411e-07,
  2.986728e-05, 1.103538e-05, 1.030925e-05, 1.193648e-05, 1.369841e-05, 
    1.085532e-05, 8.580066e-06, 8.937765e-06, 1.64112e-05, 1.041705e-05, 
    8.126878e-06, 1.224948e-05, 6.971083e-06, 6.116763e-07, 8.282745e-09,
  6.607635e-06, 2.125458e-07, 2.785012e-08, 7.492371e-08, 4.398102e-06, 
    2.066878e-05, 1.282213e-05, 5.245375e-06, 7.872985e-06, 7.268103e-06, 
    7.635869e-06, 5.66121e-06, 1.058756e-05, 2.362747e-05, 3.812885e-05,
  1.90378e-06, 3.708344e-07, 1.04083e-07, 3.391265e-07, 1.909752e-06, 
    1.373915e-05, 1.134152e-05, 4.403176e-06, 3.818216e-06, 4.122018e-06, 
    6.108969e-06, 7.867166e-06, 6.391823e-06, 1.126034e-05, 2.330612e-05,
  1.889085e-05, 3.994734e-06, 2.192639e-06, 1.180042e-06, 1.184242e-06, 
    1.557324e-05, 7.648276e-06, 6.401814e-06, 2.028099e-06, 3.113584e-06, 
    8.206164e-06, 1.004037e-05, 8.613671e-06, 9.121035e-06, 1.143439e-05,
  2.434197e-05, 2.999737e-05, 2.294804e-05, 2.148646e-06, 1.60997e-06, 
    7.410611e-06, 1.219802e-05, 5.060331e-06, 2.637071e-06, 6.730004e-06, 
    8.58821e-06, 1.118646e-05, 1.055054e-05, 1.2076e-05, 1.096156e-05,
  2.587703e-05, 3.021942e-05, 3.187018e-05, 2.859549e-06, 1.594139e-06, 
    2.406332e-06, 8.714184e-06, 3.446839e-06, 1.699565e-05, 8.363882e-06, 
    9.987151e-06, 1.383155e-05, 1.084549e-05, 7.119776e-06, 7.983376e-06,
  3.125373e-05, 3.334905e-05, 3.285695e-05, 9.025805e-06, 2.372536e-06, 
    2.422983e-06, 4.973431e-06, 5.214021e-06, 2.976991e-06, 1.179669e-05, 
    8.523619e-06, 1.05623e-05, 1.030235e-05, 4.359851e-06, 3.034301e-06,
  2.725951e-05, 4.327426e-05, 4.492772e-05, 1.350278e-05, 3.154659e-06, 
    2.265656e-06, 2.026268e-06, 2.471129e-06, 2.328946e-06, 4.54286e-06, 
    9.010092e-06, 1.038079e-05, 7.873236e-06, 2.130791e-06, 3.477297e-07,
  1.771883e-05, 2.341048e-05, 2.06271e-05, 1.472146e-05, 5.924024e-06, 
    3.005916e-06, 1.571931e-06, 1.99982e-06, 1.58743e-06, 4.259709e-06, 
    6.42828e-06, 6.715696e-06, 3.376934e-06, 2.406562e-07, 6.35125e-08,
  8.103398e-06, 1.308263e-05, 1.154724e-05, 1.414536e-05, 9.459099e-06, 
    4.535834e-06, 2.292271e-06, 2.808212e-06, 4.400434e-06, 4.75193e-06, 
    4.885818e-06, 3.100638e-06, 3.353226e-07, 1.185335e-07, 1.183013e-07,
  3.864111e-06, 3.660641e-06, 4.450253e-06, 4.324278e-06, 4.596581e-06, 
    5.834619e-06, 4.925723e-06, 3.659024e-06, 4.849994e-06, 4.143268e-06, 
    3.032139e-06, 3.781487e-07, 1.690023e-07, 1.938869e-07, 2.811093e-08,
  2.857191e-06, 5.346594e-07, 1.018487e-06, 3.544548e-06, 3.12978e-06, 
    4.81503e-06, 2.807589e-06, 7.934032e-06, 4.042604e-06, 4.73671e-06, 
    4.413885e-06, 7.094928e-06, 1.284469e-05, 1.618195e-05, 2.085001e-05,
  9.88438e-07, 4.376413e-07, 7.632441e-07, 2.576837e-06, 1.473213e-06, 
    1.277459e-06, 1.165012e-06, 5.494247e-06, 2.31569e-06, 3.299954e-06, 
    3.065879e-06, 7.529067e-06, 1.269657e-05, 1.160607e-05, 1.981632e-05,
  7.517819e-06, 2.262272e-06, 3.633168e-06, 4.092271e-06, 1.360018e-06, 
    4.11438e-06, 7.791501e-07, 6.342854e-06, 5.29449e-06, 3.549571e-06, 
    3.108519e-06, 3.975685e-06, 5.920167e-06, 1.093358e-05, 2.057857e-05,
  6.336073e-06, 1.269551e-05, 1.519842e-05, 6.266868e-06, 3.913744e-06, 
    1.283425e-06, 1.569684e-06, 1.237406e-06, 1.226707e-06, 4.308298e-06, 
    1.580506e-06, 1.403533e-06, 1.284495e-06, 1.874241e-06, 4.085938e-06,
  7.653063e-06, 1.011568e-05, 1.365362e-05, 2.694714e-06, 3.143737e-06, 
    3.32889e-06, 2.485794e-07, 7.563926e-07, 4.831329e-06, 3.421967e-06, 
    1.493111e-06, 6.539587e-07, 2.414693e-07, 2.475111e-07, 4.331943e-07,
  6.284085e-06, 8.299573e-06, 1.107776e-05, 5.578059e-06, 3.240955e-06, 
    2.519808e-06, 3.444077e-06, 2.977996e-06, 2.083112e-06, 2.298547e-06, 
    1.278447e-06, 4.85706e-07, 5.277755e-07, 3.209139e-07, 4.682665e-07,
  5.667449e-06, 9.084449e-06, 1.113338e-05, 1.023215e-05, 4.777486e-06, 
    3.118325e-06, 1.304222e-06, 9.321028e-07, 1.306599e-06, 2.005176e-06, 
    7.785719e-07, 7.175892e-07, 5.512348e-07, 4.537835e-07, 4.422032e-07,
  4.472454e-06, 6.322271e-06, 1.14048e-05, 1.159712e-05, 1.071348e-05, 
    7.451675e-06, 3.450014e-06, 1.143211e-06, 6.235186e-07, 4.78601e-07, 
    5.927112e-07, 5.075577e-07, 4.805089e-07, 4.390865e-07, 4.3637e-07,
  1.630206e-06, 3.181437e-06, 6.266865e-06, 1.486956e-05, 1.863558e-05, 
    1.418427e-05, 1.010827e-05, 4.587484e-06, 9.418278e-07, 2.991382e-07, 
    2.34524e-07, 3.202003e-07, 3.589327e-07, 3.916416e-07, 5.183081e-07,
  6.41131e-07, 1.683331e-06, 6.492434e-06, 2.12884e-05, 3.302706e-05, 
    2.687819e-05, 1.629229e-05, 1.139107e-05, 4.484291e-06, 9.588658e-07, 
    3.746926e-07, 3.49707e-07, 3.265016e-07, 1.595646e-07, 5.14249e-07,
  1.47573e-06, 4.681267e-06, 1.096231e-05, 1.867182e-05, 2.005293e-05, 
    2.12676e-05, 2.307491e-05, 1.911818e-05, 1.607486e-05, 1.444973e-05, 
    8.315509e-06, 6.12312e-06, 6.3127e-06, 7.124946e-06, 1.162888e-05,
  2.324768e-06, 5.893228e-06, 9.977083e-06, 1.795271e-05, 1.989312e-05, 
    1.618533e-05, 1.820699e-05, 2.225043e-05, 1.833913e-05, 1.678139e-05, 
    1.318427e-05, 6.906214e-06, 3.855583e-06, 5.020598e-06, 5.64721e-06,
  2.961664e-06, 4.809544e-06, 8.928617e-06, 1.824091e-05, 2.773656e-05, 
    2.330862e-05, 9.512338e-06, 1.372136e-05, 2.082867e-05, 2.164031e-05, 
    1.712713e-05, 1.144661e-05, 4.140995e-06, 7.719232e-07, 1.304104e-06,
  4.829899e-06, 6.863836e-06, 1.299045e-05, 2.016821e-05, 3.093778e-05, 
    3.403832e-05, 2.499657e-05, 9.493758e-06, 1.23764e-05, 1.914739e-05, 
    2.207797e-05, 1.517006e-05, 7.069396e-06, 1.623893e-06, 1.405448e-07,
  4.950021e-06, 8.538244e-06, 1.319024e-05, 2.05941e-05, 3.252845e-05, 
    3.424469e-05, 3.582356e-05, 2.98941e-05, 1.405257e-05, 1.020829e-05, 
    2.216998e-05, 1.734244e-05, 9.578234e-06, 1.949431e-06, 4.327527e-07,
  1.036081e-05, 9.171087e-06, 1.179108e-05, 1.898813e-05, 3.115443e-05, 
    3.548579e-05, 4.542008e-05, 4.144385e-05, 2.589331e-05, 2.081293e-05, 
    1.893556e-05, 1.516937e-05, 1.15919e-05, 3.001192e-06, 1.034431e-06,
  1.029333e-05, 1.029146e-05, 1.026155e-05, 1.598244e-05, 3.049712e-05, 
    3.306435e-05, 4.00658e-05, 4.503851e-05, 3.962109e-05, 2.78166e-05, 
    1.909394e-05, 1.582813e-05, 1.293234e-05, 3.302793e-06, 1.595655e-06,
  1.086769e-05, 7.851952e-06, 7.468249e-06, 1.392239e-05, 3.282418e-05, 
    3.330136e-05, 3.895648e-05, 4.494853e-05, 3.96005e-05, 3.265101e-05, 
    2.580519e-05, 1.954489e-05, 1.265498e-05, 2.905529e-06, 1.296804e-06,
  7.232183e-06, 4.765081e-06, 5.13095e-06, 1.060454e-05, 2.717554e-05, 
    2.785868e-05, 3.011778e-05, 3.958883e-05, 4.081932e-05, 3.512866e-05, 
    2.844026e-05, 2.151632e-05, 1.057615e-05, 2.788373e-06, 1.391776e-06,
  4.65598e-06, 2.958412e-06, 1.869267e-06, 3.818021e-06, 8.458086e-06, 
    1.030271e-05, 1.555328e-05, 2.550311e-05, 3.388518e-05, 3.088626e-05, 
    2.844049e-05, 2.07881e-05, 9.294458e-06, 3.4123e-06, 1.841372e-06,
  9.733226e-06, 1.875568e-05, 2.651564e-05, 2.304172e-05, 1.272898e-05, 
    9.729786e-06, 9.520051e-06, 7.494637e-06, 7.103237e-06, 1.037166e-05, 
    1.898014e-05, 2.832575e-05, 3.325667e-05, 3.550378e-05, 3.058705e-05,
  7.763367e-06, 1.213667e-05, 1.662779e-05, 1.153484e-05, 5.994943e-06, 
    3.006253e-06, 4.228052e-06, 6.557891e-06, 3.647682e-06, 4.179559e-06, 
    8.185476e-06, 2.009327e-05, 3.054514e-05, 2.855056e-05, 2.503689e-05,
  7.515002e-06, 1.28927e-05, 1.14329e-05, 7.15745e-06, 3.609601e-06, 
    6.09406e-06, 1.681594e-06, 4.555905e-06, 5.776456e-06, 3.290057e-06, 
    4.625274e-06, 1.239697e-05, 2.416136e-05, 2.497244e-05, 2.340945e-05,
  7.804935e-06, 1.288256e-05, 1.581812e-05, 8.004167e-06, 3.433952e-06, 
    5.514425e-06, 8.027847e-06, 2.483973e-06, 2.76999e-06, 3.255914e-06, 
    3.303554e-06, 8.285539e-06, 1.769989e-05, 2.529624e-05, 2.410843e-05,
  6.310185e-06, 9.406443e-06, 9.276744e-06, 3.511243e-06, 3.896857e-06, 
    6.158067e-06, 8.561957e-06, 1.516191e-05, 2.861026e-05, 8.464671e-06, 
    4.195615e-06, 6.184771e-06, 1.717815e-05, 2.349467e-05, 1.832574e-05,
  4.235699e-06, 5.524889e-06, 6.871463e-06, 4.358541e-06, 7.908058e-06, 
    1.264859e-05, 9.754162e-06, 1.193614e-05, 1.890591e-05, 1.093329e-05, 
    7.395244e-06, 5.494631e-06, 1.724666e-05, 1.391357e-05, 6.551376e-06,
  5.68476e-06, 3.668855e-06, 6.026113e-06, 9.007333e-06, 9.011469e-06, 
    7.040855e-06, 9.246983e-06, 9.58131e-06, 8.591444e-06, 6.703292e-06, 
    4.7662e-06, 4.726931e-06, 9.971376e-06, 6.376828e-06, 1.776155e-06,
  3.432311e-06, 2.191285e-06, 7.256084e-06, 7.374222e-06, 8.216655e-06, 
    4.075862e-06, 3.641343e-06, 5.203771e-06, 6.831413e-06, 7.614181e-06, 
    1.262799e-06, 4.38916e-06, 4.447214e-06, 2.453785e-06, 1.305363e-06,
  2.62367e-06, 2.521291e-06, 3.868792e-06, 4.745079e-06, 7.172675e-06, 
    3.788321e-06, 2.045917e-06, 1.754687e-06, 4.381861e-06, 4.971848e-06, 
    4.031809e-06, 3.25722e-06, 2.191298e-06, 1.574767e-06, 5.740289e-07,
  3.140642e-06, 2.410171e-06, 2.835434e-06, 4.17163e-06, 5.493984e-06, 
    6.114498e-06, 3.638081e-06, 2.885893e-06, 3.424661e-06, 3.027928e-06, 
    3.590222e-06, 2.712324e-06, 1.343521e-06, 1.057863e-06, 7.29107e-07,
  6.031657e-07, 1.94382e-06, 3.410537e-06, 4.938014e-06, 5.027573e-06, 
    5.831987e-06, 4.758986e-06, 2.792258e-06, 4.627833e-06, 5.826408e-06, 
    3.46825e-06, 4.841118e-06, 3.235692e-06, 5.692445e-07, 3.738388e-06,
  5.795418e-07, 1.629186e-06, 3.52746e-06, 5.99646e-06, 9.114502e-06, 
    9.48582e-06, 9.81892e-06, 7.166051e-06, 7.011585e-06, 4.677683e-06, 
    1.511134e-06, 3.331346e-06, 1.243811e-06, 2.872758e-06, 3.267209e-07,
  9.452701e-07, 2.546745e-06, 4.160592e-06, 6.845165e-06, 1.462973e-05, 
    2.779147e-05, 9.089025e-06, 1.166943e-05, 1.222739e-05, 7.492119e-06, 
    3.872279e-06, 2.206101e-06, 2.138923e-06, 5.066991e-06, 1.570892e-06,
  2.129821e-06, 5.353869e-06, 6.735141e-06, 9.347216e-06, 1.728749e-05, 
    2.363886e-05, 2.898831e-05, 1.047337e-05, 1.259775e-05, 1.164794e-05, 
    8.356772e-06, 3.753139e-06, 4.394614e-06, 3.573502e-06, 4.118218e-06,
  3.623582e-06, 5.799456e-06, 8.645906e-06, 1.21087e-05, 1.838479e-05, 
    2.239284e-05, 2.676448e-05, 3.112967e-05, 1.996907e-05, 1.212694e-05, 
    1.40082e-05, 6.826506e-06, 4.064396e-06, 2.444458e-06, 5.434849e-06,
  6.456984e-06, 9.351489e-06, 1.261726e-05, 1.383309e-05, 1.789056e-05, 
    2.250986e-05, 3.320343e-05, 2.49549e-05, 2.007926e-05, 2.543923e-05, 
    2.014254e-05, 1.082849e-05, 5.305354e-06, 2.66434e-06, 2.830016e-06,
  7.804975e-06, 8.765212e-06, 1.31097e-05, 1.553636e-05, 2.051566e-05, 
    2.574728e-05, 3.293706e-05, 3.804691e-05, 3.631381e-05, 3.400521e-05, 
    3.049661e-05, 1.93004e-05, 8.791612e-06, 3.469265e-06, 1.369635e-06,
  7.71608e-06, 7.050313e-06, 1.086156e-05, 1.428533e-05, 1.800622e-05, 
    2.426667e-05, 3.35074e-05, 3.668338e-05, 3.93657e-05, 4.757883e-05, 
    4.763911e-05, 2.974239e-05, 1.325197e-05, 4.295082e-06, 1.245787e-06,
  9.319819e-06, 1.00787e-05, 1.29644e-05, 1.550233e-05, 1.671849e-05, 
    2.183804e-05, 3.235508e-05, 4.351713e-05, 5.341333e-05, 5.798023e-05, 
    5.21623e-05, 3.524373e-05, 1.556818e-05, 4.215314e-06, 1.078931e-06,
  1.008973e-05, 1.493605e-05, 1.685692e-05, 1.725286e-05, 1.690627e-05, 
    1.81432e-05, 2.709248e-05, 4.661396e-05, 6.857825e-05, 7.167758e-05, 
    5.696597e-05, 3.455849e-05, 1.19796e-05, 2.402789e-06, 1.132654e-06,
  6.638101e-06, 1.301942e-05, 1.782543e-05, 2.534626e-05, 2.907985e-05, 
    3.178216e-05, 3.381485e-05, 3.40043e-05, 3.841773e-05, 3.806161e-05, 
    2.752172e-05, 2.280989e-05, 1.840255e-05, 7.980732e-06, 2.107726e-06,
  6.158331e-06, 9.597584e-06, 1.545364e-05, 2.167601e-05, 2.038195e-05, 
    1.895581e-05, 2.530723e-05, 2.447783e-05, 2.11715e-05, 2.53448e-05, 
    3.069444e-05, 3.189598e-05, 2.547427e-05, 1.704046e-05, 9.442443e-06,
  5.017254e-06, 8.856165e-06, 1.329597e-05, 1.968556e-05, 2.390478e-05, 
    3.343881e-05, 1.409842e-05, 2.202973e-05, 2.487752e-05, 2.165356e-05, 
    2.435174e-05, 2.882192e-05, 3.017202e-05, 2.44482e-05, 2.298088e-05,
  5.98784e-06, 9.637763e-06, 1.741905e-05, 1.720458e-05, 2.334792e-05, 
    2.606469e-05, 3.442667e-05, 9.60217e-06, 1.584214e-05, 2.589181e-05, 
    2.743678e-05, 2.668694e-05, 3.397054e-05, 3.953476e-05, 3.369067e-05,
  5.072397e-06, 5.444701e-06, 1.310047e-05, 1.128843e-05, 1.354665e-05, 
    1.884197e-05, 2.447491e-05, 4.525565e-05, 3.229326e-05, 1.54449e-05, 
    2.218269e-05, 2.665855e-05, 3.638975e-05, 4.991259e-05, 4.753424e-05,
  5.772853e-06, 5.985385e-06, 1.033504e-05, 8.9901e-06, 8.447533e-06, 
    1.106621e-05, 1.649515e-05, 2.615687e-05, 2.328879e-05, 2.098322e-05, 
    2.40832e-05, 3.449217e-05, 5.279537e-05, 6.314324e-05, 5.560234e-05,
  7.536327e-06, 9.849145e-06, 7.960937e-06, 8.109299e-06, 6.285924e-06, 
    5.2246e-06, 6.717226e-06, 1.129161e-05, 1.338691e-05, 1.873858e-05, 
    2.850707e-05, 4.820794e-05, 6.713028e-05, 7.130772e-05, 4.782142e-05,
  1.143997e-05, 1.257395e-05, 9.801111e-06, 8.646679e-06, 6.033489e-06, 
    7.181767e-06, 4.738357e-06, 5.243964e-06, 6.67086e-06, 1.598077e-05, 
    3.030236e-05, 5.653385e-05, 8.246356e-05, 6.431402e-05, 2.46858e-05,
  1.568762e-05, 2.093203e-05, 1.19412e-05, 6.450409e-06, 4.943589e-06, 
    3.751538e-06, 3.309372e-06, 2.665819e-06, 5.97453e-06, 1.256368e-05, 
    2.302296e-05, 5.474315e-05, 5.482605e-05, 2.258072e-05, 3.99523e-06,
  1.615375e-05, 2.131334e-05, 1.489193e-05, 6.682694e-06, 4.159382e-06, 
    3.944489e-06, 3.437529e-06, 2.347167e-06, 4.853558e-06, 1.155209e-05, 
    1.946909e-05, 2.767286e-05, 1.818673e-05, 2.763691e-06, 4.463305e-07,
  4.101512e-05, 3.133074e-05, 2.57897e-05, 1.857648e-05, 9.792497e-06, 
    4.089478e-06, 3.961394e-06, 1.963772e-06, 6.483915e-06, 1.018852e-05, 
    1.775774e-05, 3.282847e-05, 3.984452e-05, 2.646388e-05, 1.063493e-05,
  4.14328e-05, 2.873408e-05, 2.162288e-05, 1.692032e-05, 1.024103e-05, 
    3.806688e-06, 2.175893e-06, 9.934391e-07, 1.750088e-06, 3.924121e-06, 
    9.03964e-06, 2.035352e-05, 2.824403e-05, 2.290268e-05, 2.156869e-05,
  3.803498e-05, 3.216425e-05, 2.395353e-05, 1.707575e-05, 1.112399e-05, 
    7.389408e-06, 1.732106e-06, 1.260554e-06, 3.015616e-06, 5.387753e-06, 
    7.448266e-06, 1.120346e-05, 1.593324e-05, 2.278015e-05, 3.73276e-05,
  3.938888e-05, 3.486237e-05, 2.75401e-05, 2.239769e-05, 1.197531e-05, 
    4.690702e-06, 3.687309e-06, 4.944704e-07, 5.355678e-07, 2.80055e-06, 
    4.339315e-06, 5.797706e-06, 1.162503e-05, 1.856421e-05, 3.396555e-05,
  4.30659e-05, 3.924857e-05, 3.195913e-05, 2.603415e-05, 1.750872e-05, 
    6.323052e-06, 3.976286e-06, 3.716373e-06, 6.83831e-06, 2.884454e-06, 
    5.072425e-06, 6.368673e-06, 6.990531e-06, 1.10531e-05, 3.025123e-05,
  4.477098e-05, 4.128373e-05, 3.466855e-05, 3.092836e-05, 2.254233e-05, 
    9.554949e-06, 9.21378e-06, 3.886159e-06, 3.719564e-06, 3.547747e-06, 
    3.352349e-06, 5.740018e-06, 7.484824e-06, 1.35696e-05, 3.697495e-05,
  3.856458e-05, 4.085762e-05, 3.604017e-05, 3.031586e-05, 2.750986e-05, 
    1.406261e-05, 8.285342e-06, 5.242468e-06, 1.917005e-06, 9.820038e-07, 
    3.329853e-06, 5.168516e-06, 1.064854e-05, 2.363082e-05, 3.947963e-05,
  3.346894e-05, 4.297211e-05, 3.737487e-05, 2.776522e-05, 2.617969e-05, 
    1.721402e-05, 8.585906e-06, 5.213619e-06, 2.027785e-06, 1.252404e-06, 
    2.887381e-06, 1.354412e-06, 3.892639e-06, 9.236095e-06, 1.191479e-05,
  2.917784e-05, 3.858234e-05, 3.012253e-05, 2.325791e-05, 2.1916e-05, 
    1.889723e-05, 1.216116e-05, 6.770893e-06, 4.00053e-06, 2.555603e-06, 
    1.662173e-06, 1.523119e-06, 1.367869e-06, 1.157944e-06, 1.861623e-06,
  2.025328e-05, 2.366154e-05, 2.109369e-05, 2.015796e-05, 1.74276e-05, 
    1.704446e-05, 1.408262e-05, 9.34011e-06, 8.745174e-06, 1.104247e-05, 
    8.11157e-06, 3.61347e-06, 1.644223e-06, 1.041105e-06, 6.044559e-07,
  3.889613e-05, 4.117163e-05, 4.374503e-05, 3.295602e-05, 1.796316e-05, 
    8.894998e-06, 4.047855e-06, 4.508968e-06, 2.520714e-06, 3.133598e-06, 
    5.248157e-06, 4.943696e-06, 3.532622e-06, 6.722124e-06, 1.425048e-05,
  3.598855e-05, 3.733556e-05, 4.268298e-05, 3.206674e-05, 1.660696e-05, 
    5.61484e-06, 4.23752e-06, 3.602456e-06, 1.177572e-06, 3.418594e-07, 
    1.108947e-06, 3.577455e-06, 5.80003e-06, 6.092935e-06, 7.500123e-06,
  2.591107e-05, 3.39742e-05, 3.995591e-05, 3.338035e-05, 2.344384e-05, 
    1.678593e-05, 3.896346e-06, 5.369693e-06, 2.418677e-06, 7.122343e-07, 
    1.172658e-06, 2.306061e-06, 3.439695e-06, 3.581982e-06, 3.295255e-06,
  2.303939e-05, 2.741561e-05, 3.64737e-05, 3.621188e-05, 2.147714e-05, 
    1.876957e-05, 2.200099e-05, 3.607297e-06, 3.594878e-06, 1.795983e-06, 
    1.472443e-06, 1.384547e-06, 2.727595e-06, 3.715613e-06, 3.154121e-06,
  1.460509e-05, 2.108531e-05, 3.129655e-05, 3.04531e-05, 1.947203e-05, 
    1.428495e-05, 2.022769e-05, 2.776962e-05, 7.999642e-06, 1.798253e-06, 
    2.061307e-06, 1.857879e-06, 3.446252e-06, 5.965988e-06, 6.494792e-06,
  1.006728e-05, 1.258265e-05, 2.490653e-05, 2.407088e-05, 1.525813e-05, 
    1.068547e-05, 1.273063e-05, 1.194606e-05, 6.227807e-06, 6.395406e-06, 
    5.623945e-06, 4.213111e-06, 4.251625e-06, 4.853247e-06, 5.560096e-06,
  7.860331e-06, 1.352633e-05, 2.021242e-05, 1.922524e-05, 1.450123e-05, 
    9.149779e-06, 7.660852e-06, 9.469903e-06, 8.367711e-06, 5.869184e-06, 
    7.839971e-06, 9.727079e-06, 7.599115e-06, 7.589967e-06, 3.810824e-06,
  1.200404e-05, 1.341312e-05, 1.631941e-05, 1.468135e-05, 1.159511e-05, 
    8.448323e-06, 8.014434e-06, 7.353605e-06, 7.203326e-06, 9.405928e-06, 
    1.287964e-05, 1.288467e-05, 1.227618e-05, 1.078916e-05, 8.249416e-06,
  1.055901e-05, 1.295019e-05, 1.46495e-05, 8.415638e-06, 6.028593e-06, 
    6.719053e-06, 8.023253e-06, 7.712202e-06, 5.832712e-06, 9.469477e-06, 
    1.601327e-05, 1.90663e-05, 1.684608e-05, 1.286778e-05, 1.007646e-05,
  3.715172e-06, 9.530222e-06, 1.100721e-05, 6.094502e-06, 4.448116e-06, 
    5.125815e-06, 4.408828e-06, 5.145233e-06, 4.792059e-06, 7.750371e-06, 
    1.920909e-05, 2.666587e-05, 2.475762e-05, 1.927682e-05, 1.416791e-05,
  1.439743e-05, 1.192392e-05, 1.245272e-05, 9.383219e-06, 3.219293e-06, 
    4.963544e-06, 6.567281e-06, 6.815436e-06, 1.556924e-05, 1.71741e-05, 
    8.469676e-06, 3.56599e-06, 5.689407e-06, 4.914103e-06, 5.438765e-06,
  1.019714e-05, 1.05648e-05, 1.179964e-05, 7.093552e-06, 1.537817e-06, 
    2.009106e-06, 6.853895e-06, 7.140505e-06, 1.135985e-05, 1.909482e-05, 
    2.007678e-05, 1.17695e-05, 5.602792e-06, 6.108985e-06, 4.572797e-06,
  9.197968e-06, 1.050248e-05, 1.017436e-05, 5.201524e-06, 2.462209e-06, 
    8.972913e-06, 3.371903e-06, 1.009156e-05, 1.45952e-05, 2.250028e-05, 
    2.582111e-05, 2.325742e-05, 1.432057e-05, 6.51588e-06, 4.255116e-06,
  1.102068e-05, 1.261986e-05, 1.40299e-05, 7.50139e-06, 3.516194e-06, 
    7.932478e-06, 8.234923e-06, 3.980907e-06, 7.364662e-06, 1.412486e-05, 
    1.918843e-05, 2.466567e-05, 2.628754e-05, 1.815756e-05, 9.966549e-06,
  1.183686e-05, 1.099616e-05, 1.211055e-05, 7.232907e-06, 4.052902e-06, 
    4.564081e-06, 5.427207e-06, 9.233634e-06, 1.271872e-05, 9.297801e-06, 
    1.403614e-05, 1.957972e-05, 2.795052e-05, 2.849449e-05, 2.24433e-05,
  1.161815e-05, 1.016236e-05, 1.052998e-05, 8.818809e-06, 6.866701e-06, 
    3.930336e-06, 4.154159e-06, 9.433869e-06, 1.220731e-05, 9.187334e-06, 
    8.967043e-06, 1.198132e-05, 1.713449e-05, 2.53968e-05, 2.971306e-05,
  1.64255e-05, 1.471155e-05, 9.100119e-06, 8.152577e-06, 6.290172e-06, 
    4.756052e-06, 4.342132e-06, 2.696957e-06, 3.256094e-06, 3.327058e-06, 
    4.064829e-06, 5.303519e-06, 8.289448e-06, 1.503204e-05, 2.376429e-05,
  1.847534e-05, 1.780826e-05, 1.051144e-05, 6.323956e-06, 3.919811e-06, 
    3.470754e-06, 2.769641e-06, 3.105492e-06, 3.135676e-06, 2.599355e-06, 
    2.823292e-06, 3.322484e-06, 4.056401e-06, 6.919201e-06, 1.488002e-05,
  2.089241e-05, 1.916016e-05, 7.797305e-06, 3.713711e-06, 1.398799e-06, 
    3.352866e-06, 2.999853e-06, 1.828931e-06, 1.780411e-06, 2.347998e-06, 
    3.041642e-06, 2.834437e-06, 3.425802e-06, 5.319316e-06, 1.049865e-05,
  1.96816e-05, 1.166406e-05, 4.822872e-06, 2.600563e-06, 2.331818e-06, 
    2.684914e-06, 1.80937e-06, 4.229384e-06, 3.939029e-06, 1.533045e-06, 
    1.775857e-06, 1.92466e-06, 2.155235e-06, 3.326262e-06, 8.052419e-06,
  3.823036e-06, 1.722837e-06, 2.204176e-06, 2.273771e-06, 1.405613e-06, 
    2.315569e-06, 2.078667e-06, 2.647844e-06, 3.857057e-06, 1.059463e-05, 
    2.449346e-05, 3.355649e-05, 3.444398e-05, 1.858728e-05, 1.108764e-05,
  5.232086e-06, 2.482222e-06, 2.120563e-06, 9.907995e-07, 4.684273e-07, 
    2.670209e-07, 9.218193e-07, 1.665502e-06, 2.605895e-06, 4.361797e-06, 
    1.326324e-05, 2.732466e-05, 3.239726e-05, 2.653765e-05, 1.551077e-05,
  1.469253e-05, 1.40163e-05, 9.697645e-06, 2.069293e-06, 7.75413e-07, 
    2.253259e-06, 5.82697e-08, 2.958585e-07, 7.874264e-07, 1.629659e-06, 
    2.906928e-06, 1.164672e-05, 2.451922e-05, 3.267221e-05, 2.197865e-05,
  1.727625e-05, 1.787983e-05, 1.610623e-05, 2.155446e-06, 1.018584e-06, 
    1.060212e-06, 1.487366e-06, 8.257927e-08, 8.39409e-08, 1.500305e-06, 
    1.614224e-06, 3.215107e-06, 1.070458e-05, 2.531942e-05, 2.790932e-05,
  2.503722e-05, 1.91714e-05, 2.041499e-05, 2.967036e-06, 2.198851e-06, 
    1.826794e-06, 2.044904e-06, 2.151331e-06, 3.415986e-06, 2.049169e-06, 
    2.687041e-06, 1.864304e-06, 2.848835e-06, 1.544285e-05, 2.835187e-05,
  3.044366e-05, 2.771818e-05, 2.079203e-05, 6.830613e-06, 9.339456e-06, 
    1.881258e-06, 2.889221e-06, 3.549088e-06, 2.335091e-06, 1.35121e-06, 
    1.074721e-06, 1.068414e-06, 1.184083e-06, 4.810095e-06, 2.195123e-05,
  3.564577e-05, 3.625392e-05, 2.317411e-05, 1.352968e-05, 9.56525e-06, 
    2.860366e-06, 2.665161e-06, 3.26491e-06, 2.920588e-06, 1.656448e-06, 
    1.049178e-06, 1.191714e-06, 1.072693e-06, 1.542606e-06, 8.505226e-06,
  3.979902e-05, 4.084666e-05, 3.001386e-05, 9.130778e-06, 8.880575e-06, 
    4.07709e-06, 3.380457e-06, 3.002475e-06, 2.808185e-06, 1.848268e-06, 
    1.405174e-06, 1.070136e-06, 1.221202e-06, 8.560918e-07, 4.147924e-06,
  4.423504e-05, 4.132604e-05, 2.842616e-05, 2.443813e-06, 3.22052e-06, 
    6.298375e-06, 4.001747e-06, 4.490335e-06, 4.33632e-06, 3.725397e-06, 
    1.550007e-06, 1.142719e-06, 9.107201e-07, 9.147846e-07, 3.854056e-06,
  3.296093e-05, 2.239185e-05, 1.072381e-05, 8.602588e-07, 1.359883e-06, 
    4.440075e-06, 5.437851e-06, 9.599296e-06, 8.575014e-06, 3.751373e-06, 
    1.571621e-06, 7.843593e-07, 5.573798e-07, 8.179219e-07, 2.622607e-06,
  1.036346e-05, 1.360376e-05, 2.481936e-05, 1.585209e-05, 1.685585e-05, 
    1.81655e-05, 8.874928e-06, 1.084374e-06, 4.586457e-07, 7.286239e-07, 
    4.338559e-07, 3.284416e-07, 6.252796e-06, 1.510548e-05, 1.615662e-05,
  1.119172e-05, 9.357195e-06, 1.37781e-05, 1.758245e-05, 1.509957e-05, 
    2.341924e-05, 8.253883e-06, 3.759668e-07, 3.184863e-07, 5.120792e-07, 
    4.087873e-07, 3.89433e-07, 4.326457e-07, 3.312893e-06, 9.599643e-06,
  2.73434e-05, 2.76329e-05, 2.314893e-05, 1.005164e-05, 1.553409e-05, 
    2.752692e-05, 1.889557e-05, 1.38869e-06, 1.049718e-06, 4.142709e-07, 
    5.936309e-07, 5.095709e-07, 3.250611e-07, 8.352626e-07, 7.032056e-06,
  4.083438e-05, 4.346398e-05, 3.969638e-05, 1.491101e-05, 1.549417e-05, 
    2.102976e-05, 2.26428e-05, 5.385126e-06, 2.836296e-06, 1.285035e-06, 
    1.507062e-06, 6.126218e-07, 6.446154e-07, 5.317975e-07, 5.187976e-06,
  4.286005e-05, 3.804749e-05, 3.836197e-05, 4.25552e-06, 1.182079e-05, 
    2.357537e-05, 1.580712e-05, 8.805299e-06, 5.517543e-06, 5.925048e-07, 
    2.183015e-06, 6.358276e-07, 3.411167e-07, 3.716581e-07, 5.011133e-06,
  4.719413e-05, 3.620649e-05, 3.188103e-05, 1.500135e-05, 1.513138e-05, 
    1.395509e-05, 2.14386e-05, 8.585695e-06, 8.529556e-07, 2.062883e-07, 
    5.028103e-07, 5.299337e-07, 3.795314e-07, 2.961817e-07, 1.864357e-06,
  4.610274e-05, 4.705646e-05, 3.886412e-05, 2.32709e-05, 1.45475e-05, 
    5.466135e-06, 1.093817e-05, 1.077893e-05, 3.9524e-06, 1.245871e-06, 
    1.098131e-06, 1.041297e-06, 7.719915e-07, 2.390306e-07, 4.621059e-07,
  5.787944e-05, 5.332554e-05, 4.313867e-05, 2.293134e-05, 1.379623e-05, 
    6.400764e-06, 5.807088e-06, 4.203606e-06, 2.729658e-06, 2.172636e-06, 
    1.320552e-06, 1.497271e-06, 7.790243e-07, 2.273655e-07, 4.042923e-07,
  5.795346e-05, 5.514608e-05, 3.714349e-05, 1.305042e-05, 7.986494e-06, 
    5.546428e-06, 6.445732e-06, 6.040099e-06, 4.095583e-06, 2.31147e-06, 
    1.050234e-06, 1.416139e-06, 4.471771e-07, 2.420637e-07, 5.058898e-07,
  3.879571e-05, 2.271585e-05, 2.327551e-05, 1.447414e-05, 6.821438e-06, 
    6.990836e-06, 6.644602e-06, 6.919451e-06, 5.254493e-06, 2.16782e-06, 
    7.922299e-07, 1.209045e-06, 4.952789e-07, 2.184421e-07, 4.751644e-07,
  7.528243e-06, 1.446315e-06, 2.434826e-06, 2.262369e-06, 2.14769e-06, 
    3.616951e-06, 1.114268e-05, 1.523413e-05, 1.13557e-05, 5.034968e-06, 
    2.546715e-06, 1.195922e-06, 4.745231e-06, 1.49068e-05, 7.316783e-06,
  1.612865e-05, 5.285975e-06, 1.544466e-06, 4.129111e-06, 6.624329e-06, 
    1.567154e-05, 2.456007e-05, 1.935913e-05, 1.404894e-05, 6.90858e-06, 
    2.06976e-06, 4.734865e-07, 5.382559e-06, 1.561649e-05, 1.027983e-05,
  3.255886e-05, 3.482883e-05, 2.705075e-05, 8.844693e-06, 2.117623e-05, 
    2.549434e-05, 3.965773e-05, 3.366292e-05, 1.71038e-05, 4.894079e-06, 
    9.385685e-07, 6.146185e-07, 5.733202e-06, 1.871468e-05, 9.504618e-06,
  4.249178e-05, 4.442212e-05, 4.354524e-05, 1.545418e-05, 1.371496e-05, 
    1.383258e-05, 2.945132e-05, 3.001557e-05, 7.30953e-06, 2.535631e-06, 
    1.187597e-06, 7.591621e-07, 6.387875e-06, 1.52229e-05, 6.707423e-06,
  5.130782e-05, 4.902794e-05, 4.162485e-05, 7.452168e-06, 1.577248e-06, 
    7.344394e-06, 1.735911e-05, 1.096811e-05, 2.531563e-06, 1.161019e-06, 
    1.361019e-06, 9.949189e-07, 7.918285e-06, 1.171788e-05, 5.437718e-06,
  5.455736e-05, 5.70782e-05, 4.628299e-05, 1.621962e-05, 5.839102e-06, 
    2.34199e-06, 1.892278e-05, 9.405491e-06, 6.244283e-07, 8.754186e-07, 
    9.740389e-07, 1.506899e-06, 5.372193e-06, 6.859064e-06, 5.384763e-06,
  5.459883e-05, 6.420424e-05, 6.116135e-05, 3.364755e-05, 1.261837e-05, 
    2.751327e-06, 1.202968e-05, 1.459076e-05, 1.72946e-06, 1.265919e-06, 
    1.814428e-06, 2.113854e-06, 3.503101e-06, 5.650661e-06, 6.927757e-06,
  5.457462e-05, 6.151434e-05, 5.422429e-05, 3.39173e-05, 1.866792e-05, 
    1.137819e-05, 1.029524e-05, 5.164635e-06, 6.677683e-07, 2.411643e-06, 
    2.451962e-06, 3.694953e-06, 5.828005e-06, 7.242197e-06, 7.300567e-06,
  3.81868e-05, 4.593965e-05, 3.345068e-05, 1.938471e-05, 1.32838e-05, 
    1.129551e-05, 7.065895e-06, 1.463857e-06, 3.223007e-07, 1.818908e-06, 
    2.232792e-06, 4.461019e-06, 6.912608e-06, 6.498795e-06, 3.839779e-06,
  1.557918e-05, 1.257006e-05, 1.240801e-05, 1.092262e-05, 5.17454e-06, 
    2.648219e-06, 2.15417e-06, 2.020126e-06, 1.057492e-06, 1.542339e-06, 
    2.248254e-06, 3.781749e-06, 5.182141e-06, 4.588097e-06, 3.386362e-06,
  3.292527e-06, 5.734955e-08, 1.295232e-07, 4.857708e-08, 4.048519e-06, 
    9.66181e-06, 4.655707e-06, 6.025221e-07, 1.055885e-05, 5.452209e-05, 
    3.57853e-05, 1.541386e-05, 1.061291e-05, 5.460783e-06, 1.19437e-06,
  1.398212e-05, 1.995626e-06, 3.662454e-07, 8.472109e-07, 7.871649e-06, 
    1.457547e-05, 9.66577e-06, 4.810332e-06, 2.114518e-05, 3.879038e-05, 
    1.999221e-05, 9.277997e-06, 4.778016e-06, 1.723537e-06, 1.136958e-06,
  2.905924e-05, 2.161065e-05, 1.277884e-05, 2.657395e-06, 6.045068e-06, 
    1.604977e-05, 1.615227e-05, 1.762682e-05, 2.464797e-05, 2.484825e-05, 
    6.413655e-06, 3.556189e-06, 1.963622e-06, 4.906129e-07, 4.249999e-07,
  3.069475e-05, 2.692691e-05, 1.578927e-05, 4.813944e-06, 4.433013e-06, 
    1.151461e-05, 2.308534e-05, 2.71505e-05, 3.037892e-05, 2.154262e-05, 
    2.589233e-06, 7.534198e-07, 1.24184e-06, 7.932331e-07, 1.417205e-06,
  3.36261e-05, 2.104814e-05, 1.324541e-05, 2.321099e-06, 2.316746e-06, 
    9.134583e-06, 1.233277e-05, 4.76415e-06, 1.28316e-05, 9.238175e-06, 
    1.423202e-06, 3.864123e-07, 1.674765e-06, 2.289295e-06, 2.220255e-06,
  3.803916e-05, 2.679455e-05, 1.709909e-05, 7.768039e-06, 4.523618e-06, 
    2.01426e-06, 3.734376e-06, 2.652005e-06, 1.118229e-06, 1.641779e-06, 
    9.941945e-07, 1.318152e-06, 6.676422e-06, 6.72483e-06, 2.84363e-06,
  3.887402e-05, 3.898483e-05, 2.520305e-05, 1.005716e-05, 4.871879e-06, 
    1.7516e-06, 1.563863e-06, 1.951823e-06, 1.850995e-06, 8.076502e-07, 
    7.973737e-07, 3.836462e-06, 9.452622e-06, 7.071502e-06, 2.533354e-06,
  3.634424e-05, 4.086846e-05, 2.373827e-05, 1.00171e-05, 7.350951e-06, 
    2.432289e-06, 1.902244e-06, 1.25948e-06, 8.820438e-07, 1.217381e-06, 
    4.050309e-06, 9.4794e-06, 9.987806e-06, 6.120271e-06, 5.163393e-06,
  2.26961e-05, 2.465637e-05, 1.502509e-05, 8.206363e-06, 3.787861e-06, 
    3.544382e-06, 2.947006e-06, 2.878321e-06, 4.304604e-06, 9.443647e-06, 
    1.674718e-05, 1.775188e-05, 1.026903e-05, 5.180252e-06, 5.46927e-06,
  8.251242e-06, 7.844588e-06, 7.819345e-06, 6.827952e-06, 3.389176e-06, 
    4.48139e-06, 7.553874e-06, 1.301371e-05, 1.835902e-05, 2.525477e-05, 
    2.709822e-05, 1.88154e-05, 7.553695e-06, 5.883565e-06, 5.267404e-06,
  2.898717e-06, 1.357256e-07, 6.958245e-08, 1.498683e-06, 9.395266e-06, 
    2.625244e-05, 4.793517e-05, 4.216493e-05, 2.572031e-05, 2.124036e-05, 
    2.918977e-05, 7.369843e-05, 7.74613e-05, 3.925146e-05, 1.843908e-05,
  7.558808e-06, 1.718726e-07, 2.851523e-07, 2.631039e-06, 9.051459e-06, 
    2.2169e-05, 4.720248e-05, 4.903386e-05, 3.50634e-05, 3.856812e-05, 
    6.266893e-05, 7.064889e-05, 4.054882e-05, 2.24851e-05, 1.129477e-05,
  2.608262e-05, 1.055124e-05, 5.150415e-06, 2.695944e-06, 3.469645e-06, 
    9.905069e-06, 3.618771e-05, 6.261298e-05, 5.257616e-05, 3.955854e-05, 
    3.326119e-05, 3.008116e-05, 2.404346e-05, 1.745535e-05, 1.385699e-05,
  3.005619e-05, 1.721676e-05, 1.112396e-05, 2.949321e-06, 3.431205e-06, 
    8.475981e-06, 1.827267e-05, 1.671576e-05, 2.145009e-05, 2.374686e-05, 
    1.599407e-05, 8.070751e-06, 7.323173e-06, 1.226444e-05, 1.313567e-05,
  2.646152e-05, 2.123364e-05, 1.226498e-05, 1.728546e-06, 2.95703e-06, 
    9.203402e-06, 6.175153e-06, 2.395293e-06, 4.217765e-06, 2.557856e-06, 
    1.47339e-06, 4.541643e-07, 3.693925e-07, 2.158342e-06, 6.016266e-06,
  3.054748e-05, 2.623643e-05, 1.834208e-05, 7.762389e-06, 4.935257e-06, 
    4.009736e-06, 4.077767e-06, 3.141953e-06, 2.297615e-06, 2.329092e-06, 
    2.088267e-06, 1.210866e-06, 3.566193e-07, 4.22934e-07, 1.829853e-06,
  2.849091e-05, 2.739203e-05, 2.336584e-05, 1.194727e-05, 6.981873e-06, 
    4.693655e-06, 1.840367e-06, 3.268515e-06, 2.995027e-06, 1.88779e-06, 
    1.866536e-06, 2.009608e-06, 9.329672e-07, 1.421984e-07, 2.09325e-06,
  2.397311e-05, 2.581124e-05, 1.230213e-05, 1.134372e-05, 8.555475e-06, 
    5.064493e-06, 8.829943e-07, 2.140609e-06, 3.618506e-06, 3.328185e-06, 
    2.81244e-06, 2.153495e-06, 7.539465e-07, 9.696142e-07, 3.112848e-06,
  1.472081e-05, 1.406697e-05, 6.995674e-06, 6.233252e-06, 5.861046e-06, 
    3.408277e-06, 2.790145e-06, 1.436311e-06, 3.554064e-06, 4.574599e-06, 
    3.799669e-06, 2.988626e-06, 3.258891e-06, 3.187959e-06, 3.916128e-06,
  3.794487e-06, 2.22587e-06, 2.022351e-06, 2.389183e-06, 5.468324e-06, 
    1.046363e-05, 1.277559e-05, 1.568698e-05, 9.398338e-06, 5.462684e-06, 
    3.713042e-06, 4.550453e-06, 3.515921e-06, 5.01868e-06, 4.296347e-06,
  5.323516e-07, 1.277419e-07, 1.644544e-06, 2.779366e-06, 3.593812e-06, 
    2.2623e-06, 1.184345e-06, 1.184347e-06, 4.142381e-06, 9.64064e-06, 
    2.005407e-05, 1.024778e-05, 4.500026e-06, 4.953749e-06, 3.961036e-06,
  3.876926e-06, 6.246534e-07, 6.358787e-07, 2.020022e-06, 1.745354e-06, 
    7.481898e-07, 5.653611e-07, 6.476265e-07, 1.395245e-06, 8.743399e-06, 
    2.0474e-05, 2.585025e-05, 6.080733e-06, 4.775279e-06, 4.319269e-06,
  1.117965e-05, 1.07573e-05, 7.46861e-06, 2.036048e-06, 6.64049e-07, 
    1.064054e-06, 3.02207e-07, 6.397585e-07, 6.841312e-07, 2.103672e-06, 
    1.675206e-05, 4.346582e-05, 2.010099e-05, 2.783993e-06, 3.076174e-06,
  1.369987e-05, 1.615334e-05, 1.430994e-05, 2.385181e-06, 1.722708e-06, 
    2.877811e-06, 5.027799e-06, 6.570021e-07, 4.258827e-07, 1.088411e-06, 
    5.50501e-06, 3.0867e-05, 4.223803e-05, 2.087944e-05, 9.370398e-06,
  1.368079e-05, 1.485728e-05, 1.297178e-05, 1.336365e-06, 2.93399e-06, 
    6.847153e-06, 8.461397e-06, 1.280995e-05, 1.196139e-05, 1.991645e-06, 
    6.985001e-06, 1.433353e-05, 3.181936e-05, 2.604738e-05, 1.770886e-05,
  1.103966e-05, 1.318467e-05, 1.050242e-05, 7.093404e-06, 6.157145e-06, 
    7.542047e-06, 1.298965e-05, 1.047669e-05, 6.346706e-06, 5.749377e-06, 
    5.252555e-06, 7.565513e-06, 1.820781e-05, 2.153951e-05, 1.751746e-05,
  6.866665e-06, 1.193934e-05, 1.190734e-05, 1.331869e-05, 1.051227e-05, 
    6.707584e-06, 1.113318e-05, 1.121063e-05, 6.362132e-06, 3.704291e-06, 
    3.727654e-06, 5.603398e-06, 1.142532e-05, 1.596005e-05, 1.626657e-05,
  5.567697e-06, 1.29756e-05, 2.23788e-05, 2.66888e-05, 1.130455e-05, 
    4.56928e-06, 8.986112e-06, 1.202879e-05, 7.521045e-06, 5.151893e-06, 
    4.120964e-06, 3.658136e-06, 8.810186e-06, 1.170538e-05, 1.624058e-05,
  1.3009e-05, 2.256759e-05, 3.963885e-05, 2.78499e-05, 6.567406e-06, 
    2.491728e-06, 9.122941e-06, 1.287135e-05, 8.972473e-06, 6.291833e-06, 
    4.350223e-06, 3.868162e-06, 5.257569e-06, 7.575064e-06, 9.833291e-06,
  2.076958e-05, 2.294534e-05, 2.222091e-05, 8.940188e-06, 1.204208e-06, 
    1.691511e-06, 8.059924e-06, 1.453837e-05, 1.022704e-05, 5.22073e-06, 
    4.976749e-06, 4.303528e-06, 4.227956e-06, 6.664054e-06, 5.534073e-06,
  3.156184e-07, 1.807282e-06, 3.808477e-06, 2.495993e-06, 1.536956e-06, 
    5.40334e-06, 1.890624e-05, 1.560808e-05, 2.781654e-06, 4.877565e-06, 
    1.467418e-05, 9.73091e-06, 3.083955e-06, 3.649606e-06, 1.111391e-05,
  1.109473e-06, 2.385802e-06, 2.106078e-06, 1.473223e-06, 2.313792e-06, 
    1.075905e-05, 2.62326e-05, 1.251777e-05, 1.539587e-06, 6.058102e-06, 
    1.124377e-05, 9.292037e-06, 2.639526e-06, 9.103175e-07, 2.71025e-06,
  1.485218e-06, 2.916562e-06, 2.63963e-06, 3.619959e-06, 8.633775e-06, 
    2.50631e-05, 2.096622e-05, 1.084777e-05, 1.131901e-06, 6.215093e-06, 
    1.148469e-05, 9.11693e-06, 3.109155e-06, 4.740142e-07, 9.75034e-08,
  1.793386e-06, 3.264255e-06, 5.083843e-06, 6.068235e-06, 2.30153e-05, 
    3.382811e-05, 2.771163e-05, 3.728297e-06, 5.117324e-07, 5.346499e-06, 
    1.080153e-05, 1.092712e-05, 6.84836e-06, 2.687164e-06, 1.443574e-07,
  2.0328e-06, 3.284924e-06, 6.291843e-06, 1.031499e-05, 3.816497e-05, 
    3.892391e-05, 1.070317e-05, 2.735153e-06, 6.280241e-06, 5.040283e-06, 
    1.104317e-05, 9.732056e-06, 1.413611e-05, 9.937722e-06, 4.742109e-06,
  2.797538e-06, 4.239166e-06, 6.940984e-06, 2.478969e-05, 4.472362e-05, 
    2.620594e-05, 5.022292e-06, 2.088542e-06, 2.457344e-06, 5.733789e-06, 
    5.627317e-06, 7.49123e-06, 1.174361e-05, 1.94632e-05, 2.184172e-05,
  7.579746e-06, 6.419939e-06, 1.400986e-05, 4.066253e-05, 3.627884e-05, 
    6.666571e-06, 1.907922e-06, 3.543454e-06, 4.33141e-06, 5.16989e-06, 
    5.057566e-06, 5.865274e-06, 7.341663e-06, 1.611346e-05, 3.272553e-05,
  1.037792e-05, 1.147903e-05, 2.047236e-05, 3.02731e-05, 1.18384e-05, 
    3.225928e-07, 1.020043e-06, 4.704448e-06, 3.704356e-06, 4.49757e-06, 
    5.267837e-06, 5.125835e-06, 6.293076e-06, 9.224111e-06, 2.148271e-05,
  1.290395e-05, 1.217902e-05, 8.397769e-06, 5.692709e-06, 1.035192e-06, 
    9.06909e-08, 2.641946e-06, 5.693264e-06, 6.326152e-06, 5.144697e-06, 
    5.554875e-06, 4.600591e-06, 7.124866e-06, 7.713465e-06, 1.018028e-05,
  5.731024e-06, 5.556336e-06, 3.141272e-06, 1.402443e-06, 1.059724e-06, 
    1.429849e-07, 3.54666e-06, 7.389069e-06, 8.435556e-06, 4.354943e-06, 
    4.437004e-06, 3.443902e-06, 8.486231e-06, 7.837415e-06, 8.496941e-06,
  1.543435e-06, 2.992006e-06, 5.688071e-06, 7.348355e-06, 7.208627e-06, 
    1.062819e-05, 9.920059e-06, 7.316326e-06, 5.313528e-06, 1.480563e-06, 
    8.239836e-07, 4.082977e-06, 3.325903e-06, 5.521421e-07, 2.083148e-06,
  2.118912e-06, 5.076282e-06, 6.902759e-06, 5.965581e-06, 5.025163e-06, 
    6.528333e-06, 6.376831e-06, 3.224033e-06, 2.701555e-06, 8.132173e-07, 
    7.604668e-07, 4.780743e-06, 5.446217e-06, 4.082616e-06, 1.110587e-06,
  3.324517e-06, 4.685681e-06, 5.6463e-06, 4.135304e-06, 2.035418e-06, 
    5.215838e-06, 2.293768e-06, 2.947083e-06, 7.330193e-07, 3.80613e-07, 
    1.087998e-06, 4.415562e-06, 7.34359e-06, 8.922819e-06, 5.602761e-06,
  3.542878e-06, 5.473011e-06, 5.210865e-06, 2.051257e-06, 5.475555e-07, 
    7.967345e-07, 1.021923e-06, 1.095975e-06, 3.209103e-07, 6.213775e-07, 
    6.349459e-07, 3.836683e-06, 1.065308e-05, 1.251287e-05, 7.600436e-06,
  3.680271e-06, 3.480943e-06, 2.131875e-06, 6.486439e-07, 7.430297e-07, 
    1.303543e-06, 2.02777e-06, 2.455876e-06, 2.057217e-06, 1.147098e-06, 
    5.751916e-06, 4.154211e-06, 8.738986e-06, 1.305961e-05, 1.336543e-05,
  8.344194e-06, 4.390176e-06, 4.389308e-06, 2.498998e-06, 1.365588e-06, 
    2.101776e-06, 4.046542e-06, 4.479223e-06, 4.776629e-06, 2.696555e-06, 
    4.073824e-06, 1.861382e-06, 9.150152e-06, 1.297634e-05, 1.151874e-05,
  7.582512e-06, 8.601054e-06, 1.195515e-05, 7.924447e-06, 3.328704e-06, 
    2.349566e-06, 4.116174e-06, 5.963641e-06, 7.375565e-06, 6.737183e-06, 
    7.047554e-06, 2.648663e-06, 1.032465e-05, 1.149508e-05, 1.167878e-05,
  1.07683e-05, 1.150683e-05, 1.017349e-05, 1.220003e-05, 3.887095e-06, 
    1.515062e-06, 4.064539e-06, 5.93732e-06, 4.892334e-06, 7.734679e-06, 
    6.948925e-06, 5.350943e-06, 9.208563e-06, 9.549319e-06, 1.358778e-05,
  1.173609e-05, 1.43891e-05, 6.674452e-06, 1.264869e-05, 7.791195e-06, 
    1.095246e-06, 3.278209e-06, 7.646722e-06, 5.042938e-06, 6.55714e-06, 
    1.01525e-05, 8.209398e-06, 1.119622e-05, 1.298343e-05, 1.111334e-05,
  6.639925e-06, 6.761882e-06, 6.656212e-06, 1.10782e-05, 8.05979e-06, 
    7.406612e-07, 3.617925e-06, 1.002968e-05, 8.472523e-06, 7.362145e-06, 
    1.029738e-05, 9.979448e-06, 1.352283e-05, 1.19502e-05, 4.452745e-06,
  3.215561e-07, 2.049615e-07, 1.09823e-06, 4.217547e-06, 1.008369e-05, 
    7.587405e-06, 1.407202e-06, 2.149964e-06, 3.373489e-06, 5.395998e-06, 
    5.635868e-06, 5.075245e-06, 6.816713e-06, 5.009585e-06, 5.985041e-06,
  1.42725e-07, 8.464364e-07, 3.521363e-06, 1.386715e-05, 1.957349e-05, 
    1.212835e-05, 2.247518e-06, 5.933703e-07, 1.705629e-06, 3.798267e-06, 
    5.780422e-06, 7.845866e-06, 6.828348e-06, 6.862384e-06, 5.004872e-06,
  6.646462e-07, 3.289919e-06, 7.186494e-06, 1.754973e-05, 1.992434e-05, 
    1.637798e-05, 1.284353e-06, 8.500168e-07, 2.047139e-06, 2.119529e-06, 
    3.675501e-06, 9.123585e-06, 9.501859e-06, 8.948919e-06, 6.656277e-06,
  1.220261e-06, 3.689985e-06, 1.199091e-05, 2.12032e-05, 1.917678e-05, 
    9.321382e-06, 4.747669e-06, 5.176364e-07, 1.74738e-06, 5.477984e-06, 
    8.154086e-06, 8.883001e-06, 9.441746e-06, 5.856224e-06, 6.998355e-06,
  2.722694e-06, 5.738849e-06, 1.726977e-05, 2.401865e-05, 1.436975e-05, 
    4.76159e-06, 4.966053e-06, 7.16611e-06, 1.220599e-05, 7.358246e-06, 
    1.226996e-05, 7.429725e-06, 7.505235e-06, 3.451752e-06, 7.68579e-06,
  4.740108e-06, 6.953398e-06, 1.777113e-05, 1.980248e-05, 1.020475e-05, 
    3.285646e-06, 3.275134e-06, 6.449662e-06, 8.743288e-06, 8.059457e-06, 
    9.291128e-06, 8.199452e-06, 8.079075e-06, 8.303552e-06, 7.174278e-06,
  6.195709e-06, 5.925664e-06, 1.076247e-05, 1.418046e-05, 7.500093e-06, 
    2.659126e-06, 1.687099e-06, 5.864336e-06, 5.820405e-06, 8.107652e-06, 
    8.390381e-06, 8.26736e-06, 1.052028e-05, 1.122275e-05, 9.616949e-06,
  1.00384e-05, 5.380807e-06, 5.975739e-06, 4.954682e-06, 4.987147e-06, 
    1.16215e-06, 2.052053e-06, 4.981421e-06, 5.626207e-06, 9.050165e-06, 
    9.793655e-06, 1.337881e-05, 1.675383e-05, 1.600675e-05, 1.371636e-05,
  1.345146e-05, 5.611921e-06, 2.884998e-06, 3.506012e-06, 2.883068e-06, 
    7.580072e-07, 2.925286e-06, 4.460692e-06, 5.053355e-06, 7.386171e-06, 
    1.088366e-05, 1.693357e-05, 2.202123e-05, 2.303777e-05, 2.277378e-05,
  1.065421e-05, 7.786193e-06, 1.653294e-06, 3.117382e-06, 4.938846e-07, 
    8.283479e-07, 2.446548e-06, 6.464751e-06, 5.981298e-06, 5.231069e-06, 
    7.713187e-06, 1.46416e-05, 2.35733e-05, 2.920553e-05, 3.863197e-05,
  8.713056e-07, 3.954883e-06, 6.830134e-06, 7.684704e-06, 7.732163e-06, 
    9.361038e-06, 7.482475e-06, 3.003411e-06, 1.450124e-06, 2.861144e-06, 
    4.800856e-06, 5.6202e-06, 8.911518e-06, 7.826965e-06, 6.687508e-06,
  1.131194e-06, 3.136627e-06, 4.462481e-06, 4.778419e-06, 3.399985e-06, 
    4.025989e-06, 3.339464e-06, 8.293194e-07, 5.893386e-07, 1.085762e-06, 
    4.296339e-06, 8.350937e-06, 8.210082e-06, 1.242846e-05, 6.363053e-06,
  2.485856e-06, 2.826721e-06, 4.358097e-06, 2.771756e-06, 7.270388e-07, 
    2.617711e-06, 3.009385e-07, 1.251122e-06, 1.336609e-06, 4.956204e-06, 
    7.996295e-06, 1.013023e-05, 9.430782e-06, 1.084886e-05, 9.6763e-06,
  3.743073e-06, 2.305869e-06, 6.004716e-06, 1.76225e-06, 9.05417e-07, 
    1.503785e-06, 2.497504e-06, 3.455023e-07, 6.267672e-07, 1.646435e-06, 
    7.793597e-06, 1.14632e-05, 1.205789e-05, 1.196875e-05, 1.426607e-05,
  7.599352e-06, 3.445971e-06, 6.539876e-06, 1.476099e-06, 2.474324e-07, 
    2.402804e-06, 1.897871e-06, 5.197558e-06, 7.976014e-06, 1.832977e-06, 
    1.143505e-05, 1.004454e-05, 1.255554e-05, 1.242007e-05, 1.335429e-05,
  1.064481e-05, 3.519277e-06, 5.536758e-06, 2.249839e-06, 2.542722e-06, 
    1.607096e-06, 9.395628e-07, 9.723568e-07, 1.661518e-06, 4.196352e-06, 
    1.026087e-05, 1.202447e-05, 1.208792e-05, 1.364161e-05, 1.335686e-05,
  9.970053e-06, 3.715864e-06, 5.727615e-06, 2.113938e-06, 2.740554e-06, 
    9.714699e-07, 3.193143e-07, 8.108063e-07, 8.00518e-07, 2.142213e-06, 
    5.567463e-06, 1.194963e-05, 1.005626e-05, 1.189651e-05, 1.190699e-05,
  1.380317e-05, 3.951166e-06, 3.398557e-07, 2.76038e-06, 2.622786e-06, 
    1.413825e-06, 1.557217e-07, 2.661444e-07, 6.877062e-07, 1.360234e-06, 
    2.317289e-06, 1.045231e-05, 1.013445e-05, 1.301333e-05, 1.029672e-05,
  1.497143e-05, 4.21616e-06, 1.957247e-07, 1.077453e-06, 3.228658e-06, 
    9.361463e-07, 2.260387e-07, 2.467196e-07, 4.737921e-07, 7.546746e-07, 
    1.169522e-06, 6.708837e-06, 1.393417e-05, 1.487375e-05, 2.319506e-05,
  1.155281e-05, 5.454936e-06, 7.921876e-07, 9.157948e-07, 3.819666e-06, 
    2.826215e-06, 2.458816e-07, 4.678452e-07, 2.649e-07, 4.283511e-07, 
    8.023864e-07, 3.631927e-06, 1.367452e-05, 1.563034e-05, 2.782737e-05,
  1.755342e-07, 3.693575e-08, 1.885437e-07, 7.12518e-08, 7.839323e-08, 
    1.153617e-07, 3.756604e-07, 2.201743e-07, 1.646792e-07, 9.542601e-07, 
    1.534558e-06, 8.300324e-07, 4.097426e-06, 5.851371e-06, 5.770988e-06,
  6.078334e-07, 1.401939e-07, 8.603056e-08, 1.242806e-07, 1.170803e-07, 
    1.738134e-07, 1.628842e-07, 2.527306e-07, 1.302392e-07, 1.221857e-07, 
    4.17927e-07, 2.283653e-06, 1.709856e-06, 5.726914e-06, 4.167016e-06,
  1.34336e-06, 1.735068e-06, 1.811736e-06, 9.192192e-07, 3.916518e-07, 
    6.76639e-07, 5.152517e-07, 2.343245e-07, 1.70104e-07, 2.08597e-07, 
    3.414819e-07, 1.609587e-06, 4.333059e-06, 6.224974e-06, 5.628613e-06,
  1.486276e-06, 4.192633e-06, 8.552086e-06, 4.656338e-06, 2.678532e-06, 
    1.433068e-06, 2.069253e-06, 4.22362e-07, 9.788252e-08, 3.873157e-07, 
    7.073596e-07, 1.957204e-06, 3.780631e-06, 6.101679e-06, 9.189072e-06,
  1.090016e-06, 5.950302e-06, 1.074602e-05, 7.50811e-06, 5.407789e-06, 
    5.103831e-06, 6.57358e-06, 4.924271e-06, 7.018867e-07, 1.350637e-06, 
    3.61635e-06, 3.883139e-06, 4.395656e-06, 5.64284e-06, 8.020791e-06,
  8.601058e-07, 7.749246e-06, 1.138645e-05, 9.781375e-06, 9.76143e-06, 
    9.307299e-06, 8.4825e-06, 5.000875e-06, 3.578432e-06, 6.956227e-06, 
    9.028734e-06, 7.070536e-06, 7.912556e-06, 6.301764e-06, 6.286053e-06,
  3.720542e-06, 7.930032e-06, 9.092426e-06, 5.923579e-06, 6.152767e-06, 
    6.329199e-06, 7.385226e-06, 1.052425e-05, 1.24207e-05, 1.167609e-05, 
    1.272003e-05, 9.956096e-06, 7.487959e-06, 7.223181e-06, 8.114638e-06,
  9.478859e-06, 8.69725e-06, 6.604937e-06, 4.855015e-06, 5.722913e-06, 
    6.159935e-06, 9.909905e-06, 1.240159e-05, 1.459995e-05, 1.448463e-05, 
    1.400151e-05, 9.169143e-06, 6.72277e-06, 1.057852e-05, 1.131189e-05,
  5.943016e-06, 4.651089e-06, 7.436043e-06, 6.276094e-06, 5.703423e-06, 
    7.839858e-06, 1.199107e-05, 1.630815e-05, 1.76372e-05, 1.383997e-05, 
    9.00082e-06, 7.580625e-06, 7.730479e-06, 1.167245e-05, 1.867656e-05,
  2.588337e-06, 5.354013e-06, 6.7889e-06, 6.552552e-06, 6.995861e-06, 
    7.911104e-06, 1.170765e-05, 1.752873e-05, 1.537549e-05, 1.096089e-05, 
    8.005075e-06, 6.478224e-06, 4.577631e-06, 1.128874e-05, 1.930935e-05,
  3.781741e-07, 1.237963e-06, 5.5337e-06, 9.679648e-06, 1.058393e-05, 
    7.191661e-06, 2.328265e-06, 9.259577e-07, 7.80928e-07, 1.005733e-06, 
    1.394693e-06, 8.390703e-07, 1.392735e-06, 2.496672e-06, 1.073756e-06,
  6.936139e-07, 2.113649e-06, 6.35909e-06, 1.162598e-05, 8.834611e-06, 
    4.87803e-06, 2.151424e-06, 1.084619e-06, 8.616763e-07, 7.855396e-07, 
    6.258423e-07, 9.599573e-07, 2.264525e-06, 3.999279e-06, 1.839546e-06,
  1.850352e-07, 1.521264e-06, 6.811038e-06, 1.223476e-05, 1.069279e-05, 
    6.14494e-06, 1.14749e-06, 3.208836e-06, 4.374134e-06, 3.290597e-06, 
    2.217723e-06, 2.211757e-06, 3.538829e-06, 4.442336e-06, 3.524817e-06,
  1.694048e-07, 1.299836e-07, 3.713213e-06, 9.598549e-06, 9.461483e-06, 
    7.527732e-06, 1.79858e-05, 3.367695e-06, 3.23946e-06, 5.198206e-06, 
    4.276774e-06, 2.936624e-06, 4.064075e-06, 6.506683e-06, 7.591039e-06,
  1.52554e-07, 8.887751e-08, 2.168337e-06, 6.03025e-06, 7.514971e-06, 
    1.331357e-05, 2.049797e-05, 3.521379e-05, 1.578509e-05, 6.52827e-06, 
    1.206431e-05, 1.036293e-05, 1.163945e-05, 1.426775e-05, 1.852617e-05,
  9.501427e-08, 6.571656e-07, 3.393928e-06, 6.406227e-06, 5.064465e-06, 
    5.966905e-06, 1.42519e-05, 2.021734e-05, 2.37644e-05, 2.804364e-05, 
    2.054597e-05, 1.822551e-05, 2.106415e-05, 2.245636e-05, 2.640003e-05,
  1.365918e-06, 4.748534e-06, 7.796994e-06, 8.216205e-06, 7.757308e-06, 
    1.408096e-05, 2.75617e-05, 4.014324e-05, 2.618998e-05, 1.641056e-05, 
    1.529979e-05, 1.874015e-05, 2.512732e-05, 2.848938e-05, 2.984308e-05,
  2.876123e-06, 4.093572e-06, 6.365388e-06, 7.374272e-06, 1.250982e-05, 
    2.642126e-05, 2.666043e-05, 8.545364e-06, 8.934364e-06, 1.354417e-05, 
    1.51343e-05, 1.566887e-05, 1.532614e-05, 1.548521e-05, 1.512192e-05,
  2.995182e-06, 3.656126e-06, 8.103116e-06, 1.054137e-05, 1.932532e-05, 
    2.505996e-05, 5.20964e-06, 5.910249e-06, 1.246048e-05, 1.417072e-05, 
    6.100379e-06, 4.975809e-06, 6.591538e-06, 1.172803e-05, 1.399344e-05,
  7.077655e-06, 8.897893e-06, 8.415237e-06, 1.390506e-05, 1.871489e-05, 
    6.488202e-06, 4.928981e-06, 9.80918e-06, 1.600453e-05, 1.028984e-05, 
    4.527337e-06, 4.063413e-06, 7.961256e-06, 1.321169e-05, 1.408649e-05,
  4.878432e-06, 6.320469e-06, 6.645233e-06, 7.40355e-06, 1.143562e-05, 
    9.865056e-06, 9.7685e-06, 4.379702e-06, 6.862185e-06, 7.441257e-06, 
    5.191076e-06, 3.299039e-06, 5.713394e-06, 5.302712e-06, 5.915094e-06,
  3.775703e-06, 3.85386e-06, 3.991315e-06, 5.83247e-06, 6.89032e-06, 
    4.662371e-06, 4.420113e-06, 3.850755e-06, 5.443421e-06, 1.125489e-05, 
    1.485787e-05, 1.390562e-05, 9.914324e-06, 1.302014e-05, 7.436976e-06,
  1.654487e-06, 2.910497e-06, 2.908676e-06, 3.787831e-06, 6.819105e-06, 
    7.252257e-06, 1.306007e-06, 4.979522e-06, 8.458135e-06, 1.499947e-05, 
    2.029667e-05, 2.686299e-05, 2.723608e-05, 2.293644e-05, 1.785007e-05,
  2.480451e-06, 2.664902e-06, 3.16429e-06, 5.384321e-06, 4.033062e-06, 
    1.102181e-05, 1.598501e-05, 2.197985e-06, 1.291084e-05, 3.049559e-05, 
    3.208499e-05, 3.232689e-05, 3.648525e-05, 3.719882e-05, 3.418984e-05,
  4.738322e-06, 4.408664e-06, 3.481152e-06, 3.312801e-06, 8.127306e-06, 
    1.346566e-05, 1.876798e-05, 2.594959e-05, 2.752894e-05, 2.614243e-05, 
    3.204732e-05, 1.965209e-05, 1.063513e-05, 4.829596e-06, 6.84815e-06,
  6.965286e-06, 5.373375e-06, 3.910638e-06, 3.489382e-06, 8.140807e-06, 
    1.152998e-05, 2.087715e-05, 2.699587e-05, 2.297563e-05, 1.220204e-05, 
    4.237481e-06, 1.482675e-06, 5.825194e-07, 1.958806e-07, 8.853519e-07,
  9.606641e-06, 5.824074e-06, 3.878974e-06, 5.420557e-06, 3.859335e-06, 
    4.491857e-06, 5.924459e-06, 4.773492e-06, 2.766624e-06, 1.391779e-06, 
    8.925024e-07, 7.913793e-07, 9.695102e-07, 9.702567e-07, 7.744725e-07,
  8.102078e-06, 2.857011e-06, 3.44958e-06, 2.658855e-06, 1.004491e-06, 
    4.073128e-07, 2.236381e-07, 1.204115e-06, 2.519202e-06, 3.761427e-06, 
    4.252487e-06, 6.806961e-06, 7.697318e-06, 9.84108e-06, 1.06753e-05,
  8.264749e-06, 4.315871e-06, 1.116037e-06, 9.709373e-07, 1.512068e-06, 
    9.425627e-07, 8.31017e-07, 4.954389e-06, 6.418692e-06, 1.067037e-05, 
    6.201181e-06, 4.854137e-06, 8.075305e-06, 8.4648e-06, 7.691016e-06,
  7.241079e-06, 3.186321e-06, 4.590457e-07, 8.051169e-07, 6.424104e-07, 
    4.179838e-07, 2.989645e-06, 5.476466e-06, 1.440994e-05, 1.085338e-05, 
    6.913308e-06, 3.892073e-06, 6.791963e-06, 1.131631e-05, 1.012695e-05,
  2.514019e-06, 2.028581e-06, 1.528356e-06, 2.473746e-06, 4.108772e-06, 
    3.619026e-06, 1.791916e-06, 1.805208e-06, 2.437225e-06, 4.805061e-06, 
    1.284084e-05, 1.865854e-05, 2.011748e-05, 1.914101e-05, 1.981994e-05,
  2.952366e-06, 2.539735e-06, 3.709131e-07, 1.354706e-07, 1.019088e-06, 
    1.439373e-06, 1.046597e-06, 8.951375e-07, 1.736801e-06, 3.038384e-06, 
    3.29926e-06, 1.153653e-05, 1.765662e-05, 2.337819e-05, 2.366644e-05,
  5.653335e-06, 4.611266e-06, 3.360344e-06, 1.475835e-07, 5.041271e-08, 
    1.721783e-06, 6.882274e-08, 1.625781e-07, 2.367506e-06, 1.000242e-06, 
    5.540012e-07, 2.863908e-06, 6.952709e-06, 1.685214e-05, 1.707135e-05,
  7.899918e-06, 6.101635e-06, 5.828168e-06, 3.601881e-06, 1.891268e-06, 
    5.997113e-07, 3.138584e-06, 9.546986e-08, 5.538513e-07, 5.555424e-06, 
    1.409214e-06, 5.677595e-07, 5.549257e-07, 2.830157e-06, 7.967198e-06,
  7.188409e-06, 6.538898e-06, 7.197375e-06, 3.856665e-06, 3.385531e-06, 
    4.288583e-06, 3.652533e-06, 4.874527e-06, 1.343093e-05, 8.630304e-06, 
    4.783438e-06, 2.358521e-06, 2.724985e-07, 6.325507e-08, 8.04164e-07,
  9.371713e-06, 7.485931e-06, 7.000785e-06, 5.849617e-06, 4.692403e-06, 
    1.828198e-06, 4.389577e-06, 7.398023e-06, 9.798255e-06, 5.874771e-06, 
    1.371107e-06, 4.93573e-06, 3.773073e-06, 4.078771e-07, 1.45044e-07,
  7.95854e-06, 7.256165e-06, 9.175111e-06, 5.404362e-06, 5.576398e-06, 
    1.002513e-06, 3.653444e-06, 5.088924e-06, 3.545601e-06, 5.372989e-06, 
    4.72202e-06, 4.639247e-06, 8.307076e-06, 4.530646e-06, 4.183126e-07,
  7.298588e-06, 1.284558e-05, 1.08886e-05, 5.420007e-06, 5.971358e-06, 
    1.301265e-06, 5.836954e-06, 6.572974e-06, 3.421313e-06, 3.709273e-06, 
    4.334709e-06, 6.58624e-06, 6.579597e-06, 5.451142e-06, 6.063033e-06,
  1.207949e-05, 1.392345e-05, 9.280138e-06, 4.269275e-06, 8.605283e-06, 
    3.168313e-06, 5.617103e-06, 7.77081e-06, 8.829566e-06, 1.185977e-05, 
    5.445032e-06, 6.861902e-06, 4.158199e-06, 6.155454e-06, 8.272576e-06,
  1.022263e-05, 1.248589e-05, 6.898865e-06, 5.656462e-06, 1.140926e-05, 
    6.031389e-06, 6.604143e-06, 6.243949e-06, 9.002672e-06, 1.035217e-05, 
    6.630079e-06, 8.306211e-06, 1.363605e-06, 3.270536e-06, 3.502376e-06,
  3.862832e-06, 4.650759e-06, 3.768082e-06, 1.262223e-06, 3.919595e-06, 
    1.786157e-05, 2.678162e-05, 2.391565e-05, 1.413255e-05, 4.223184e-06, 
    1.083457e-06, 1.807675e-07, 9.319e-07, 4.10453e-06, 6.886479e-06,
  2.926439e-06, 3.492507e-06, 4.067575e-06, 2.95474e-06, 1.071337e-05, 
    2.066267e-05, 2.302523e-05, 2.457367e-05, 1.823842e-05, 7.629724e-06, 
    1.248147e-06, 1.711647e-07, 2.958026e-07, 2.482692e-06, 4.277709e-06,
  3.189126e-06, 3.656513e-06, 4.314562e-06, 7.878569e-06, 2.549024e-05, 
    4.898949e-05, 1.668707e-05, 3.013343e-05, 3.132698e-05, 1.508874e-05, 
    3.586172e-06, 4.282727e-07, 6.700711e-08, 8.950472e-07, 3.958863e-07,
  3.421615e-06, 4.504378e-06, 5.561319e-06, 1.621624e-05, 3.369983e-05, 
    4.639975e-05, 6.169933e-05, 2.987337e-05, 3.297358e-05, 2.503394e-05, 
    9.560295e-06, 1.013428e-06, 1.916907e-07, 1.242021e-06, 1.388064e-07,
  5.940767e-06, 5.06184e-06, 7.4186e-06, 2.084322e-05, 3.144327e-05, 
    4.736938e-05, 7.549708e-05, 8.74094e-05, 3.567924e-05, 1.914168e-05, 
    1.409155e-05, 2.182309e-06, 4.285555e-07, 1.911415e-06, 2.153766e-06,
  4.536085e-06, 3.883431e-06, 8.66048e-06, 1.754519e-05, 2.59201e-05, 
    4.882933e-05, 6.966646e-05, 6.261593e-05, 3.626464e-05, 2.218886e-05, 
    1.321459e-05, 2.073848e-06, 5.102925e-07, 7.965907e-07, 1.791912e-06,
  1.192388e-06, 3.564452e-06, 9.639432e-06, 1.623474e-05, 3.250649e-05, 
    4.036534e-05, 4.338711e-05, 4.458096e-05, 3.011992e-05, 1.476266e-05, 
    9.648266e-06, 2.889169e-06, 5.785329e-07, 8.928534e-07, 2.336401e-06,
  1.432983e-06, 4.782587e-06, 1.136311e-05, 2.373198e-05, 3.508971e-05, 
    3.306643e-05, 3.54153e-05, 3.117997e-05, 1.958219e-05, 1.016191e-05, 
    8.019207e-06, 2.931979e-06, 1.399179e-06, 3.096168e-06, 3.988133e-06,
  2.262047e-06, 5.272163e-06, 1.782321e-05, 3.132492e-05, 2.718845e-05, 
    2.433518e-05, 3.066314e-05, 2.989906e-05, 1.97521e-05, 8.996923e-06, 
    2.709129e-06, 2.213173e-06, 2.213236e-06, 2.26789e-06, 8.466697e-06,
  3.955232e-06, 1.286214e-05, 2.569641e-05, 2.970359e-05, 1.551822e-05, 
    1.776408e-05, 2.413248e-05, 2.524105e-05, 1.477588e-05, 4.193634e-06, 
    2.421665e-06, 2.968536e-06, 2.95919e-06, 2.031678e-06, 7.447518e-06,
  6.461377e-05, 6.507822e-05, 5.986479e-05, 5.402783e-05, 5.923898e-05, 
    7.78544e-05, 8.169987e-05, 7.956062e-05, 9.130304e-05, 8.39505e-05, 
    6.52397e-05, 4.943591e-05, 3.067562e-05, 9.44105e-06, 2.401593e-06,
  6.417975e-05, 2.838288e-05, 3.64703e-05, 4.607282e-05, 4.977719e-05, 
    5.512065e-05, 5.717625e-05, 5.027973e-05, 4.748543e-05, 4.472793e-05, 
    3.959297e-05, 4.082702e-05, 3.010405e-05, 1.767065e-05, 4.290698e-06,
  2.080155e-05, 1.996842e-05, 2.600208e-05, 3.275987e-05, 2.975375e-05, 
    1.682398e-05, 1.608102e-05, 3.28491e-05, 3.203885e-05, 2.561113e-05, 
    2.608112e-05, 3.18099e-05, 3.223883e-05, 1.796887e-05, 5.078018e-06,
  1.431001e-05, 1.810461e-05, 2.21465e-05, 1.681119e-05, 1.691286e-05, 
    1.393882e-05, 1.625338e-05, 6.685225e-06, 6.051623e-06, 2.285291e-05, 
    2.432314e-05, 3.395477e-05, 3.342493e-05, 1.672774e-05, 5.451942e-06,
  1.19985e-05, 1.25202e-05, 1.231426e-05, 7.662401e-06, 1.115774e-05, 
    2.306164e-05, 1.939345e-05, 1.745769e-05, 1.962989e-05, 1.309996e-05, 
    2.799822e-05, 3.817716e-05, 2.930619e-05, 1.189763e-05, 5.138241e-06,
  8.602404e-06, 7.569498e-06, 7.725691e-06, 6.356518e-06, 1.039707e-05, 
    1.316196e-05, 9.195706e-06, 9.53128e-06, 6.596741e-06, 6.205194e-06, 
    1.475851e-05, 2.616756e-05, 1.801352e-05, 8.004384e-06, 2.844504e-06,
  8.602453e-06, 7.850917e-06, 8.701125e-06, 8.911398e-06, 9.183531e-06, 
    4.35107e-06, 1.508443e-06, 4.442307e-06, 2.108636e-06, 6.207292e-07, 
    5.636314e-06, 9.130522e-06, 7.912977e-06, 5.510292e-06, 2.526419e-06,
  1.551147e-05, 1.147526e-05, 9.422093e-06, 7.659754e-06, 4.935473e-06, 
    5.208264e-06, 4.853966e-06, 5.614264e-06, 4.293328e-06, 1.399319e-06, 
    1.031833e-06, 2.490117e-06, 3.18157e-06, 3.472348e-06, 5.307211e-06,
  1.649235e-05, 9.016857e-06, 6.444661e-06, 4.607419e-06, 3.89109e-06, 
    4.377793e-06, 5.886901e-06, 7.247306e-06, 5.786321e-06, 4.678986e-06, 
    2.167106e-06, 1.601072e-06, 1.682475e-06, 2.816206e-06, 8.796897e-06,
  1.28925e-05, 8.043104e-06, 5.117885e-06, 3.741282e-06, 2.963866e-06, 
    3.137131e-06, 3.730607e-06, 5.464627e-06, 6.250188e-06, 2.74299e-06, 
    1.726156e-06, 1.451052e-06, 1.559048e-06, 3.297399e-06, 5.020292e-06,
  3.359725e-06, 6.03348e-06, 4.303819e-06, 2.324897e-06, 1.877393e-06, 
    2.273445e-06, 1.733497e-06, 2.760112e-06, 6.894362e-06, 1.721251e-05, 
    3.363118e-05, 5.572694e-05, 6.968444e-05, 5.985574e-05, 3.298965e-05,
  6.269426e-06, 5.953673e-06, 3.567141e-06, 3.205713e-06, 3.87944e-07, 
    6.184524e-07, 4.938087e-07, 1.706442e-06, 3.178325e-06, 6.164846e-06, 
    6.391213e-06, 2.096638e-05, 5.59963e-05, 6.087698e-05, 3.850452e-05,
  9.065649e-06, 1.111895e-05, 8.463851e-06, 1.475339e-06, 1.392365e-07, 
    1.356421e-06, 1.495328e-07, 1.165369e-06, 2.876144e-06, 7.954432e-06, 
    1.224587e-05, 1.298626e-05, 3.321913e-05, 6.280216e-05, 5.219805e-05,
  1.173317e-05, 1.175566e-05, 1.100042e-05, 5.118707e-06, 5.06315e-07, 
    3.477321e-07, 1.813039e-06, 1.245782e-07, 7.889429e-07, 8.33144e-06, 
    2.177875e-05, 3.236045e-05, 5.693999e-05, 7.879869e-05, 5.59507e-05,
  1.464674e-05, 1.238633e-05, 1.214291e-05, 7.160526e-06, 5.906104e-06, 
    5.965382e-06, 2.129646e-06, 5.020975e-06, 1.789345e-05, 1.041693e-05, 
    2.300761e-05, 3.717156e-05, 6.320227e-05, 6.656095e-05, 3.978308e-05,
  1.82848e-05, 1.203602e-05, 1.060639e-05, 8.487829e-06, 8.21758e-06, 
    6.613093e-06, 8.592815e-06, 8.112135e-06, 9.654927e-06, 6.554472e-06, 
    5.792043e-06, 1.707795e-05, 3.441784e-05, 3.448162e-05, 1.44177e-05,
  2.144331e-05, 1.282136e-05, 1.021438e-05, 9.254536e-06, 6.164056e-06, 
    6.230129e-06, 6.350104e-06, 8.05849e-06, 9.578451e-06, 3.372919e-06, 
    2.310569e-06, 7.019619e-06, 9.986312e-06, 9.721003e-06, 3.733622e-06,
  2.006228e-05, 1.214473e-05, 9.479532e-06, 7.323357e-06, 5.310974e-06, 
    7.037753e-06, 6.775839e-06, 7.315845e-06, 7.481306e-06, 2.933258e-06, 
    1.937417e-06, 3.005122e-06, 5.410015e-06, 5.495407e-06, 6.340781e-06,
  1.558215e-05, 1.144097e-05, 7.398492e-06, 5.335171e-06, 6.035847e-06, 
    6.778323e-06, 7.170054e-06, 9.161747e-06, 8.694434e-06, 6.543021e-06, 
    3.652082e-06, 2.354643e-06, 2.290107e-06, 2.292288e-06, 1.950452e-06,
  7.788136e-06, 8.656011e-06, 5.568119e-06, 4.62207e-06, 5.583302e-06, 
    6.06863e-06, 7.872999e-06, 1.208101e-05, 1.089694e-05, 3.422396e-06, 
    1.502841e-06, 1.160206e-06, 3.287708e-06, 1.901703e-06, 6.451165e-07,
  2.845214e-06, 5.396534e-06, 1.182744e-05, 1.489051e-05, 1.182591e-05, 
    6.380966e-06, 1.685761e-06, 1.418815e-07, 2.515129e-08, 6.231208e-06, 
    7.566636e-06, 4.726092e-06, 8.309521e-06, 5.814773e-06, 7.722375e-06,
  7.493979e-06, 4.923939e-06, 8.529282e-06, 1.007786e-05, 5.451554e-06, 
    2.708955e-06, 1.310354e-06, 1.139693e-06, 7.068342e-07, 1.77273e-06, 
    7.5666e-06, 7.090767e-06, 6.949012e-06, 1.405779e-05, 8.521966e-06,
  1.154778e-05, 1.51161e-05, 1.316927e-05, 8.123363e-06, 4.62918e-06, 
    7.193065e-06, 6.797027e-07, 3.443915e-06, 2.567739e-06, 4.539624e-06, 
    1.181261e-05, 1.470166e-05, 1.643124e-05, 1.324899e-05, 1.18981e-05,
  1.141203e-05, 2.03815e-05, 2.20015e-05, 8.394721e-06, 6.42352e-06, 
    4.948467e-06, 7.182133e-06, 1.374579e-06, 1.027474e-06, 4.633133e-06, 
    1.558213e-05, 2.54884e-05, 2.815473e-05, 2.215511e-05, 2.443428e-05,
  1.756067e-05, 1.807823e-05, 2.287497e-05, 1.179774e-05, 8.070798e-06, 
    8.225065e-06, 6.4192e-06, 8.882375e-06, 1.381452e-05, 7.287821e-06, 
    1.714361e-05, 3.233731e-05, 4.297637e-05, 4.162932e-05, 3.981017e-05,
  2.14276e-05, 2.287844e-05, 1.977942e-05, 1.505577e-05, 8.04585e-06, 
    8.874482e-06, 9.081114e-06, 4.928652e-06, 6.43767e-06, 1.076298e-05, 
    1.491195e-05, 2.751815e-05, 4.075731e-05, 4.945203e-05, 4.599309e-05,
  1.87864e-05, 1.914364e-05, 1.951267e-05, 1.264083e-05, 7.711642e-06, 
    8.659074e-06, 7.095453e-06, 6.069449e-06, 3.489412e-06, 4.612597e-06, 
    1.047411e-05, 2.019438e-05, 3.119526e-05, 3.620093e-05, 3.144771e-05,
  1.919834e-05, 1.925062e-05, 1.561718e-05, 1.04055e-05, 9.018997e-06, 
    8.798526e-06, 6.040141e-06, 3.940791e-06, 2.323787e-06, 4.173093e-06, 
    4.432208e-06, 9.502231e-06, 1.547135e-05, 1.90258e-05, 1.837428e-05,
  2.011809e-05, 1.865637e-05, 9.398602e-06, 7.82988e-06, 6.203267e-06, 
    6.613338e-06, 6.818678e-06, 8.016848e-06, 5.113476e-06, 5.978412e-06, 
    7.21035e-06, 6.778709e-06, 6.821499e-06, 1.452486e-05, 2.070841e-05,
  1.273336e-05, 1.072904e-05, 2.702808e-06, 4.456861e-06, 4.378082e-06, 
    7.166221e-06, 3.651907e-06, 1.132792e-05, 9.766618e-06, 4.985898e-06, 
    3.790623e-06, 3.759085e-06, 5.019163e-06, 7.89492e-06, 1.91533e-05,
  9.389407e-06, 4.923389e-06, 2.33367e-06, 4.257169e-06, 3.288059e-06, 
    3.417835e-06, 2.553482e-07, 3.314005e-07, 5.075444e-07, 3.560409e-06, 
    3.170666e-06, 1.799695e-06, 9.516944e-06, 3.764661e-05, 6.742976e-05,
  1.903616e-05, 4.682043e-06, 7.517605e-07, 3.709709e-06, 2.831196e-06, 
    1.754399e-06, 4.620528e-07, 1.246545e-06, 1.51343e-06, 1.349563e-06, 
    2.493294e-06, 5.077207e-06, 5.165042e-06, 1.661293e-05, 3.600595e-05,
  2.742939e-05, 4.106066e-06, 5.212498e-06, 2.359099e-06, 1.445039e-06, 
    5.325367e-06, 4.127486e-07, 5.768156e-06, 9.148152e-06, 3.978858e-06, 
    1.47957e-06, 6.947022e-06, 6.237659e-06, 8.77788e-06, 1.555931e-05,
  1.842362e-05, 4.711033e-06, 8.872401e-06, 6.503246e-06, 2.246325e-06, 
    7.116068e-07, 3.352368e-06, 2.419495e-06, 5.429523e-06, 1.107076e-05, 
    4.448295e-06, 6.391241e-06, 4.816054e-06, 3.907436e-06, 5.488695e-06,
  8.549784e-06, 6.228712e-06, 9.792414e-06, 7.274047e-06, 4.503674e-06, 
    3.079495e-06, 6.503979e-07, 6.919499e-06, 1.545094e-05, 1.870832e-05, 
    1.845104e-05, 8.897237e-06, 5.334015e-06, 5.608882e-06, 4.389419e-06,
  6.928535e-06, 6.734562e-06, 8.793344e-06, 7.602413e-06, 7.374924e-06, 
    5.326502e-06, 2.846697e-06, 4.340938e-06, 1.423411e-05, 2.739145e-05, 
    3.411393e-05, 2.248124e-05, 8.959225e-06, 2.819704e-06, 4.275845e-06,
  8.584811e-06, 8.952844e-06, 6.862953e-06, 6.645283e-06, 6.480727e-06, 
    5.409923e-06, 3.935086e-06, 4.481546e-06, 7.502397e-06, 1.95835e-05, 
    4.067889e-05, 4.866456e-05, 2.453122e-05, 1.034355e-05, 4.316948e-06,
  8.286435e-06, 1.043514e-05, 6.112895e-06, 6.029956e-06, 6.459568e-06, 
    5.812283e-06, 4.058685e-06, 4.127491e-06, 6.032338e-06, 1.231752e-05, 
    3.431906e-05, 5.859361e-05, 5.80564e-05, 2.705385e-05, 1.146482e-05,
  1.358285e-05, 5.995799e-06, 4.934856e-06, 4.691866e-06, 4.963572e-06, 
    6.269283e-06, 5.489763e-06, 6.080716e-06, 6.405039e-06, 1.056082e-05, 
    2.339522e-05, 5.37753e-05, 6.96634e-05, 5.706725e-05, 2.392282e-05,
  9.629186e-06, 4.804518e-06, 4.166627e-07, 5.699289e-06, 6.934064e-06, 
    6.763335e-06, 7.090568e-06, 1.041666e-05, 1.050823e-05, 9.015092e-06, 
    1.422628e-05, 3.322393e-05, 5.854638e-05, 6.618677e-05, 5.102866e-05,
  2.838961e-05, 4.293687e-05, 1.286352e-05, 1.923257e-07, 6.803951e-07, 
    4.265347e-07, 1.831827e-06, 3.788339e-06, 4.46395e-06, 2.998645e-06, 
    5.219167e-06, 5.09348e-06, 4.574867e-06, 2.367142e-05, 3.462048e-05,
  5.276811e-05, 4.2183e-05, 1.612191e-06, 1.562236e-08, 6.942684e-07, 
    2.055875e-07, 1.933013e-06, 4.497392e-06, 5.154453e-06, 1.362628e-06, 
    4.492301e-06, 5.068258e-06, 1.199078e-06, 9.91334e-06, 1.323074e-05,
  3.302747e-05, 8.940449e-06, 3.224037e-06, 1.143672e-06, 5.992043e-07, 
    2.544583e-06, 2.518903e-06, 2.019903e-05, 2.855547e-05, 1.228235e-05, 
    2.911834e-06, 4.834078e-06, 2.18011e-06, 1.621031e-06, 6.9292e-06,
  1.465577e-05, 8.114616e-06, 7.788531e-06, 5.097275e-06, 4.404361e-06, 
    9.917136e-07, 7.774606e-06, 1.228641e-05, 2.142596e-05, 2.506648e-05, 
    7.757378e-06, 6.512585e-06, 4.000954e-06, 3.504094e-07, 4.045992e-06,
  1.33218e-05, 1.086862e-05, 1.085247e-05, 6.340147e-06, 5.743324e-06, 
    8.077638e-06, 5.424725e-06, 1.576309e-05, 2.777896e-05, 2.954742e-05, 
    2.444868e-05, 8.265697e-06, 5.024435e-06, 6.606811e-07, 9.088951e-07,
  1.484656e-05, 9.999098e-06, 1.040249e-05, 8.48972e-06, 6.4598e-06, 
    7.052226e-06, 8.763221e-06, 1.432985e-05, 3.580184e-05, 5.419345e-05, 
    3.362312e-05, 9.54183e-06, 5.752278e-06, 2.711237e-06, 3.152865e-07,
  1.536469e-05, 1.150616e-05, 1.019974e-05, 8.377626e-06, 6.411725e-06, 
    8.383535e-06, 6.740983e-06, 8.230184e-06, 1.933781e-05, 3.111472e-05, 
    3.120402e-05, 1.597647e-05, 5.565149e-06, 5.318601e-06, 2.804229e-07,
  1.766537e-05, 1.277791e-05, 7.092728e-06, 7.165505e-06, 6.945709e-06, 
    7.831264e-06, 3.268345e-06, 2.962955e-06, 5.264912e-06, 1.278364e-05, 
    2.304449e-05, 1.729121e-05, 5.796038e-06, 2.614139e-06, 2.357514e-06,
  1.386916e-05, 8.690902e-06, 3.909901e-06, 6.233429e-06, 6.612791e-06, 
    1.767547e-06, 2.220731e-06, 5.502704e-06, 4.323792e-06, 8.566977e-06, 
    1.244704e-05, 1.878849e-05, 8.908642e-06, 2.703116e-06, 5.614037e-06,
  9.952251e-06, 7.690353e-06, 5.604056e-07, 5.931749e-06, 5.349448e-06, 
    5.528561e-07, 2.281944e-06, 6.77284e-06, 7.883456e-06, 3.596257e-06, 
    5.285882e-06, 1.168526e-05, 1.365869e-05, 8.34545e-06, 2.739745e-06,
  3.989811e-05, 2.413897e-05, 3.638578e-06, 1.412971e-07, 3.915336e-07, 
    6.779588e-07, 1.341254e-06, 1.513547e-06, 4.188093e-06, 1.050763e-05, 
    1.168858e-05, 5.694007e-06, 6.355109e-06, 7.173945e-06, 2.029438e-05,
  1.743335e-05, 8.551776e-06, 4.894281e-07, 6.508861e-07, 4.315931e-07, 
    2.564081e-07, 2.220632e-06, 2.979275e-06, 3.712224e-06, 5.289214e-06, 
    8.760476e-06, 7.598447e-06, 6.856458e-06, 6.52363e-06, 1.438404e-05,
  1.107205e-05, 1.115702e-05, 7.580691e-06, 1.912974e-06, 8.936844e-07, 
    3.027986e-06, 1.814738e-06, 1.071057e-05, 1.672846e-05, 1.359904e-05, 
    4.139702e-06, 5.128421e-06, 6.173279e-06, 3.129782e-06, 1.982566e-05,
  1.418445e-05, 1.376191e-05, 1.211515e-05, 4.69484e-06, 4.168801e-06, 
    3.490268e-06, 4.156155e-06, 5.271762e-06, 1.080165e-05, 1.153084e-05, 
    6.900013e-06, 6.217233e-06, 6.371837e-06, 2.524052e-06, 2.236203e-05,
  1.395991e-05, 1.29161e-05, 1.132093e-05, 7.142793e-06, 6.916533e-06, 
    5.377354e-06, 1.700053e-06, 1.158965e-05, 2.741596e-05, 1.307032e-05, 
    7.732603e-06, 1.040722e-05, 5.40429e-06, 6.424003e-06, 1.94738e-05,
  1.153432e-05, 1.00639e-05, 9.275299e-06, 8.227691e-06, 6.88167e-06, 
    4.941586e-06, 3.199269e-06, 5.904402e-06, 1.53815e-05, 2.094056e-05, 
    8.361374e-06, 9.122399e-06, 4.763739e-06, 5.732988e-06, 1.502902e-05,
  1.059946e-05, 9.333927e-06, 7.998836e-06, 5.684186e-06, 3.924346e-06, 
    4.906349e-06, 2.466575e-06, 2.240974e-06, 8.411208e-06, 1.114641e-05, 
    8.334076e-06, 5.215964e-06, 2.36861e-06, 5.020339e-06, 1.158219e-05,
  1.018485e-05, 6.658588e-06, 2.952958e-06, 2.154654e-06, 2.107293e-06, 
    5.886133e-06, 3.69111e-06, 1.086924e-06, 2.432814e-06, 4.880168e-06, 
    8.282212e-06, 5.362387e-06, 2.04608e-06, 4.981138e-06, 7.508297e-06,
  8.40073e-06, 8.193314e-06, 1.572888e-06, 1.034046e-06, 1.174002e-07, 
    3.282769e-06, 4.868092e-06, 7.330556e-06, 9.492485e-06, 7.399083e-06, 
    6.501946e-06, 6.270732e-06, 3.435731e-06, 2.527366e-06, 3.679643e-06,
  6.184221e-06, 4.218939e-06, 3.23161e-07, 1.341632e-06, 3.710132e-08, 
    1.931183e-06, 4.236612e-06, 1.11407e-05, 1.582171e-05, 6.908372e-06, 
    1.904617e-06, 5.834456e-06, 4.196407e-06, 1.977476e-06, 2.601492e-06,
  6.056479e-07, 2.13069e-06, 1.743898e-06, 1.623723e-06, 9.577798e-07, 
    1.132442e-06, 5.834523e-07, 3.110098e-06, 4.37123e-06, 8.45628e-06, 
    1.444106e-05, 1.066454e-05, 9.194448e-06, 1.036927e-05, 1.038049e-05,
  7.288066e-07, 9.081153e-07, 2.717202e-06, 3.832453e-06, 1.724363e-06, 
    5.163744e-07, 2.861252e-07, 2.156581e-06, 3.736128e-06, 7.83951e-06, 
    1.148922e-05, 1.038634e-05, 7.142264e-06, 1.380672e-05, 9.95038e-06,
  5.79082e-06, 8.380599e-06, 3.961726e-06, 4.848121e-06, 2.586926e-06, 
    5.379894e-06, 1.814268e-07, 2.282043e-06, 6.965292e-06, 8.364095e-06, 
    1.084264e-05, 9.994698e-06, 6.591789e-06, 7.377065e-06, 1.0306e-05,
  5.834726e-06, 1.02177e-05, 7.104295e-06, 5.410906e-06, 2.895097e-06, 
    1.199247e-06, 3.662365e-06, 7.290485e-07, 4.050084e-06, 8.606365e-06, 
    9.257197e-06, 1.191007e-05, 7.87401e-06, 4.936049e-06, 1.379013e-05,
  6.235086e-06, 8.206705e-06, 7.543603e-06, 7.477081e-06, 4.11795e-06, 
    7.256714e-06, 4.860563e-06, 1.149099e-05, 2.574859e-05, 1.045803e-05, 
    9.264287e-06, 9.072e-06, 8.422388e-06, 5.513799e-06, 1.442384e-05,
  8.136131e-06, 8.379619e-06, 6.21716e-06, 6.556558e-06, 5.108728e-06, 
    6.348198e-06, 6.423345e-06, 5.189011e-06, 6.839606e-06, 9.622095e-06, 
    8.187149e-06, 8.182608e-06, 7.771333e-06, 6.001315e-06, 1.583472e-05,
  9.020778e-06, 7.040358e-06, 2.418379e-06, 1.5075e-06, 5.519734e-06, 
    4.857622e-06, 6.885512e-06, 5.491183e-06, 4.1839e-06, 6.040667e-06, 
    8.361265e-06, 7.722088e-06, 7.352641e-06, 5.840513e-06, 1.239284e-05,
  1.056075e-05, 6.483214e-06, 2.589122e-07, 1.221089e-08, 3.927523e-06, 
    4.443479e-06, 6.89566e-06, 5.415431e-06, 4.619128e-06, 5.821777e-06, 
    7.364273e-06, 6.793421e-06, 5.745113e-06, 8.790387e-06, 1.270546e-05,
  1.00984e-05, 7.050213e-06, 3.247074e-07, 1.901261e-08, 1.323229e-06, 
    4.439068e-06, 3.230183e-06, 7.52968e-06, 1.206934e-05, 9.842935e-06, 
    7.104733e-06, 6.168612e-06, 7.793624e-06, 8.939269e-06, 1.105671e-05,
  7.285989e-06, 3.098031e-06, 2.002163e-07, 1.631011e-08, 1.977538e-06, 
    3.031299e-06, 1.109105e-06, 1.375479e-05, 1.530847e-05, 7.484025e-06, 
    8.941593e-06, 7.562183e-06, 7.559953e-06, 8.445249e-06, 8.70114e-06,
  2.611773e-07, 4.337942e-06, 4.208377e-06, 3.761073e-06, 3.420587e-06, 
    3.441579e-06, 2.771427e-06, 2.111887e-06, 8.020303e-07, 4.468932e-06, 
    8.306841e-06, 1.095987e-05, 1.570445e-05, 1.077637e-05, 1.271455e-05,
  3.698739e-06, 3.098672e-06, 3.782154e-06, 4.79585e-06, 4.257683e-06, 
    2.720651e-06, 2.047976e-06, 2.269103e-07, 3.93218e-07, 4.622375e-06, 
    7.306754e-06, 7.859457e-06, 1.648674e-05, 1.498587e-05, 1.137283e-05,
  5.801015e-06, 6.245021e-06, 3.814876e-06, 5.687535e-06, 4.479904e-06, 
    8.597227e-06, 3.61167e-07, 7.938921e-07, 2.622192e-06, 5.160054e-06, 
    5.881831e-06, 7.135762e-06, 9.404992e-06, 8.470261e-06, 9.900173e-06,
  4.196726e-06, 4.143412e-06, 7.819132e-06, 6.016027e-06, 6.031475e-06, 
    3.021594e-06, 7.449645e-06, 1.732298e-07, 1.020722e-06, 5.154212e-06, 
    7.434706e-06, 5.850917e-06, 9.010485e-06, 7.43258e-06, 9.410864e-06,
  3.742164e-06, 3.869968e-06, 6.211324e-06, 5.952541e-06, 6.554128e-06, 
    7.961448e-06, 5.141805e-06, 7.80449e-06, 1.604802e-05, 5.43488e-06, 
    8.053631e-06, 5.474173e-06, 8.599882e-06, 6.145081e-06, 7.185337e-06,
  4.679287e-06, 4.029462e-06, 4.657964e-06, 6.566689e-06, 4.325641e-06, 
    7.222531e-06, 7.503176e-06, 6.959099e-06, 6.732367e-06, 7.027473e-06, 
    8.380153e-06, 5.64817e-06, 5.447398e-06, 6.705685e-06, 5.579553e-06,
  8.35373e-06, 6.833466e-06, 4.918893e-06, 3.605372e-06, 4.410154e-06, 
    8.320009e-06, 7.291238e-06, 5.901411e-06, 5.807071e-06, 6.453925e-06, 
    6.545053e-06, 4.957339e-06, 6.123102e-06, 3.650779e-06, 6.252352e-06,
  9.46384e-06, 8.022608e-06, 1.785473e-06, 3.404444e-06, 5.111402e-06, 
    3.815979e-06, 6.557791e-06, 4.749054e-06, 3.556216e-06, 6.454394e-06, 
    3.640192e-06, 5.157017e-06, 4.744413e-06, 5.572864e-06, 8.861061e-06,
  6.687053e-06, 4.588681e-06, 8.367055e-07, 4.61829e-06, 6.218947e-06, 
    4.811147e-06, 5.28841e-06, 7.487231e-06, 8.95105e-06, 9.952866e-06, 
    8.176257e-06, 6.493965e-06, 5.119073e-06, 4.340986e-06, 5.971518e-06,
  2.835211e-06, 3.821602e-07, 1.310176e-06, 1.622634e-06, 4.511311e-06, 
    1.509542e-06, 4.347524e-06, 1.006876e-05, 1.247458e-05, 3.668493e-06, 
    6.761957e-06, 6.773733e-06, 8.315877e-06, 5.233764e-06, 6.16075e-06,
  2.095979e-06, 3.067616e-06, 4.874391e-06, 4.581895e-06, 4.768546e-06, 
    5.74298e-06, 5.780656e-06, 1.55817e-06, 2.282394e-07, 6.492478e-06, 
    9.642883e-06, 8.572297e-06, 7.311778e-06, 6.268122e-06, 7.689195e-06,
  1.884853e-06, 1.799058e-06, 4.161214e-06, 4.603378e-06, 5.485687e-06, 
    4.241877e-06, 5.149102e-06, 5.643259e-07, 8.69593e-08, 2.35404e-06, 
    6.779997e-06, 7.682668e-06, 5.645602e-06, 1.001784e-05, 1.511874e-05,
  4.578945e-06, 6.462405e-06, 3.282389e-06, 4.304963e-06, 6.035822e-06, 
    1.249601e-05, 3.871674e-06, 3.907481e-06, 1.130625e-06, 3.803997e-06, 
    5.747557e-06, 4.915524e-06, 4.7435e-06, 6.620992e-06, 1.034022e-05,
  6.652499e-06, 8.914006e-06, 7.015916e-06, 6.299372e-06, 9.344161e-06, 
    1.490736e-05, 1.909305e-05, 5.936425e-06, 3.092047e-06, 2.329433e-06, 
    5.575994e-06, 4.407123e-06, 4.990393e-06, 5.904996e-06, 9.93608e-06,
  1.199119e-05, 1.087057e-05, 1.282865e-05, 1.123883e-05, 1.225617e-05, 
    1.633364e-05, 2.244075e-05, 2.639715e-05, 1.253168e-05, 7.958913e-06, 
    8.494752e-06, 4.401197e-06, 5.165242e-06, 8.296392e-06, 3.761277e-06,
  2.163738e-05, 2.322283e-05, 1.749081e-05, 1.207661e-05, 1.397617e-05, 
    1.701125e-05, 2.309536e-05, 2.140637e-05, 1.334351e-05, 1.182065e-05, 
    7.856927e-06, 6.100754e-06, 4.734115e-06, 5.337135e-06, 4.400919e-06,
  2.735102e-05, 2.520279e-05, 1.821167e-05, 1.153253e-05, 1.695701e-05, 
    1.654068e-05, 1.796387e-05, 2.14131e-05, 2.268322e-05, 1.464193e-05, 
    6.17554e-06, 5.023048e-06, 6.000335e-06, 4.735313e-06, 5.857567e-06,
  2.422906e-05, 2.353912e-05, 1.569389e-05, 1.45913e-05, 1.707527e-05, 
    1.883429e-05, 1.906126e-05, 2.016446e-05, 1.960277e-05, 1.351131e-05, 
    8.141598e-06, 6.591441e-06, 7.015998e-06, 7.522758e-06, 7.467049e-06,
  2.085529e-05, 2.108236e-05, 8.984331e-06, 1.660191e-05, 1.680727e-05, 
    1.792167e-05, 1.928013e-05, 1.859755e-05, 1.064125e-05, 8.687392e-06, 
    4.589583e-06, 7.477478e-06, 7.65428e-06, 8.113688e-06, 6.657326e-06,
  1.721837e-05, 1.016369e-05, 8.952329e-06, 9.471502e-06, 1.12613e-05, 
    1.151969e-05, 1.411113e-05, 1.107e-05, 6.383593e-06, 5.563375e-06, 
    8.938476e-06, 1.105803e-05, 7.595227e-06, 7.015813e-06, 1.017228e-05,
  1.782578e-06, 3.22923e-06, 6.918455e-06, 6.804899e-06, 8.347937e-06, 
    9.176383e-06, 4.155751e-06, 2.951112e-06, 4.689839e-06, 8.074616e-06, 
    7.178495e-06, 6.392584e-06, 6.593618e-06, 6.771851e-06, 6.037263e-06,
  3.215257e-06, 5.725815e-06, 1.065847e-05, 1.301614e-05, 1.77361e-05, 
    1.406376e-05, 1.326245e-05, 1.195667e-05, 6.900247e-06, 4.924406e-06, 
    3.42282e-06, 4.218472e-06, 4.379473e-06, 5.771277e-06, 5.573941e-06,
  1.399526e-05, 1.933587e-05, 2.011687e-05, 2.685711e-05, 3.032076e-05, 
    2.903551e-05, 1.457189e-05, 2.40553e-05, 1.651247e-05, 6.410206e-06, 
    4.530044e-06, 4.219682e-06, 4.929037e-06, 4.007073e-06, 4.549105e-06,
  2.203258e-05, 2.631875e-05, 3.175759e-05, 2.86388e-05, 2.640731e-05, 
    2.479604e-05, 2.707212e-05, 1.199603e-05, 1.383608e-05, 1.257739e-05, 
    1.036582e-05, 6.99467e-06, 5.034933e-06, 5.500086e-06, 4.420331e-06,
  3.372532e-05, 2.374452e-05, 2.673326e-05, 1.659183e-05, 9.951003e-06, 
    9.550849e-06, 1.043408e-05, 2.519083e-05, 1.900613e-05, 1.433172e-05, 
    2.258677e-05, 1.111355e-05, 4.939542e-06, 4.883922e-06, 4.403716e-06,
  2.478356e-05, 2.00882e-05, 1.644239e-05, 1.038278e-05, 8.898221e-06, 
    1.088945e-05, 9.925691e-06, 7.520319e-06, 8.963007e-06, 9.258461e-06, 
    1.014453e-05, 8.676429e-06, 5.957372e-06, 2.675794e-06, 4.491417e-06,
  1.926636e-05, 1.917187e-05, 1.886822e-05, 8.165467e-06, 1.278935e-05, 
    1.452134e-05, 1.420452e-05, 9.85033e-06, 1.177458e-05, 5.927822e-06, 
    5.473451e-06, 1.045551e-05, 6.20706e-06, 5.628861e-07, 3.771422e-06,
  1.870147e-05, 2.218678e-05, 1.40896e-05, 8.274948e-06, 1.339558e-05, 
    1.589059e-05, 1.392011e-05, 1.453043e-05, 1.050091e-05, 4.643707e-06, 
    7.51995e-06, 9.942572e-06, 5.922609e-06, 4.098054e-06, 8.869508e-06,
  1.644109e-05, 1.476475e-05, 1.133932e-05, 5.876432e-06, 1.362282e-05, 
    1.591509e-05, 1.632928e-05, 1.792258e-05, 9.353378e-06, 4.506242e-06, 
    6.540481e-06, 8.380321e-06, 5.453115e-06, 6.010367e-06, 5.963785e-06,
  1.112557e-05, 1.159018e-05, 5.104506e-06, 7.193107e-06, 1.248466e-05, 
    1.642607e-05, 1.721589e-05, 1.790713e-05, 1.820265e-05, 8.182139e-06, 
    3.566142e-06, 1.141517e-05, 8.83361e-06, 6.150678e-06, 7.928998e-06,
  1.113531e-06, 1.029691e-07, 3.108016e-06, 1.897409e-06, 2.159002e-06, 
    2.839541e-06, 2.581419e-06, 3.057695e-06, 4.257372e-06, 7.50464e-06, 
    1.01566e-05, 1.02192e-05, 8.178878e-06, 6.02294e-06, 6.571536e-06,
  1.521334e-06, 8.371508e-07, 2.325548e-06, 1.84644e-06, 3.948257e-06, 
    5.237966e-06, 6.702269e-06, 4.989425e-06, 6.006117e-06, 9.835803e-06, 
    9.008456e-06, 8.456307e-06, 7.223276e-06, 5.353216e-06, 5.237839e-06,
  4.095622e-06, 3.728219e-06, 2.986538e-06, 3.954819e-06, 6.024413e-06, 
    1.435775e-05, 6.235713e-06, 4.19664e-06, 4.875905e-06, 7.704435e-06, 
    1.111856e-05, 9.777211e-06, 5.988908e-06, 3.489962e-06, 3.627544e-06,
  9.832254e-06, 1.293861e-05, 8.624815e-06, 7.881592e-06, 1.331988e-05, 
    1.86185e-05, 2.079032e-05, 6.284899e-06, 1.48224e-06, 5.849969e-06, 
    8.92803e-06, 9.904407e-06, 8.718639e-06, 4.275557e-06, 3.033398e-06,
  2.178335e-05, 1.008813e-05, 1.156358e-05, 8.417145e-06, 1.502638e-05, 
    2.31608e-05, 2.201376e-05, 2.019151e-05, 5.547063e-06, 1.378546e-06, 
    8.810755e-06, 8.739399e-06, 9.309953e-06, 3.948394e-06, 7.489896e-07,
  1.975764e-05, 1.515233e-05, 7.454674e-06, 1.13223e-05, 1.423967e-05, 
    1.882553e-05, 2.665962e-05, 1.46603e-05, 5.277146e-06, 1.327995e-06, 
    3.385115e-06, 9.459944e-06, 1.205812e-05, 1.853093e-06, 6.922648e-07,
  1.792643e-05, 1.59898e-05, 9.812662e-06, 1.120771e-05, 1.062295e-05, 
    1.16221e-05, 1.581112e-05, 1.861501e-05, 1.050499e-05, 6.7088e-07, 
    1.382568e-06, 1.31514e-05, 1.512929e-05, 4.767173e-07, 1.395008e-06,
  2.013841e-05, 2.21958e-05, 1.407341e-05, 1.055352e-05, 1.138855e-05, 
    1.334688e-05, 1.713566e-05, 1.063736e-05, 8.333321e-06, 1.531126e-06, 
    3.490821e-06, 1.265936e-05, 1.326678e-05, 3.75521e-07, 3.496927e-06,
  2.21475e-05, 2.183869e-05, 7.165751e-06, 7.188112e-06, 1.569237e-05, 
    1.194859e-05, 1.176899e-05, 1.409728e-05, 1.153341e-05, 8.197136e-06, 
    5.970841e-06, 1.259525e-05, 9.063008e-06, 4.314562e-07, 6.82112e-06,
  1.894101e-05, 1.562858e-05, 6.498307e-06, 6.224376e-06, 1.343714e-05, 
    1.492066e-05, 1.047722e-05, 1.300403e-05, 1.347983e-05, 9.206179e-06, 
    6.496903e-06, 1.193048e-05, 1.892327e-06, 4.85328e-07, 5.265168e-06,
  1.338008e-05, 1.322545e-05, 1.47536e-05, 1.365724e-05, 1.430145e-05, 
    5.741347e-06, 1.126747e-06, 2.276434e-06, 1.400954e-06, 1.378734e-06, 
    1.256712e-06, 1.556993e-06, 5.624585e-06, 5.090664e-06, 9.993593e-06,
  4.664325e-06, 4.018085e-06, 5.847404e-06, 9.652461e-06, 1.410705e-05, 
    1.326486e-05, 5.814594e-06, 4.912898e-06, 3.288699e-06, 2.685129e-06, 
    1.045434e-06, 8.029342e-07, 9.097098e-07, 5.326046e-06, 8.206428e-06,
  2.515197e-06, 4.940296e-06, 6.293445e-06, 9.243849e-06, 2.302832e-05, 
    4.502611e-05, 1.926744e-05, 1.75374e-05, 7.844334e-06, 5.628972e-06, 
    3.770931e-06, 1.310221e-06, 1.475646e-06, 1.876325e-06, 6.230901e-06,
  1.075402e-05, 9.283735e-06, 8.901518e-06, 6.498615e-06, 1.111579e-05, 
    2.053784e-05, 4.180365e-05, 2.619596e-05, 7.133768e-06, 8.335394e-06, 
    4.546348e-06, 1.642582e-06, 2.760889e-06, 1.668976e-06, 7.007174e-06,
  1.350217e-05, 7.549202e-06, 7.32409e-06, 2.160784e-06, 2.288017e-06, 
    1.252095e-05, 1.749264e-05, 2.820432e-05, 2.095336e-05, 2.7495e-06, 
    7.2868e-06, 1.714735e-06, 2.035854e-06, 2.498359e-06, 1.122495e-06,
  1.683163e-05, 1.454685e-05, 5.683569e-06, 5.295418e-06, 4.214345e-06, 
    1.862306e-06, 1.232847e-05, 8.709054e-06, 7.803201e-06, 3.674023e-06, 
    8.101571e-06, 4.045035e-06, 5.195822e-06, 6.994046e-07, 1.191702e-06,
  2.130992e-05, 1.880686e-05, 8.234084e-06, 4.410213e-06, 7.521577e-06, 
    9.892415e-07, 3.575002e-06, 1.011248e-05, 8.493947e-06, 2.957126e-06, 
    8.584131e-06, 4.713784e-06, 3.905498e-06, 7.184983e-07, 2.800818e-06,
  2.594156e-05, 2.084652e-05, 7.949171e-06, 4.117465e-06, 9.78106e-06, 
    4.241623e-06, 4.288946e-06, 5.524353e-06, 1.450774e-06, 3.113849e-06, 
    8.22205e-06, 4.757394e-06, 1.687705e-06, 2.973543e-06, 9.178653e-06,
  2.994456e-05, 2.574921e-05, 1.030277e-05, 9.29489e-06, 5.910275e-06, 
    1.002e-05, 1.216551e-05, 1.065707e-05, 4.779045e-06, 7.121593e-06, 
    4.790232e-06, 2.601917e-06, 6.130936e-07, 8.676553e-06, 9.026505e-06,
  2.561211e-05, 2.326172e-05, 5.299088e-06, 1.074412e-05, 8.677855e-06, 
    9.844896e-06, 1.181205e-05, 1.313489e-05, 6.024266e-06, 7.44326e-06, 
    4.555445e-06, 4.853513e-06, 4.866965e-07, 7.100963e-06, 7.215333e-06,
  3.167338e-06, 1.231235e-06, 2.935558e-07, 7.732265e-08, 7.340853e-07, 
    3.356865e-06, 5.017556e-06, 4.178977e-06, 3.261609e-06, 4.778559e-06, 
    2.022744e-06, 1.818585e-06, 2.473961e-06, 4.598301e-06, 2.020742e-05,
  1.047694e-06, 3.203615e-07, 7.57004e-08, 1.863919e-07, 5.584192e-06, 
    9.170856e-06, 8.432019e-06, 7.015666e-06, 3.304082e-06, 4.798489e-06, 
    2.82751e-06, 5.326272e-07, 8.717445e-07, 7.697642e-06, 2.603401e-05,
  2.9417e-07, 2.917097e-07, 2.075009e-07, 5.396617e-06, 9.323279e-06, 
    2.310076e-05, 1.240488e-05, 1.673812e-05, 1.000012e-05, 7.010097e-06, 
    2.775061e-06, 7.355273e-07, 1.253131e-06, 6.106121e-06, 2.098424e-05,
  1.08731e-05, 4.698024e-06, 4.478209e-06, 1.442063e-06, 7.1043e-06, 
    2.144379e-05, 2.985759e-05, 2.113099e-05, 1.188741e-05, 8.334438e-06, 
    3.420341e-06, 2.035585e-06, 1.718545e-06, 5.542941e-06, 1.477594e-05,
  1.424782e-05, 1.004057e-05, 1.371094e-05, 7.790535e-06, 2.956083e-06, 
    1.2277e-05, 1.247535e-05, 2.713626e-05, 2.111318e-05, 3.831128e-06, 
    5.221447e-06, 3.518086e-06, 1.894795e-06, 4.305618e-06, 8.801993e-06,
  1.849227e-05, 1.420247e-05, 8.19851e-06, 1.198515e-05, 6.29809e-06, 
    1.274391e-06, 1.055663e-05, 8.844759e-06, 7.445094e-06, 2.318687e-06, 
    4.904097e-06, 6.137117e-06, 4.143594e-06, 4.647893e-06, 7.835031e-06,
  1.876107e-05, 1.407945e-05, 5.750503e-06, 6.813788e-06, 1.321155e-05, 
    1.542098e-06, 4.045587e-06, 7.956153e-06, 8.024434e-06, 2.272338e-06, 
    6.652273e-06, 5.595378e-06, 7.387211e-06, 4.904846e-06, 7.982475e-06,
  2.183854e-05, 1.99401e-05, 5.50461e-06, 5.728175e-06, 9.841597e-06, 
    5.385994e-06, 3.528418e-06, 4.311667e-06, 3.07005e-06, 2.377793e-06, 
    6.136239e-06, 6.323168e-06, 2.954612e-06, 3.313041e-06, 7.894871e-06,
  2.798026e-05, 2.743454e-05, 8.273474e-06, 8.771637e-06, 4.894625e-06, 
    3.96203e-06, 4.938634e-06, 7.947272e-06, 7.534205e-06, 3.370069e-06, 
    8.410346e-06, 7.379105e-06, 1.594463e-06, 4.277339e-06, 7.113137e-06,
  3.022443e-05, 2.690999e-05, 9.369484e-06, 9.860248e-06, 5.533958e-06, 
    6.870958e-06, 1.049187e-05, 1.377318e-05, 8.839231e-06, 4.004863e-06, 
    1.322694e-05, 8.582563e-06, 1.488507e-06, 7.397462e-06, 6.212709e-06,
  2.705026e-06, 5.509025e-07, 5.167341e-07, 3.263452e-06, 2.21005e-06, 
    2.655246e-06, 3.336198e-06, 1.007403e-06, 3.306345e-06, 7.397969e-06, 
    6.833525e-06, 1.657771e-06, 2.648073e-06, 2.790493e-06, 1.337134e-05,
  2.217421e-06, 7.248319e-08, 6.554799e-07, 8.274841e-07, 6.919846e-06, 
    3.135047e-06, 3.367897e-06, 4.979512e-06, 4.940514e-06, 2.252444e-06, 
    5.297505e-06, 1.742022e-06, 1.13315e-06, 1.470647e-05, 3.466002e-05,
  1.020594e-06, 6.130541e-08, 8.123749e-08, 6.578584e-07, 1.246181e-06, 
    2.797118e-05, 3.054624e-06, 7.35909e-06, 3.530355e-06, 2.466744e-06, 
    4.595498e-06, 1.659958e-06, 3.396638e-06, 2.555001e-05, 4.20639e-05,
  7.854394e-07, 3.047339e-06, 1.012519e-05, 8.677314e-06, 5.468737e-06, 
    9.702086e-06, 3.119441e-05, 1.042654e-05, 3.41678e-06, 2.293918e-06, 
    8.789527e-07, 1.039416e-06, 1.427552e-05, 3.043073e-05, 2.813967e-05,
  9.612903e-06, 7.313115e-06, 8.749026e-06, 6.504634e-06, 4.751564e-06, 
    6.633546e-06, 8.340253e-06, 2.484023e-05, 6.669411e-06, 2.285504e-06, 
    2.546715e-06, 7.423231e-06, 3.143702e-05, 2.770609e-05, 1.010619e-05,
  1.456901e-05, 1.255861e-05, 4.216918e-06, 2.779554e-06, 3.996735e-06, 
    4.963079e-06, 9.385041e-06, 4.437075e-06, 5.877404e-06, 3.199579e-06, 
    8.614017e-06, 2.35326e-05, 3.714504e-05, 1.629694e-05, 4.179299e-06,
  1.401956e-05, 1.164742e-05, 4.646233e-06, 1.963739e-06, 5.081511e-06, 
    4.083122e-06, 6.245573e-06, 5.136423e-06, 5.23856e-06, 5.648236e-06, 
    2.179679e-05, 3.522647e-05, 2.858627e-05, 1.241017e-05, 3.893031e-06,
  1.771029e-05, 1.283893e-05, 5.842081e-06, 9.900863e-07, 9.405692e-06, 
    5.1204e-06, 9.029779e-06, 9.67828e-06, 8.319872e-06, 2.030364e-05, 
    3.698111e-05, 3.2961e-05, 2.152696e-05, 1.173722e-05, 5.940464e-06,
  1.981996e-05, 1.450448e-05, 4.332986e-06, 6.567584e-06, 1.076185e-05, 
    9.925618e-06, 1.082913e-05, 1.057583e-05, 1.429966e-05, 2.483502e-05, 
    3.033044e-05, 2.337012e-05, 1.629036e-05, 8.863473e-06, 4.115205e-06,
  1.598857e-05, 1.179625e-05, 5.821536e-06, 7.596353e-06, 7.219906e-06, 
    9.06383e-06, 9.440597e-06, 1.4108e-05, 1.440219e-05, 2.106159e-05, 
    2.274917e-05, 1.449874e-05, 8.004317e-06, 5.697449e-06, 3.120522e-06,
  9.83459e-05, 8.600657e-05, 6.056247e-05, 3.148778e-05, 2.166172e-05, 
    1.29587e-05, 8.394814e-06, 5.575288e-06, 7.284473e-06, 1.196236e-05, 
    8.232824e-06, 8.147053e-06, 1.213531e-05, 1.009125e-05, 6.123435e-06,
  8.887391e-05, 3.467713e-05, 1.065405e-05, 7.17457e-06, 1.904907e-06, 
    3.003553e-06, 4.047192e-06, 7.483589e-06, 1.086461e-05, 1.451018e-05, 
    9.743354e-06, 5.300002e-06, 4.947787e-06, 1.61653e-05, 5.748785e-06,
  1.407395e-05, 1.681872e-06, 2.181979e-07, 7.735151e-07, 1.884857e-06, 
    1.868234e-05, 4.09733e-06, 3.600416e-06, 5.920359e-06, 4.293547e-06, 
    7.639688e-06, 7.060587e-06, 7.494187e-06, 3.602851e-06, 4.136344e-06,
  6.341827e-08, 1.402778e-06, 2.272358e-06, 1.006471e-07, 5.158839e-08, 
    5.343267e-07, 2.011364e-05, 2.399097e-06, 2.090733e-06, 3.460385e-06, 
    2.596579e-06, 1.793696e-06, 1.81578e-06, 1.681128e-06, 4.335522e-06,
  4.66903e-06, 3.734839e-06, 8.434731e-06, 3.558075e-06, 1.760604e-07, 
    3.008622e-06, 7.421188e-06, 2.332532e-05, 8.932428e-06, 1.501242e-06, 
    1.273029e-06, 8.062237e-07, 8.524834e-07, 2.688192e-06, 8.200792e-06,
  6.57438e-06, 9.688406e-06, 3.516534e-06, 3.528587e-06, 4.612958e-06, 
    6.206918e-06, 7.058266e-06, 5.540864e-06, 4.017062e-06, 9.227006e-07, 
    6.222254e-07, 7.796302e-07, 5.217145e-06, 9.982228e-06, 1.120683e-05,
  7.400231e-06, 8.293876e-06, 6.52246e-06, 2.97463e-06, 5.832438e-06, 
    9.00729e-06, 8.350464e-06, 1.425896e-06, 1.442042e-06, 3.874963e-06, 
    5.196844e-06, 9.602774e-06, 1.309053e-05, 1.26223e-05, 1.091024e-05,
  1.057393e-05, 1.059877e-05, 8.606714e-06, 2.295533e-06, 7.039107e-06, 
    5.870631e-06, 3.770297e-06, 4.152185e-06, 4.658227e-06, 1.229055e-05, 
    1.566284e-05, 1.530758e-05, 1.224301e-05, 1.323733e-05, 1.394434e-05,
  1.403623e-05, 9.939935e-06, 4.946573e-06, 1.009161e-05, 1.093905e-05, 
    1.070393e-05, 1.003589e-05, 1.644451e-05, 2.626995e-05, 2.623618e-05, 
    1.888651e-05, 1.272741e-05, 1.189145e-05, 1.164125e-05, 1.240221e-05,
  9.686781e-06, 9.23746e-06, 6.624244e-06, 1.353198e-05, 1.476709e-05, 
    1.66987e-05, 2.241367e-05, 3.082293e-05, 3.159871e-05, 2.261946e-05, 
    1.551885e-05, 1.070955e-05, 1.031375e-05, 1.124889e-05, 1.057466e-05,
  9.587196e-06, 7.552876e-06, 8.060745e-06, 1.563116e-05, 3.096406e-05, 
    1.962835e-05, 1.054713e-05, 7.498156e-06, 9.033e-06, 1.492964e-05, 
    7.848799e-06, 7.153686e-06, 1.063166e-05, 1.05718e-05, 9.599272e-06,
  4.787671e-05, 4.5596e-05, 5.048017e-05, 7.78712e-05, 6.591436e-05, 
    2.93002e-05, 1.158016e-05, 8.017913e-06, 1.140831e-05, 2.368347e-05, 
    1.456639e-05, 5.079435e-06, 7.608837e-06, 1.565873e-05, 9.652244e-06,
  0.0001853494, 0.00016551, 0.0001502272, 0.0001159967, 5.652727e-05, 
    2.914749e-05, 4.248236e-06, 2.485376e-06, 1.627474e-06, 4.768667e-06, 
    7.763819e-06, 7.987446e-06, 7.131525e-06, 5.101707e-06, 7.447324e-06,
  0.0002372157, 0.0001987353, 0.0001318293, 6.254038e-05, 1.667865e-05, 
    1.059621e-05, 1.892553e-05, 7.003916e-07, 7.121612e-07, 1.33557e-06, 
    4.403883e-06, 8.592147e-06, 1.199303e-05, 9.347177e-06, 5.379097e-06,
  0.0001243226, 8.670025e-05, 3.908065e-05, 7.869057e-06, 1.625046e-06, 
    2.079536e-06, 7.328568e-06, 1.868432e-05, 9.860069e-06, 3.649432e-06, 
    6.584254e-06, 6.147208e-06, 1.105916e-05, 6.73159e-06, 4.271153e-06,
  2.90577e-05, 1.064268e-05, 2.239528e-06, 1.163224e-06, 4.35257e-07, 
    4.548715e-06, 1.014712e-05, 5.702609e-06, 7.510783e-06, 5.413701e-06, 
    4.983461e-06, 5.644318e-06, 4.255181e-06, 6.375798e-06, 5.979365e-06,
  2.712655e-06, 2.446426e-06, 8.506669e-07, 1.376108e-06, 3.403319e-06, 
    7.334986e-06, 9.281921e-06, 8.161323e-06, 6.348349e-06, 4.392113e-06, 
    6.185484e-06, 9.632561e-06, 6.703734e-06, 4.92425e-06, 4.696521e-06,
  1.601808e-06, 6.2657e-06, 6.814994e-07, 6.544915e-07, 7.74722e-06, 
    7.873925e-06, 5.020844e-06, 2.353286e-06, 3.670817e-07, 3.316751e-06, 
    3.98971e-06, 6.254033e-06, 5.571103e-06, 6.924374e-06, 7.148537e-06,
  4.063202e-06, 6.151064e-06, 2.297738e-07, 5.765382e-06, 1.065606e-05, 
    5.411837e-06, 5.915958e-07, 2.586339e-07, 3.134697e-06, 5.526545e-06, 
    5.06995e-06, 4.204615e-06, 7.259145e-06, 9.081195e-06, 9.414553e-06,
  5.901187e-06, 8.285924e-06, 4.514608e-06, 1.081144e-05, 8.690403e-06, 
    2.004875e-06, 8.480116e-07, 2.254305e-06, 6.559288e-06, 7.871101e-06, 
    4.699438e-06, 6.875561e-06, 9.454657e-06, 9.669971e-06, 1.058072e-05,
  3.568546e-06, 8.26111e-06, 7.987193e-06, 5.507056e-06, 1.029102e-05, 
    3.660446e-05, 4.707001e-05, 7.075619e-05, 0.0001199011, 0.0001488983, 
    0.0001396842, 0.0001218911, 9.484539e-05, 6.629421e-05, 3.387565e-05,
  9.218155e-06, 1.122503e-05, 8.58357e-06, 1.172148e-05, 5.635448e-05, 
    0.000117571, 0.0001281546, 0.0001654076, 0.0001716862, 0.0001481969, 
    0.0001162965, 0.0001010821, 7.325471e-05, 5.300889e-05, 2.157334e-05,
  7.979922e-06, 1.201097e-05, 3.699036e-05, 0.0001059424, 0.0001739289, 
    0.0002317273, 0.0001870005, 0.000178798, 0.0001394646, 0.0001187425, 
    8.892706e-05, 6.676853e-05, 4.681418e-05, 2.104954e-05, 9.243106e-06,
  1.313164e-05, 4.378114e-05, 0.0001020789, 0.0001571442, 0.0002049163, 
    0.0001436152, 0.0001850918, 0.0001433026, 0.0001022208, 6.103663e-05, 
    3.614201e-05, 2.312106e-05, 1.793017e-05, 1.146345e-05, 4.231832e-06,
  4.409558e-05, 9.722313e-05, 0.0001539169, 0.0001691248, 0.0001517255, 
    9.197403e-05, 3.633395e-05, 3.269333e-05, 3.605777e-05, 9.89392e-06, 
    3.678322e-06, 4.885484e-06, 6.630637e-06, 6.880437e-06, 2.511879e-06,
  0.0001301694, 0.0001481312, 0.000118559, 6.852249e-05, 3.725644e-05, 
    1.692784e-05, 3.445118e-06, 1.218507e-06, 6.219471e-07, 2.355329e-07, 
    5.869523e-07, 2.85412e-07, 5.501387e-06, 7.189607e-06, 3.425575e-06,
  8.625799e-05, 5.453044e-05, 2.686353e-05, 9.263142e-06, 2.068513e-06, 
    3.64856e-07, 7.599544e-08, 1.819801e-07, 2.970512e-06, 3.702066e-06, 
    3.290276e-06, 4.038485e-06, 7.204895e-06, 3.92659e-06, 2.951364e-06,
  2.715626e-05, 1.324635e-05, 4.85328e-06, 4.51887e-07, 1.082575e-07, 
    8.159549e-07, 3.794767e-07, 3.281727e-06, 3.918165e-06, 3.321026e-06, 
    3.285598e-06, 3.331346e-06, 5.760868e-06, 6.059668e-06, 3.821711e-06,
  1.852764e-05, 9.548067e-06, 7.036572e-07, 7.522431e-07, 2.167524e-06, 
    1.645066e-06, 2.102948e-06, 2.974133e-06, 4.606984e-06, 3.831485e-06, 
    3.69954e-06, 3.509846e-06, 4.55956e-06, 5.333847e-06, 3.835213e-06,
  1.516815e-05, 1.071506e-05, 2.989555e-06, 1.76292e-06, 4.043978e-06, 
    4.877214e-06, 4.463232e-06, 5.278631e-06, 6.226782e-06, 5.386793e-06, 
    4.844779e-06, 6.295631e-06, 5.611012e-06, 4.911853e-06, 3.764132e-06,
  1.864037e-07, 8.37636e-08, 1.599357e-07, 5.347224e-07, 2.953401e-06, 
    7.325123e-06, 1.068988e-05, 1.394263e-05, 1.424042e-05, 1.611154e-05, 
    8.798511e-06, 9.111786e-06, 2.437213e-05, 5.014108e-05, 7.534603e-05,
  2.617798e-07, 6.733438e-07, 1.474709e-06, 4.117542e-06, 9.890023e-06, 
    1.667921e-05, 2.531116e-05, 3.204885e-05, 2.937405e-05, 2.834685e-05, 
    2.594483e-05, 1.965735e-05, 2.641913e-05, 6.088919e-05, 7.129172e-05,
  2.798221e-06, 6.449861e-06, 7.264181e-06, 1.078117e-05, 1.81405e-05, 
    5.091878e-05, 5.046092e-05, 8.169937e-05, 6.424828e-05, 4.318147e-05, 
    2.64106e-05, 2.461978e-05, 2.901283e-05, 4.031639e-05, 5.393052e-05,
  1.135992e-05, 1.363341e-05, 1.860282e-05, 2.09661e-05, 3.361756e-05, 
    4.547169e-05, 0.0001173486, 6.715429e-05, 4.630395e-05, 2.932688e-05, 
    1.474123e-05, 1.814204e-05, 3.549201e-05, 5.625163e-05, 5.71764e-05,
  2.531081e-05, 3.406168e-05, 4.213412e-05, 3.773408e-05, 3.358505e-05, 
    4.177201e-05, 2.409408e-05, 2.530681e-05, 3.833271e-05, 1.024245e-05, 
    1.055454e-05, 1.711839e-05, 4.133104e-05, 5.993967e-05, 4.139381e-05,
  2.7548e-05, 3.872777e-05, 3.524408e-05, 2.264243e-05, 1.461882e-05, 
    7.99047e-06, 2.123951e-06, 9.295869e-07, 1.13813e-06, 4.557402e-06, 
    5.468539e-06, 1.521501e-05, 3.136032e-05, 3.207885e-05, 1.698028e-05,
  2.133838e-05, 1.930087e-05, 1.163292e-05, 2.234577e-06, 5.954727e-07, 
    1.102299e-07, 1.137677e-08, 2.403904e-08, 4.303616e-07, 4.587824e-06, 
    1.179572e-05, 1.624703e-05, 1.986742e-05, 1.108106e-05, 5.576657e-06,
  1.72904e-05, 1.15861e-05, 7.684321e-06, 2.703666e-06, 9.712857e-07, 
    2.835212e-08, 3.807921e-08, 4.06495e-07, 4.613568e-07, 3.12106e-06, 
    6.532793e-06, 1.161108e-05, 1.797538e-05, 1.143634e-05, 4.240003e-06,
  1.630093e-05, 7.662548e-06, 7.623943e-06, 8.552048e-06, 7.25488e-06, 
    4.582305e-06, 3.749743e-06, 5.196272e-06, 3.186084e-06, 3.828278e-06, 
    7.149869e-06, 1.037165e-05, 1.054104e-05, 7.119992e-06, 8.427669e-06,
  1.644615e-05, 6.85081e-06, 6.220307e-06, 7.975323e-06, 6.710323e-06, 
    6.573245e-06, 5.468386e-06, 4.064951e-06, 4.132105e-06, 7.01453e-06, 
    9.559807e-06, 8.450765e-06, 7.165743e-06, 8.042894e-06, 7.384329e-06,
  1.138042e-05, 5.56817e-06, 9.122266e-06, 1.259913e-05, 1.587942e-05, 
    1.093583e-05, 3.799849e-06, 2.725312e-06, 4.732253e-06, 6.760184e-06, 
    5.77969e-06, 5.993655e-06, 1.043235e-05, 1.251102e-05, 1.647177e-05,
  5.520193e-05, 4.585877e-05, 4.459174e-05, 4.559851e-05, 3.95675e-05, 
    1.494856e-05, 3.703307e-06, 2.575638e-06, 4.734699e-06, 6.640323e-06, 
    1.075846e-05, 1.641598e-05, 1.639021e-05, 2.196054e-05, 1.450328e-05,
  0.0001203476, 0.0001040955, 9.111509e-05, 8.665041e-05, 4.297456e-05, 
    1.443993e-05, 2.607836e-06, 5.319735e-07, 7.146675e-07, 4.294249e-06, 
    3.06062e-06, 1.119028e-05, 2.020544e-05, 2.567252e-05, 2.217399e-05,
  0.0001187038, 0.0001124142, 0.0001061657, 7.614818e-05, 2.477719e-05, 
    3.708239e-06, 6.569343e-06, 5.044822e-07, 1.005484e-06, 2.198793e-06, 
    1.584113e-06, 3.657867e-06, 1.013808e-05, 2.760497e-05, 2.723501e-05,
  0.0001274411, 0.0001006393, 6.049286e-05, 2.393078e-05, 5.639853e-06, 
    1.174086e-06, 3.488727e-06, 9.113613e-06, 2.408612e-05, 1.665473e-06, 
    4.380242e-06, 3.148002e-06, 1.422245e-05, 3.808331e-05, 2.867619e-05,
  5.028414e-05, 3.299211e-05, 1.547025e-05, 4.212407e-06, 9.473141e-07, 
    1.380151e-07, 1.735811e-06, 1.490275e-06, 3.240406e-06, 9.327697e-07, 
    2.860622e-06, 6.083909e-06, 4.6213e-05, 6.620164e-05, 3.849351e-05,
  1.159275e-05, 1.203413e-05, 8.346166e-06, 1.36876e-06, 1.470639e-07, 
    2.092012e-07, 2.201945e-07, 1.949113e-06, 2.965999e-06, 2.670553e-07, 
    1.07682e-06, 1.575524e-05, 8.036332e-05, 9.124381e-05, 5.506205e-05,
  1.273245e-05, 1.302441e-05, 7.2412e-06, 5.77144e-06, 4.905639e-06, 
    5.171725e-06, 9.495715e-07, 5.518639e-08, 6.09943e-07, 9.772101e-08, 
    5.497273e-06, 2.737289e-05, 8.357732e-05, 7.688565e-05, 3.494373e-05,
  1.206407e-05, 7.354665e-06, 5.443977e-06, 6.80084e-06, 6.856766e-06, 
    7.747631e-06, 1.463869e-06, 2.625012e-08, 1.09243e-08, 1.58931e-07, 
    4.910929e-06, 3.451258e-05, 5.872103e-05, 3.839674e-05, 1.211809e-05,
  5.882516e-06, 7.849143e-06, 6.485119e-06, 4.28168e-06, 6.507201e-06, 
    7.287822e-06, 6.516727e-06, 1.709023e-07, 2.2631e-07, 1.062591e-06, 
    8.218265e-06, 2.693375e-05, 3.365298e-05, 1.583197e-05, 8.364146e-06,
  3.165079e-06, 9.103375e-07, 1.778623e-06, 6.165657e-06, 1.296933e-05, 
    3.068023e-05, 5.340554e-05, 6.11197e-05, 6.574106e-05, 7.411036e-05, 
    7.790417e-05, 4.300072e-05, 7.438287e-06, 2.588432e-06, 2.573285e-06,
  1.555576e-06, 2.78019e-06, 4.934564e-06, 8.203964e-06, 3.371295e-05, 
    9.2473e-05, 9.031992e-05, 9.827138e-05, 0.0001055145, 0.0001079094, 
    7.776615e-05, 2.372867e-05, 1.878905e-06, 3.561999e-06, 3.598973e-06,
  8.654672e-06, 8.653822e-06, 7.228685e-06, 1.018748e-05, 7.341924e-05, 
    0.0001445106, 0.0001562903, 0.000160857, 0.0001596773, 0.0001164821, 
    5.0183e-05, 9.221146e-06, 9.728079e-07, 1.754583e-06, 5.441277e-06,
  1.431254e-05, 1.86754e-05, 2.723506e-05, 6.879943e-05, 0.0001357163, 
    0.0001210498, 0.0001803959, 0.0001454892, 0.0001158177, 6.750024e-05, 
    2.117848e-05, 3.731695e-06, 5.253112e-07, 1.668527e-06, 9.807277e-06,
  1.71817e-05, 3.765064e-05, 6.054178e-05, 7.858438e-05, 9.91546e-05, 
    0.0001133616, 6.728398e-05, 4.625862e-05, 4.578352e-05, 1.969e-05, 
    5.342338e-06, 6.035143e-07, 9.437338e-07, 9.976063e-06, 1.831993e-05,
  9.253498e-06, 1.594937e-05, 2.170591e-05, 1.6259e-05, 1.323536e-05, 
    2.004354e-05, 2.745365e-05, 2.102762e-05, 1.24109e-05, 7.710801e-06, 
    2.245131e-06, 1.254019e-06, 1.037574e-05, 3.387492e-05, 1.298145e-05,
  5.6515e-06, 9.607707e-06, 8.662123e-06, 3.029857e-06, 4.383302e-06, 
    4.376709e-06, 6.423893e-06, 6.916751e-06, 7.637287e-06, 2.375422e-06, 
    3.671796e-07, 4.668406e-06, 1.985412e-05, 4.19953e-05, 1.60545e-05,
  8.972059e-06, 8.867404e-06, 7.674685e-06, 6.392791e-06, 7.738647e-06, 
    7.191852e-06, 3.547688e-06, 1.364822e-07, 2.132106e-06, 2.088547e-07, 
    1.922016e-06, 7.29585e-06, 1.817667e-05, 3.060889e-05, 2.239872e-05,
  8.895318e-06, 7.689549e-06, 5.746804e-06, 6.300641e-06, 5.003569e-06, 
    3.057291e-06, 2.510306e-06, 8.021405e-09, 4.841145e-09, 6.602769e-07, 
    1.75323e-06, 1.089565e-05, 1.782961e-05, 1.59243e-05, 7.311705e-06,
  5.766032e-06, 4.245308e-06, 4.929521e-06, 8.834838e-06, 8.029647e-06, 
    3.854436e-07, 1.687786e-08, 9.082076e-09, 2.276306e-08, 2.474569e-06, 
    1.372589e-05, 2.143398e-05, 1.276969e-05, 8.5473e-06, 7.510165e-06,
  2.903832e-09, 1.121875e-08, 4.457436e-07, 2.067718e-06, 1.121298e-06, 
    2.192375e-06, 1.602448e-05, 1.655637e-05, 1.842863e-05, 2.113633e-05, 
    2.852695e-05, 8.767148e-05, 0.0001302964, 7.704629e-05, 3.321464e-05,
  1.166713e-08, 5.975383e-07, 2.124015e-06, 2.098652e-06, 2.203652e-06, 
    2.418948e-06, 9.62842e-06, 2.129607e-05, 3.012862e-05, 4.042138e-05, 
    7.555514e-05, 0.0001180948, 7.448291e-05, 2.064769e-05, 3.442895e-06,
  2.977203e-07, 5.391788e-06, 5.220139e-06, 2.035558e-06, 2.435185e-06, 
    9.052002e-06, 8.160486e-06, 3.758724e-05, 6.115388e-05, 8.499435e-05, 
    9.217262e-05, 6.04741e-05, 1.544273e-05, 1.320418e-06, 6.449993e-07,
  2.895787e-06, 7.217696e-06, 1.655169e-06, 4.277527e-06, 3.913024e-06, 
    3.550397e-06, 1.530105e-05, 2.543669e-05, 4.222675e-05, 5.877756e-05, 
    3.86987e-05, 1.551658e-05, 2.463847e-06, 1.535141e-06, 2.674687e-06,
  3.193757e-06, 1.468341e-06, 4.777386e-07, 4.856572e-06, 5.122322e-06, 
    5.362076e-06, 1.005824e-05, 2.02166e-05, 4.011705e-05, 3.041985e-05, 
    2.081619e-05, 8.720947e-06, 5.800341e-06, 4.419519e-06, 3.834399e-06,
  5.060083e-07, 3.929165e-07, 2.143159e-06, 4.052242e-06, 5.539242e-06, 
    6.741428e-06, 5.270555e-06, 1.367423e-05, 1.511672e-05, 1.828346e-05, 
    1.273983e-05, 6.910584e-06, 5.398105e-06, 2.827742e-06, 2.269231e-06,
  1.203553e-06, 4.877533e-06, 2.902673e-06, 4.291666e-06, 6.104857e-06, 
    5.26042e-06, 3.011865e-06, 6.068834e-06, 9.612725e-06, 9.377946e-06, 
    7.647634e-06, 5.643575e-06, 5.841728e-06, 3.655308e-06, 3.076326e-06,
  5.624937e-06, 1.130001e-05, 4.766551e-06, 8.482755e-06, 1.079171e-05, 
    7.256165e-06, 4.626218e-06, 1.332008e-06, 3.473209e-06, 5.515866e-06, 
    6.249429e-06, 4.023552e-06, 5.001848e-06, 4.047665e-06, 3.335817e-06,
  1.081226e-05, 7.262755e-06, 6.467155e-06, 8.285076e-06, 1.00601e-05, 
    5.872705e-06, 4.489558e-06, 2.947012e-07, 2.031667e-06, 6.23752e-06, 
    2.513091e-06, 2.585014e-06, 3.001436e-06, 1.965459e-06, 1.857058e-06,
  5.916047e-06, 3.533484e-06, 6.569253e-06, 1.109222e-05, 1.255683e-05, 
    7.930379e-06, 2.795286e-06, 6.694068e-08, 3.910816e-06, 5.728592e-06, 
    3.289668e-06, 8.888681e-07, 2.678575e-06, 2.658744e-06, 4.428422e-06,
  2.974041e-08, 3.68083e-08, 3.172809e-08, 9.861672e-08, 7.094177e-08, 
    1.776991e-09, 2.864215e-10, 3.234124e-08, 2.536833e-06, 9.624742e-06, 
    1.278282e-05, 6.134519e-06, 7.427691e-06, 6.724117e-06, 1.238212e-05,
  4.050195e-08, 3.280584e-08, 5.449377e-08, 2.968503e-07, 1.182564e-08, 
    7.598291e-10, 2.912559e-08, 1.901451e-07, 2.98879e-06, 9.879538e-06, 
    1.307344e-05, 7.545135e-06, 3.745638e-06, 1.469295e-05, 1.022714e-05,
  3.549271e-08, 2.382785e-06, 3.015217e-07, 2.929257e-08, 1.505426e-09, 
    1.322888e-07, 1.128732e-07, 6.301052e-07, 4.352828e-06, 1.442227e-05, 
    1.178161e-05, 7.877818e-06, 5.108652e-06, 3.65082e-06, 3.057509e-06,
  4.985417e-06, 2.771944e-07, 6.474336e-07, 5.387228e-07, 9.724633e-09, 
    3.723113e-08, 5.019743e-06, 7.631716e-07, 4.464975e-06, 1.382377e-05, 
    6.86362e-06, 8.742765e-06, 6.769612e-06, 2.182856e-06, 2.240045e-06,
  7.859078e-07, 2.149204e-07, 3.194183e-06, 1.144916e-06, 2.156149e-07, 
    1.140732e-06, 3.580804e-06, 9.803568e-06, 2.183076e-05, 1.236075e-05, 
    7.757168e-06, 6.694402e-06, 6.92234e-06, 4.160401e-06, 3.02334e-06,
  1.331102e-08, 6.866301e-07, 1.628712e-06, 5.103627e-06, 2.755854e-06, 
    4.572013e-06, 5.638502e-06, 7.382097e-06, 8.342445e-06, 1.272821e-05, 
    8.938806e-06, 7.632112e-06, 7.754479e-06, 6.922778e-06, 6.510779e-06,
  1.217519e-06, 1.339245e-06, 3.457626e-07, 4.4546e-06, 1.635169e-05, 
    1.629727e-05, 1.070615e-05, 6.838774e-06, 8.943667e-06, 1.121253e-05, 
    7.422752e-06, 5.528997e-06, 7.319448e-06, 9.26195e-06, 1.072221e-05,
  1.780451e-06, 2.458364e-06, 1.359701e-06, 1.437906e-06, 6.503934e-06, 
    1.200413e-05, 7.429603e-06, 2.36396e-06, 7.798483e-06, 9.185358e-06, 
    7.518042e-06, 5.506055e-06, 6.916037e-06, 8.910984e-06, 8.143639e-06,
  3.479413e-06, 5.038539e-06, 1.129347e-06, 1.113914e-06, 5.091847e-06, 
    7.018498e-06, 5.721068e-06, 7.043824e-07, 6.714306e-06, 8.573896e-06, 
    5.654773e-06, 5.668511e-06, 6.675195e-06, 8.856972e-06, 7.095488e-06,
  2.463273e-06, 3.524227e-06, 4.823236e-06, 1.581984e-06, 2.119675e-06, 
    1.009754e-05, 3.856446e-06, 1.611738e-06, 7.42797e-06, 6.395091e-06, 
    5.67213e-06, 6.344477e-06, 6.226019e-06, 8.091512e-06, 7.492257e-06,
  7.119082e-05, 8.905376e-06, 5.920327e-07, 8.754702e-08, 4.367596e-08, 
    3.857017e-09, 2.683423e-08, 1.001368e-08, 1.467445e-07, 6.129695e-06, 
    1.057695e-05, 1.439145e-05, 1.225828e-05, 5.3303e-06, 6.55154e-06,
  3.054627e-05, 2.725055e-06, 2.278875e-07, 3.384017e-08, 4.984615e-09, 
    2.213951e-09, 9.588241e-09, 9.715385e-08, 2.722456e-07, 7.264602e-06, 
    1.17639e-05, 1.754185e-05, 1.214942e-05, 1.159219e-05, 9.251931e-06,
  6.854327e-06, 7.924968e-07, 4.896701e-08, 7.084199e-09, 6.640707e-09, 
    1.896333e-07, 1.684528e-07, 1.27012e-06, 1.708495e-06, 7.628061e-06, 
    1.025227e-05, 1.850894e-05, 1.168471e-05, 9.991859e-06, 1.003144e-05,
  1.039388e-06, 8.907348e-08, 2.021918e-08, 9.728991e-09, 1.243943e-08, 
    2.18158e-07, 5.932581e-06, 8.476618e-07, 2.667183e-06, 6.997117e-06, 
    1.321667e-05, 1.843144e-05, 1.529798e-05, 1.065983e-05, 9.071809e-06,
  1.206672e-06, 2.547682e-06, 6.915589e-07, 1.433456e-07, 1.190273e-07, 
    1.305965e-06, 2.149003e-06, 1.992414e-05, 1.963278e-05, 4.739533e-06, 
    1.028828e-05, 1.546772e-05, 1.63235e-05, 1.272315e-05, 1.024776e-05,
  4.338297e-06, 3.25868e-06, 1.526686e-06, 1.828606e-06, 9.487197e-07, 
    2.252789e-06, 2.597748e-06, 5.999513e-06, 4.271722e-06, 8.007293e-06, 
    1.01784e-05, 1.205988e-05, 1.332345e-05, 1.203004e-05, 8.859324e-06,
  7.502979e-06, 6.636025e-06, 1.862689e-06, 2.764305e-06, 5.357752e-06, 
    4.576268e-06, 3.538135e-06, 6.588414e-06, 5.475801e-06, 7.460206e-06, 
    1.063341e-05, 1.102461e-05, 1.095012e-05, 8.604708e-06, 7.12066e-06,
  6.576747e-06, 8.754219e-06, 6.871791e-06, 1.725251e-06, 5.427681e-06, 
    3.536813e-06, 3.692096e-06, 2.24785e-06, 6.732589e-06, 8.810019e-06, 
    1.013685e-05, 1.098335e-05, 9.831836e-06, 5.909075e-06, 6.525857e-06,
  8.303829e-06, 8.286767e-06, 3.957961e-06, 2.192751e-06, 5.002963e-06, 
    6.075485e-06, 3.244034e-06, 2.841919e-06, 4.401137e-06, 1.000227e-05, 
    1.080557e-05, 1.262173e-05, 9.431063e-06, 6.514853e-06, 8.047046e-06,
  8.393482e-06, 8.227054e-06, 7.522347e-06, 5.793265e-06, 3.458457e-06, 
    4.638498e-06, 5.046668e-06, 5.661121e-06, 6.473749e-06, 7.538718e-06, 
    1.114515e-05, 1.204353e-05, 1.003626e-05, 8.914363e-06, 1.147573e-05,
  8.106539e-07, 1.374883e-07, 2.925999e-08, 2.613039e-08, 2.079881e-07, 
    4.079815e-07, 7.607626e-07, 1.192991e-06, 1.007046e-06, 9.792086e-06, 
    1.086052e-05, 1.582801e-05, 1.85313e-05, 1.061585e-05, 1.044649e-05,
  2.889866e-07, 3.899455e-07, 5.592565e-07, 7.378401e-07, 1.433504e-06, 
    1.357173e-06, 1.379249e-06, 1.805432e-06, 9.758523e-07, 6.595121e-06, 
    1.166942e-05, 1.83661e-05, 1.623835e-05, 2.313665e-05, 1.912296e-05,
  8.286104e-07, 1.28145e-06, 3.063568e-06, 3.763254e-06, 2.13561e-06, 
    8.434077e-06, 8.916714e-07, 1.097831e-06, 3.543963e-06, 8.950007e-06, 
    9.60748e-06, 1.928566e-05, 1.602209e-05, 1.521196e-05, 1.578794e-05,
  1.458616e-06, 2.116213e-06, 4.362954e-06, 5.694791e-06, 5.230723e-06, 
    5.566933e-06, 7.879244e-06, 9.867703e-07, 3.006491e-06, 1.158566e-05, 
    1.060288e-05, 1.786712e-05, 1.624469e-05, 1.882386e-05, 1.902209e-05,
  1.651747e-06, 6.531037e-06, 6.3391e-06, 4.41987e-06, 4.687502e-06, 
    8.058456e-06, 9.704611e-06, 1.353548e-05, 1.969906e-05, 8.701732e-06, 
    1.508783e-05, 1.460381e-05, 1.765224e-05, 1.690563e-05, 2.287203e-05,
  6.17275e-06, 1.030234e-05, 5.224456e-06, 5.26519e-06, 6.914531e-06, 
    6.675074e-06, 8.243162e-06, 5.809993e-06, 8.391604e-06, 1.381293e-05, 
    1.629746e-05, 1.511163e-05, 1.71242e-05, 1.781108e-05, 2.208649e-05,
  9.866297e-06, 1.094008e-05, 7.197146e-06, 5.424665e-06, 7.312194e-06, 
    7.515446e-06, 6.741453e-06, 7.836456e-06, 9.326747e-06, 9.874485e-06, 
    1.332607e-05, 1.726854e-05, 1.65146e-05, 1.6652e-05, 2.087971e-05,
  1.094817e-05, 9.507081e-06, 5.971923e-06, 7.463601e-06, 7.648416e-06, 
    8.464328e-06, 7.696109e-06, 5.291489e-06, 5.261831e-06, 7.959212e-06, 
    1.303238e-05, 1.718324e-05, 1.677066e-05, 1.563942e-05, 1.356164e-05,
  9.496885e-06, 8.500595e-06, 4.235576e-06, 7.103009e-06, 7.944004e-06, 
    7.988041e-06, 6.667972e-06, 5.170024e-06, 4.051111e-06, 5.913769e-06, 
    1.028561e-05, 1.210516e-05, 1.464839e-05, 1.49274e-05, 1.212624e-05,
  8.867564e-06, 4.716073e-06, 3.80421e-06, 6.288325e-06, 6.724388e-06, 
    6.82839e-06, 9.51919e-06, 8.411502e-06, 4.402285e-06, 7.073937e-06, 
    6.779591e-06, 8.357351e-06, 1.01213e-05, 1.416344e-05, 1.136958e-05,
  3.912873e-07, 1.171671e-06, 1.111175e-06, 1.526e-06, 5.021704e-06, 
    5.751e-06, 6.948166e-06, 5.204474e-06, 4.848241e-06, 4.844692e-06, 
    7.080685e-06, 1.209478e-05, 1.654732e-05, 2.10431e-05, 2.444634e-05,
  1.535228e-06, 2.439141e-06, 3.332889e-06, 4.791045e-06, 6.134288e-06, 
    3.600889e-06, 5.730121e-06, 3.004018e-06, 3.525233e-06, 2.396465e-06, 
    6.986557e-06, 1.303162e-05, 1.655154e-05, 2.401093e-05, 2.156987e-05,
  1.896278e-06, 5.493565e-06, 6.52044e-06, 6.19809e-06, 3.534597e-06, 
    1.174894e-05, 2.303367e-06, 5.810264e-06, 4.719802e-06, 4.045287e-06, 
    6.559704e-06, 1.423777e-05, 1.602781e-05, 1.707578e-05, 1.597914e-05,
  3.977482e-06, 5.262842e-06, 6.322818e-06, 7.232093e-06, 5.284339e-06, 
    6.988974e-06, 1.078588e-05, 2.561141e-06, 3.323439e-06, 3.475985e-06, 
    9.856089e-06, 1.542322e-05, 1.482621e-05, 1.270772e-05, 1.211266e-05,
  3.14157e-06, 5.334869e-06, 6.443129e-06, 7.425245e-06, 7.408913e-06, 
    7.228713e-06, 8.17782e-06, 1.438875e-05, 1.677509e-05, 2.973055e-06, 
    1.282762e-05, 1.541071e-05, 1.355551e-05, 1.023695e-05, 1.120836e-05,
  6.315623e-06, 5.696588e-06, 8.008595e-06, 6.818971e-06, 7.334378e-06, 
    8.7322e-06, 9.742149e-06, 6.930032e-06, 7.168044e-06, 8.713221e-06, 
    1.253782e-05, 1.245592e-05, 1.117562e-05, 1.143769e-05, 1.163867e-05,
  6.454849e-06, 6.386203e-06, 8.579429e-06, 5.07842e-06, 6.818642e-06, 
    8.461419e-06, 5.75271e-06, 5.910701e-06, 6.802131e-06, 5.858045e-06, 
    1.133857e-05, 1.155081e-05, 8.400769e-06, 1.260441e-05, 1.31947e-05,
  6.296748e-06, 7.659074e-06, 7.918297e-06, 6.61858e-06, 7.419943e-06, 
    8.911768e-06, 7.209273e-06, 8.658054e-06, 7.376535e-06, 7.677558e-06, 
    1.221704e-05, 1.170561e-05, 9.650424e-06, 1.149941e-05, 1.336686e-05,
  6.744105e-06, 8.329905e-06, 4.294168e-06, 5.116076e-06, 6.959245e-06, 
    1.119035e-05, 1.20066e-05, 1.401614e-05, 1.389451e-05, 1.208746e-05, 
    1.273605e-05, 1.290032e-05, 1.116189e-05, 8.994254e-06, 8.072378e-06,
  7.01052e-06, 3.746104e-06, 3.229645e-06, 3.985587e-06, 7.679111e-06, 
    1.270544e-05, 1.716967e-05, 1.856431e-05, 1.925597e-05, 2.169897e-05, 
    1.968951e-05, 1.726751e-05, 1.104212e-05, 6.849974e-06, 6.187303e-06,
  4.523477e-07, 2.84189e-06, 2.51169e-06, 3.757545e-06, 4.665817e-06, 
    6.13571e-06, 4.631884e-06, 2.764237e-06, 3.269653e-06, 4.122027e-06, 
    5.208252e-06, 7.667778e-06, 9.380826e-06, 9.772461e-06, 8.578445e-06,
  2.086102e-06, 2.096025e-06, 3.624623e-06, 5.422108e-06, 6.990754e-06, 
    3.184972e-06, 4.832053e-06, 6.425947e-06, 3.440166e-06, 3.737045e-06, 
    5.100059e-06, 6.117238e-06, 9.949886e-06, 1.270385e-05, 8.210641e-06,
  2.463082e-06, 4.246502e-06, 5.082849e-06, 6.531872e-06, 8.10859e-06, 
    1.231325e-05, 2.580346e-06, 1.208483e-05, 1.098918e-05, 6.339234e-06, 
    3.673509e-06, 5.991854e-06, 8.970118e-06, 1.04633e-05, 1.021045e-05,
  3.302465e-06, 2.751296e-06, 7.338667e-06, 8.42078e-06, 8.907754e-06, 
    1.11565e-05, 1.91425e-05, 4.459042e-06, 7.998513e-06, 9.878951e-06, 
    7.950905e-06, 6.808222e-06, 5.420949e-06, 6.892879e-06, 1.018967e-05,
  3.605105e-06, 5.478448e-06, 8.982902e-06, 7.908493e-06, 1.074535e-05, 
    1.402369e-05, 2.538685e-05, 4.375432e-05, 2.688821e-05, 8.590778e-06, 
    1.375939e-05, 9.935065e-06, 7.519395e-06, 7.45953e-06, 1.013786e-05,
  1.532759e-06, 5.983879e-06, 9.266151e-06, 5.265761e-06, 9.648394e-06, 
    1.849179e-05, 3.069185e-05, 3.63882e-05, 2.61169e-05, 2.432897e-05, 
    1.86536e-05, 1.543636e-05, 1.254694e-05, 1.174609e-05, 1.148457e-05,
  3.951091e-06, 8.851625e-06, 5.340657e-06, 5.72618e-06, 7.905971e-06, 
    1.734627e-05, 2.330589e-05, 2.787258e-05, 2.408738e-05, 1.859874e-05, 
    1.763818e-05, 2.001421e-05, 1.919391e-05, 1.702827e-05, 1.392543e-05,
  5.790321e-06, 7.530508e-06, 4.276504e-06, 5.803855e-06, 8.476391e-06, 
    1.46066e-05, 1.709709e-05, 1.760535e-05, 1.768725e-05, 1.742369e-05, 
    1.889086e-05, 1.806882e-05, 1.863872e-05, 2.002047e-05, 1.307769e-05,
  5.659839e-06, 5.389864e-06, 2.75608e-06, 3.517599e-06, 9.146994e-06, 
    1.070963e-05, 1.177676e-05, 1.223795e-05, 1.201516e-05, 1.397621e-05, 
    1.513878e-05, 1.51312e-05, 1.585053e-05, 1.385959e-05, 1.068861e-05,
  3.276266e-06, 2.714169e-06, 1.074057e-06, 1.996846e-06, 4.898937e-06, 
    7.563874e-06, 5.799611e-06, 5.19466e-06, 7.460085e-06, 1.189172e-05, 
    1.480914e-05, 1.381238e-05, 1.405627e-05, 9.950767e-06, 1.084933e-05,
  2.646972e-08, 1.061404e-06, 2.919e-06, 4.583988e-06, 6.103596e-06, 
    6.246332e-06, 4.773686e-06, 6.214832e-06, 9.048165e-06, 1.442293e-05, 
    1.413381e-05, 1.381076e-05, 9.702833e-06, 6.784684e-06, 3.246774e-06,
  6.515451e-07, 2.189315e-06, 3.955533e-06, 5.581296e-06, 7.777316e-06, 
    4.746705e-06, 5.126178e-06, 4.722572e-06, 3.747979e-06, 6.41795e-06, 
    1.32377e-05, 1.582521e-05, 1.027565e-05, 7.3985e-06, 6.26906e-06,
  3.027919e-06, 4.880542e-06, 6.570615e-06, 6.159803e-06, 7.226404e-06, 
    1.431837e-05, 7.940042e-06, 9.692099e-06, 7.314312e-06, 3.775854e-06, 
    6.21242e-06, 1.213979e-05, 1.216251e-05, 4.896308e-06, 3.8792e-06,
  1.680103e-06, 6.837982e-06, 1.018513e-05, 6.23325e-06, 7.525481e-06, 
    1.305957e-05, 2.876801e-05, 1.136175e-05, 1.19985e-05, 6.721481e-06, 
    5.372247e-06, 8.741787e-06, 1.060633e-05, 5.507269e-06, 3.65145e-06,
  4.869759e-06, 8.259743e-06, 1.11789e-05, 4.98807e-06, 7.562994e-06, 
    2.06478e-05, 2.851612e-05, 4.32679e-05, 3.050583e-05, 1.07311e-05, 
    8.622578e-06, 9.523055e-06, 6.619201e-06, 4.35488e-06, 4.570147e-06,
  5.921286e-06, 7.172615e-06, 6.075949e-06, 3.919019e-06, 1.092046e-05, 
    2.632668e-05, 3.88147e-05, 3.465027e-05, 2.011893e-05, 1.222433e-05, 
    1.233974e-05, 8.803908e-06, 8.815192e-06, 6.138552e-06, 4.599481e-06,
  5.786156e-06, 4.835401e-06, 4.483507e-06, 4.470488e-06, 1.124583e-05, 
    2.029341e-05, 3.101377e-05, 3.291586e-05, 2.02127e-05, 1.061858e-05, 
    1.478368e-05, 1.494552e-05, 8.866962e-06, 6.291075e-06, 6.007328e-06,
  4.916373e-06, 8.098643e-06, 5.766863e-06, 2.625685e-06, 1.211312e-05, 
    1.823273e-05, 2.686824e-05, 2.666355e-05, 2.127695e-05, 1.070201e-05, 
    1.120486e-05, 1.55472e-05, 7.082154e-06, 7.264041e-06, 7.199342e-06,
  2.431976e-06, 4.370297e-06, 3.051223e-06, 1.331932e-06, 9.992367e-06, 
    1.863971e-05, 2.102923e-05, 2.756272e-05, 2.385457e-05, 1.109142e-05, 
    1.127476e-05, 1.037486e-05, 5.079833e-06, 5.482505e-06, 8.635976e-06,
  2.84333e-06, 2.152823e-06, 8.249049e-07, 1.29915e-06, 9.165445e-06, 
    1.983229e-05, 2.129568e-05, 2.145857e-05, 2.654881e-05, 2.044459e-05, 
    1.422445e-05, 1.005362e-05, 4.689422e-06, 4.823833e-06, 7.665792e-06,
  5.926337e-07, 2.80349e-06, 4.26311e-06, 2.075071e-06, 1.933895e-06, 
    3.801155e-06, 4.863788e-06, 7.03756e-06, 1.403466e-05, 1.704586e-05, 
    2.218143e-05, 1.275767e-05, 6.374897e-06, 1.320499e-06, 3.151797e-06,
  3.46861e-06, 2.468169e-06, 2.774525e-06, 9.420359e-07, 3.666332e-06, 
    3.100691e-06, 7.05311e-06, 8.890293e-06, 9.244167e-06, 1.639747e-05, 
    1.474127e-05, 1.043121e-05, 7.06135e-06, 4.58399e-06, 4.106098e-06,
  3.852278e-06, 5.926252e-06, 8.000427e-06, 2.300517e-06, 5.589896e-06, 
    2.09324e-05, 7.665009e-06, 1.628302e-05, 1.289808e-05, 1.737995e-05, 
    1.317476e-05, 5.920121e-06, 8.545002e-06, 7.935485e-07, 2.159346e-06,
  5.32653e-06, 7.183799e-06, 8.877419e-06, 3.375422e-06, 6.404915e-06, 
    1.994819e-05, 3.700584e-05, 1.923286e-05, 1.693431e-05, 1.655151e-05, 
    1.458063e-05, 7.905443e-06, 7.058634e-06, 1.870239e-06, 9.40198e-07,
  6.019833e-06, 9.035482e-06, 8.037658e-06, 4.96048e-06, 5.688147e-06, 
    1.519657e-05, 2.343924e-05, 3.60018e-05, 3.060348e-05, 1.054324e-05, 
    1.042496e-05, 6.258771e-06, 3.99692e-06, 1.585641e-06, 9.085427e-07,
  6.739318e-06, 8.608006e-06, 7.546485e-06, 7.023743e-06, 5.516451e-06, 
    9.364065e-06, 1.169902e-05, 1.37007e-05, 1.109931e-05, 6.91497e-06, 
    5.751187e-06, 3.447561e-06, 2.867047e-06, 1.674084e-06, 9.574596e-07,
  8.55896e-06, 1.00457e-05, 6.099426e-06, 6.154239e-06, 3.518101e-06, 
    3.135999e-06, 4.126988e-06, 9.019202e-06, 1.20296e-05, 5.84552e-06, 
    4.642452e-06, 3.550003e-06, 2.69675e-06, 1.814982e-06, 1.047844e-06,
  9.630337e-06, 1.188102e-05, 6.228116e-06, 6.609655e-06, 5.531047e-06, 
    1.428935e-06, 2.902945e-06, 3.575277e-06, 5.204328e-06, 6.037715e-06, 
    4.579042e-06, 5.421771e-06, 2.507439e-06, 1.870058e-06, 8.969197e-07,
  1.045207e-05, 1.037252e-05, 5.965482e-06, 5.570539e-06, 4.767401e-06, 
    9.077019e-07, 1.991374e-06, 5.844438e-06, 5.476812e-06, 4.941832e-06, 
    3.098008e-06, 4.953462e-06, 2.583526e-06, 1.759212e-06, 9.265092e-07,
  9.226315e-06, 6.563863e-06, 4.310464e-06, 3.625379e-06, 4.264242e-06, 
    2.929684e-06, 2.312097e-06, 1.987934e-06, 3.457274e-06, 3.34678e-06, 
    2.940559e-06, 3.680355e-06, 1.963259e-06, 1.762059e-06, 7.340411e-07,
  7.344276e-06, 6.389371e-06, 4.672474e-06, 5.138068e-06, 8.298674e-07, 
    1.335935e-06, 2.795095e-06, 3.885406e-06, 6.941541e-06, 9.71084e-06, 
    9.675191e-06, 3.818655e-06, 1.044008e-06, 1.013216e-07, 7.132709e-06,
  1.180529e-05, 5.146307e-06, 5.083079e-06, 5.396095e-06, 2.13254e-06, 
    1.313664e-06, 2.342632e-06, 3.948339e-06, 6.899731e-06, 9.692156e-06, 
    1.037452e-05, 4.906086e-06, 6.718473e-07, 4.401666e-06, 1.922995e-05,
  1.136784e-05, 6.483189e-06, 6.982447e-06, 7.078588e-06, 9.662381e-07, 
    1.195043e-05, 9.30196e-06, 6.409212e-06, 6.782447e-06, 1.324186e-05, 
    1.041392e-05, 4.968296e-06, 7.135702e-07, 7.795095e-06, 2.90856e-05,
  8.623593e-06, 7.195693e-06, 6.398568e-06, 6.458414e-06, 1.636325e-06, 
    6.006665e-06, 2.700777e-05, 1.524917e-05, 7.555918e-06, 1.790037e-05, 
    1.171647e-05, 5.802456e-06, 2.587439e-06, 1.552161e-05, 2.917876e-05,
  9.550244e-06, 6.896942e-06, 7.344362e-06, 4.90222e-06, 1.902663e-06, 
    3.371019e-06, 3.430805e-06, 2.117881e-05, 3.096764e-05, 1.405821e-05, 
    1.068054e-05, 4.752599e-06, 8.375962e-06, 2.973047e-05, 3.180407e-05,
  9.570016e-06, 8.584212e-06, 6.988756e-06, 3.508608e-06, 1.921092e-06, 
    3.923961e-07, 2.318787e-06, 6.187534e-06, 6.559841e-06, 8.436266e-06, 
    7.462107e-06, 4.78924e-06, 2.391591e-05, 4.501179e-05, 1.805565e-05,
  1.090533e-05, 8.029598e-06, 5.552262e-06, 2.70247e-06, 2.095837e-06, 
    2.839586e-06, 2.45448e-06, 6.28713e-06, 1.549179e-05, 1.031383e-05, 
    8.507224e-06, 2.189135e-05, 4.764558e-05, 4.418943e-05, 2.007477e-05,
  1.003507e-05, 9.480201e-06, 1.93476e-06, 1.60456e-06, 4.725126e-06, 
    3.748888e-06, 4.75888e-06, 1.012375e-05, 1.278897e-05, 1.460423e-05, 
    2.497565e-05, 4.044253e-05, 4.487316e-05, 2.450953e-05, 1.328316e-05,
  1.176642e-05, 5.682937e-06, 1.472846e-06, 3.464019e-06, 3.825111e-06, 
    5.340075e-06, 9.388621e-06, 1.391331e-05, 1.749319e-05, 2.164264e-05, 
    2.487938e-05, 2.607317e-05, 1.955969e-05, 9.470165e-06, 6.618184e-06,
  8.996812e-06, 7.258453e-06, 1.932129e-06, 3.060662e-06, 4.913995e-06, 
    6.73109e-06, 9.8066e-06, 9.060047e-06, 1.025783e-05, 1.556542e-05, 
    1.652353e-05, 1.485053e-05, 1.21573e-05, 7.876954e-06, 6.023457e-06,
  7.895542e-06, 6.709738e-06, 5.401867e-06, 5.575598e-06, 8.00717e-06, 
    8.026652e-06, 2.689595e-06, 2.497016e-06, 2.38503e-06, 1.380975e-06, 
    1.128247e-06, 5.439954e-07, 2.62303e-06, 3.840762e-08, 1.629724e-06,
  2.453137e-05, 1.273342e-05, 1.026212e-05, 9.885386e-06, 6.544662e-06, 
    2.963733e-06, 2.094437e-06, 2.277457e-06, 1.178645e-06, 1.63694e-06, 
    3.158834e-06, 4.099679e-06, 7.278701e-09, 7.264836e-07, 7.548731e-06,
  8.264324e-05, 4.1757e-05, 1.573469e-05, 7.023224e-06, 3.821232e-06, 
    3.178838e-06, 3.61398e-06, 1.32324e-06, 1.471225e-06, 1.572186e-06, 
    1.686653e-06, 2.155909e-06, 2.599735e-08, 5.876609e-07, 1.868363e-05,
  8.311804e-05, 3.066171e-05, 6.643072e-06, 3.492285e-06, 4.084097e-06, 
    3.614534e-06, 1.298233e-05, 1.317068e-05, 3.10366e-06, 1.608414e-06, 
    1.06663e-06, 6.310058e-07, 5.874281e-08, 1.742092e-06, 2.041106e-05,
  2.395574e-05, 7.261128e-06, 4.782446e-06, 3.944346e-06, 4.055746e-06, 
    4.958363e-06, 1.307482e-06, 2.746211e-05, 1.555009e-05, 2.020484e-06, 
    1.400563e-06, 8.305323e-07, 4.429626e-07, 6.453301e-06, 1.713445e-05,
  8.760189e-06, 9.93956e-06, 6.474291e-06, 4.599454e-06, 5.151265e-07, 
    1.642915e-06, 3.171521e-06, 1.69121e-06, 1.218961e-06, 6.620139e-07, 
    1.741478e-07, 3.663247e-07, 4.079476e-06, 1.769048e-05, 3.901438e-06,
  1.009894e-05, 1.024832e-05, 5.47468e-06, 5.393103e-06, 8.270485e-07, 
    9.919642e-07, 1.575261e-06, 1.249824e-06, 8.45049e-07, 1.880355e-07, 
    9.258957e-07, 6.734335e-06, 2.158974e-05, 1.20755e-05, 2.825924e-06,
  8.058072e-06, 9.066483e-06, 1.663057e-06, 1.73959e-06, 3.263511e-06, 
    5.948525e-06, 4.11133e-06, 3.915728e-06, 3.173073e-06, 4.676894e-06, 
    1.269204e-05, 2.482642e-05, 2.466742e-05, 3.751073e-06, 2.531953e-06,
  1.233086e-05, 4.98117e-06, 2.887424e-06, 4.876227e-06, 7.051634e-06, 
    1.052188e-05, 9.958942e-06, 1.129246e-05, 1.051033e-05, 2.301504e-05, 
    3.443976e-05, 3.04055e-05, 1.020596e-05, 3.812564e-06, 2.357185e-06,
  8.773099e-06, 9.077756e-06, 4.043794e-06, 6.867982e-06, 1.322332e-05, 
    1.555212e-05, 1.774566e-05, 1.708184e-05, 2.881955e-05, 4.523864e-05, 
    3.946312e-05, 1.621033e-05, 6.161652e-06, 4.186171e-06, 3.278574e-06,
  4.338736e-05, 9.652389e-06, 1.676138e-06, 8.531437e-09, 1.733245e-07, 
    6.455188e-07, 8.424939e-07, 7.555849e-07, 1.127039e-06, 2.590594e-06, 
    2.310843e-06, 3.232198e-07, 1.154162e-08, 7.019412e-07, 1.481848e-06,
  4.298279e-05, 1.069826e-05, 5.85825e-07, 7.755375e-07, 1.878989e-06, 
    1.967865e-06, 1.315584e-06, 1.274746e-06, 8.466635e-07, 1.293043e-07, 
    3.335504e-07, 1.582101e-07, 3.355454e-08, 1.978448e-06, 7.507722e-06,
  4.634236e-05, 8.830412e-06, 4.024019e-06, 4.107579e-06, 2.11275e-06, 
    4.575499e-06, 4.29191e-06, 2.768255e-06, 7.950787e-07, 4.90163e-07, 
    2.059679e-06, 4.695813e-07, 6.750079e-07, 2.996056e-06, 3.442677e-05,
  8.351645e-05, 4.738573e-05, 2.139416e-05, 1.517785e-05, 1.449024e-05, 
    2.187422e-06, 9.322008e-06, 2.783185e-06, 1.472708e-06, 7.138196e-07, 
    2.13731e-07, 1.977024e-07, 1.78261e-06, 1.149165e-05, 4.335975e-05,
  8.47785e-05, 5.10553e-05, 3.351742e-05, 2.523362e-05, 1.979493e-05, 
    9.243931e-06, 8.218272e-07, 5.464954e-06, 3.823761e-06, 3.990832e-07, 
    7.124697e-07, 1.237665e-06, 3.923798e-06, 2.252767e-05, 2.805983e-05,
  2.648435e-05, 2.697423e-05, 2.349529e-05, 1.800237e-05, 8.798283e-06, 
    4.924282e-06, 2.023671e-06, 3.659367e-07, 2.20592e-07, 8.963985e-08, 
    9.125463e-08, 1.567766e-06, 1.279836e-05, 1.975784e-05, 7.883454e-06,
  9.255647e-06, 1.009504e-05, 6.629948e-06, 4.409793e-06, 3.879672e-06, 
    3.170102e-06, 2.429147e-06, 1.76054e-07, 9.678103e-07, 3.2867e-06, 
    1.095783e-06, 6.061148e-06, 2.590096e-05, 5.498563e-06, 3.366831e-06,
  8.169873e-06, 6.452491e-06, 2.749292e-07, 2.028877e-06, 3.658773e-06, 
    2.926256e-06, 1.31694e-06, 2.122061e-07, 3.050658e-08, 5.861215e-07, 
    2.090727e-06, 2.099842e-05, 1.587204e-05, 3.760456e-06, 3.22399e-06,
  7.622808e-06, 4.409098e-06, 1.608644e-06, 2.482359e-06, 2.859235e-06, 
    1.388927e-06, 1.132063e-06, 7.64462e-07, 7.85692e-07, 1.73918e-06, 
    6.437728e-06, 2.377122e-05, 1.032071e-05, 5.833641e-06, 4.279034e-06,
  6.951736e-06, 5.874231e-06, 4.137132e-06, 4.551218e-06, 2.884079e-06, 
    6.601549e-07, 2.207081e-06, 4.440734e-07, 3.854245e-07, 3.566779e-06, 
    1.779001e-05, 1.83241e-05, 1.374272e-05, 1.168039e-05, 7.061196e-06,
  3.121014e-05, 1.350647e-06, 3.937793e-06, 1.216645e-05, 1.187108e-05, 
    3.420775e-06, 1.574205e-06, 7.805852e-08, 1.559472e-07, 5.704311e-07, 
    1.416022e-06, 8.733524e-07, 9.574451e-07, 2.052045e-06, 3.652099e-06,
  4.340641e-06, 6.136947e-06, 1.158773e-05, 2.311699e-05, 2.78405e-05, 
    7.72867e-06, 1.714813e-06, 4.937287e-07, 2.789099e-07, 9.806179e-07, 
    1.320379e-06, 1.301117e-06, 1.809396e-06, 4.929678e-06, 5.833524e-06,
  1.783823e-05, 2.767351e-05, 3.166177e-05, 3.92641e-05, 2.20303e-05, 
    1.965396e-05, 2.202906e-06, 1.211239e-06, 1.379448e-06, 1.342161e-06, 
    1.1482e-06, 1.157802e-06, 2.912061e-06, 5.942347e-06, 8.838418e-06,
  4.902093e-05, 5.37404e-05, 5.239122e-05, 4.392569e-05, 3.781723e-05, 
    2.636676e-06, 1.191288e-05, 4.043151e-06, 1.522286e-06, 5.654209e-07, 
    8.042263e-08, 2.098472e-06, 4.673119e-06, 4.011887e-06, 1.105087e-05,
  7.186081e-05, 6.428784e-05, 7.044246e-05, 4.223268e-05, 4.616623e-05, 
    7.446478e-06, 6.481993e-07, 1.805258e-06, 2.426912e-06, 1.052925e-07, 
    1.129096e-07, 1.825519e-06, 6.742845e-06, 1.434762e-05, 1.937298e-05,
  9.334298e-05, 6.406202e-05, 7.052271e-05, 3.888652e-05, 2.334073e-05, 
    5.939933e-06, 8.320415e-07, 1.995717e-07, 8.152585e-08, 9.206747e-08, 
    2.841307e-06, 3.679169e-06, 1.161034e-05, 1.874448e-05, 1.550687e-05,
  9.313328e-05, 7.941599e-05, 7.397558e-05, 3.465098e-05, 1.351281e-05, 
    2.145395e-06, 3.989206e-07, 3.212188e-07, 2.040576e-06, 2.311828e-06, 
    4.182796e-06, 8.732144e-06, 1.255106e-05, 1.580167e-05, 1.188699e-05,
  8.111116e-05, 8.233149e-05, 5.38003e-05, 2.573213e-05, 8.614518e-06, 
    1.808565e-06, 2.907703e-07, 2.70523e-07, 2.1296e-07, 2.426401e-07, 
    3.19413e-06, 9.716211e-06, 9.44778e-06, 1.201859e-05, 1.390734e-05,
  6.593615e-05, 4.521498e-05, 3.348492e-05, 2.127185e-05, 9.145507e-06, 
    3.429547e-06, 4.078375e-07, 1.956933e-08, 2.82637e-07, 1.23111e-06, 
    2.569246e-06, 7.107279e-06, 2.786697e-06, 4.643927e-06, 1.445775e-05,
  4.417586e-05, 2.812409e-05, 2.459428e-05, 1.635117e-05, 8.949819e-06, 
    4.047391e-06, 1.326214e-06, 4.656348e-09, 3.098256e-08, 8.091889e-07, 
    6.275515e-06, 6.906662e-06, 3.496206e-06, 9.555836e-06, 2.71675e-05,
  0.0002113222, 0.0001145875, 3.003439e-05, 2.609931e-05, 8.583514e-05, 
    7.893132e-05, 4.049469e-05, 3.39929e-05, 1.94006e-05, 6.343992e-06, 
    1.223202e-06, 1.464819e-07, 4.5976e-07, 7.91421e-07, 8.123135e-07,
  0.0002139223, 8.386411e-05, 3.052607e-05, 4.303544e-05, 7.994242e-05, 
    6.182535e-05, 4.798458e-05, 4.282839e-05, 2.2181e-05, 4.45474e-06, 
    1.399935e-06, 6.640398e-07, 7.22814e-07, 7.913197e-07, 7.848607e-07,
  0.0001130912, 7.127326e-05, 4.000849e-05, 5.054593e-05, 4.131992e-05, 
    7.82345e-05, 5.635581e-05, 5.163649e-05, 2.317318e-05, 3.403051e-06, 
    1.189264e-06, 7.310713e-07, 4.825101e-07, 7.829873e-07, 2.549943e-06,
  0.0001049201, 6.664647e-05, 3.136679e-05, 3.709766e-05, 3.360808e-05, 
    3.427682e-06, 6.743347e-05, 3.325725e-05, 1.039933e-05, 1.453668e-06, 
    7.356713e-07, 8.029025e-07, 6.256373e-07, 5.080493e-07, 4.714198e-06,
  8.645145e-05, 4.712394e-05, 1.482407e-05, 2.189291e-05, 3.809252e-05, 
    2.115236e-05, 9.2825e-07, 2.444664e-06, 5.641452e-06, 1.465608e-06, 
    7.282003e-07, 3.627026e-07, 4.054804e-06, 5.751867e-06, 1.116721e-05,
  3.843896e-05, 1.17567e-05, 4.442732e-06, 1.041467e-05, 1.555528e-05, 
    1.06603e-05, 1.220463e-06, 8.113168e-08, 9.215588e-08, 4.230787e-07, 
    1.26016e-06, 9.21188e-07, 9.525153e-06, 1.22102e-05, 1.266241e-05,
  2.106689e-05, 9.944149e-06, 1.233575e-05, 9.504382e-06, 5.826416e-06, 
    2.337511e-06, 9.389067e-07, 1.061066e-06, 1.127842e-06, 2.803858e-06, 
    1.742747e-06, 7.158165e-06, 1.2435e-05, 6.790042e-06, 5.069112e-06,
  2.365056e-05, 2.421536e-05, 2.213557e-05, 3.632741e-06, 2.839994e-06, 
    1.038214e-06, 5.763507e-07, 7.631073e-07, 1.435176e-06, 2.148287e-06, 
    1.007068e-05, 5.503626e-06, 7.778077e-06, 9.640227e-06, 1.15372e-05,
  4.180657e-05, 4.460938e-05, 1.430006e-05, 3.733556e-06, 3.013039e-06, 
    2.487383e-06, 2.69529e-06, 3.631697e-06, 2.964999e-06, 6.265465e-06, 
    6.079433e-06, 4.846755e-06, 6.642627e-06, 1.225938e-05, 1.898379e-05,
  6.938841e-05, 2.688162e-05, 4.730759e-06, 3.369776e-06, 2.956067e-06, 
    2.497551e-06, 3.52892e-06, 5.131539e-06, 5.528585e-06, 4.583209e-06, 
    3.423335e-06, 3.818571e-06, 6.942985e-06, 1.242567e-05, 1.337194e-05,
  1.31786e-06, 8.630015e-07, 2.020291e-06, 0.0001004908, 8.379132e-05, 
    8.287871e-06, 7.602714e-06, 3.116684e-05, 0.000115177, 0.0001267818, 
    1.9862e-05, 2.965577e-07, 1.940224e-07, 3.494416e-06, 5.768429e-06,
  5.448451e-05, 1.529499e-05, 2.313657e-06, 1.924741e-05, 1.315856e-06, 
    1.151377e-06, 6.446797e-06, 2.858551e-05, 8.983369e-05, 0.0001562026, 
    4.696885e-05, 4.680359e-06, 1.017868e-07, 1.267496e-06, 3.110017e-06,
  4.450688e-05, 9.872416e-06, 2.770097e-06, 2.530272e-06, 7.4485e-07, 
    2.30474e-06, 2.770083e-06, 3.421729e-05, 0.0001035505, 0.0001715561, 
    0.0001093117, 1.753107e-05, 3.900607e-06, 2.032632e-07, 1.7829e-06,
  1.157105e-05, 3.771173e-06, 3.273548e-06, 2.293609e-06, 1.28769e-06, 
    6.985413e-07, 2.741573e-05, 5.588908e-05, 9.963413e-05, 0.0001135662, 
    0.0001144716, 4.515129e-05, 9.150951e-06, 4.276225e-07, 1.332105e-06,
  1.09915e-05, 6.554352e-06, 7.350328e-06, 6.874904e-06, 8.742698e-06, 
    1.86186e-05, 1.163365e-05, 4.975027e-05, 8.76562e-05, 4.47849e-05, 
    7.636067e-05, 7.341934e-05, 2.384125e-05, 7.476158e-06, 2.747016e-06,
  1.536372e-05, 1.515523e-05, 1.154854e-05, 1.035507e-05, 9.283849e-06, 
    2.112604e-05, 2.424164e-05, 7.396187e-06, 1.457153e-05, 6.474983e-05, 
    4.182907e-05, 6.928142e-05, 6.403251e-05, 3.095257e-05, 8.055739e-06,
  8.802214e-06, 1.269607e-05, 1.643112e-05, 1.908315e-05, 1.878765e-05, 
    2.966009e-05, 6.071846e-05, 0.0001104034, 0.0001051587, 6.082495e-05, 
    4.421376e-05, 4.507462e-05, 3.987291e-05, 1.911724e-05, 6.644385e-06,
  5.939214e-06, 1.034955e-05, 1.771901e-05, 2.393526e-05, 2.824839e-05, 
    2.88267e-05, 2.25266e-05, 2.286982e-05, 2.188398e-05, 1.654145e-05, 
    1.16318e-05, 9.204033e-06, 7.371837e-06, 5.887997e-06, 3.694526e-06,
  6.744292e-06, 6.976892e-06, 7.919195e-06, 8.654553e-06, 6.259821e-06, 
    3.943785e-06, 3.593305e-06, 4.072404e-06, 3.614938e-06, 3.328968e-06, 
    2.433589e-06, 3.144558e-06, 4.543335e-06, 5.836301e-06, 3.825598e-06,
  2.114916e-06, 3.572456e-06, 4.460374e-06, 4.089978e-06, 4.019782e-06, 
    3.94021e-06, 3.45161e-06, 3.362335e-06, 2.661293e-06, 3.103098e-06, 
    3.780812e-06, 7.474986e-06, 5.023797e-06, 4.682877e-06, 5.787593e-06,
  8.970062e-06, 8.024747e-06, 6.715713e-06, 7.846768e-05, 0.0001478834, 
    6.235861e-05, 1.07843e-05, 2.765415e-06, 4.353412e-06, 1.82245e-05, 
    2.81722e-06, 1.308699e-06, 3.119668e-07, 2.014489e-06, 1.718482e-06,
  5.667334e-06, 5.697173e-06, 2.658954e-05, 0.00014446, 0.0001447652, 
    6.939075e-05, 3.481226e-05, 7.932595e-06, 7.956173e-06, 1.626835e-05, 
    5.959112e-06, 6.050012e-07, 3.932473e-07, 3.243607e-06, 4.291542e-06,
  7.611137e-06, 2.849901e-05, 9.448864e-05, 0.0001526904, 0.0001175295, 
    9.114653e-05, 3.647436e-05, 2.492966e-05, 2.039342e-05, 2.365303e-05, 
    6.848669e-06, 2.162995e-06, 3.412455e-07, 1.926227e-06, 3.335604e-06,
  8.050841e-06, 1.663684e-05, 5.118054e-05, 0.0001393521, 0.0001250141, 
    6.419563e-05, 6.187573e-05, 2.421743e-05, 3.000011e-05, 4.341259e-05, 
    1.101433e-05, 1.996903e-06, 1.104118e-06, 5.174729e-06, 3.341695e-06,
  5.085238e-06, 5.751572e-06, 2.042528e-05, 8.580886e-05, 8.798151e-05, 
    6.389927e-05, 9.170407e-06, 1.182843e-05, 5.902087e-05, 5.144083e-05, 
    3.161605e-05, 1.084999e-05, 3.776793e-06, 5.607359e-06, 4.167421e-06,
  7.996578e-06, 9.408252e-06, 1.401796e-05, 2.966215e-05, 4.563672e-05, 
    3.197346e-05, 9.135611e-06, 2.694302e-06, 2.035619e-06, 3.710618e-05, 
    5.930583e-05, 4.184111e-05, 2.663478e-05, 7.568274e-06, 6.530605e-06,
  8.366725e-06, 1.13026e-05, 1.281126e-05, 1.943487e-05, 3.908251e-05, 
    3.03168e-05, 1.210928e-05, 6.926763e-06, 1.42544e-05, 4.369254e-05, 
    6.418446e-05, 7.585368e-05, 5.67967e-05, 3.594166e-05, 9.981125e-06,
  8.455397e-06, 8.210334e-06, 1.362451e-05, 1.895524e-05, 3.071647e-05, 
    4.377947e-05, 2.398986e-05, 1.352184e-05, 1.910232e-05, 5.167384e-05, 
    6.519025e-05, 6.839605e-05, 9.221478e-05, 7.937625e-05, 4.971685e-05,
  6.072714e-06, 4.329478e-06, 7.604378e-06, 8.232397e-06, 1.304136e-05, 
    2.24878e-05, 2.732184e-05, 2.349389e-05, 2.164824e-05, 4.313601e-05, 
    4.641791e-05, 5.001905e-05, 6.706622e-05, 6.504409e-05, 5.856044e-05,
  2.866576e-06, 2.58372e-06, 2.793606e-06, 2.827046e-06, 3.303822e-06, 
    5.099478e-06, 8.175732e-06, 1.087401e-05, 1.112991e-05, 1.797708e-05, 
    2.167056e-05, 2.261678e-05, 2.714252e-05, 2.724957e-05, 2.862432e-05,
  8.290558e-06, 7.822549e-06, 7.262534e-06, 9.317696e-06, 6.432711e-06, 
    2.236152e-06, 4.834541e-07, 6.045839e-08, 1.269181e-08, 5.517218e-07, 
    1.523903e-06, 1.716643e-05, 5.589139e-06, 3.388943e-06, 7.732552e-07,
  1.01655e-05, 9.990745e-06, 1.078138e-05, 1.159371e-05, 8.405423e-06, 
    9.35401e-06, 8.721107e-07, 6.959448e-08, 2.49697e-08, 1.032198e-06, 
    8.459922e-07, 1.547759e-05, 5.492011e-06, 4.218291e-06, 1.077756e-06,
  8.598439e-06, 1.104004e-05, 2.572215e-05, 2.201596e-05, 1.486453e-05, 
    1.933037e-05, 3.948659e-06, 1.079047e-06, 4.39583e-07, 6.978651e-07, 
    2.637287e-07, 9.950127e-06, 3.753661e-06, 1.294217e-06, 8.661851e-08,
  9.958285e-06, 1.150108e-05, 3.725536e-05, 4.787864e-05, 3.274052e-05, 
    8.021841e-06, 1.715147e-05, 5.511195e-06, 2.010594e-06, 3.019829e-07, 
    5.265642e-07, 9.708701e-06, 3.348729e-06, 1.860299e-06, 2.013154e-07,
  8.84516e-06, 1.053314e-05, 3.724795e-05, 6.75449e-05, 5.837076e-05, 
    2.129399e-05, 2.13129e-06, 2.323383e-05, 1.222441e-05, 1.155495e-07, 
    5.880081e-07, 6.712001e-06, 5.131983e-06, 2.539621e-06, 1.221226e-06,
  1.080438e-05, 1.613595e-05, 2.919837e-05, 4.394999e-05, 4.269119e-05, 
    2.158594e-05, 2.807358e-06, 2.212151e-07, 5.185376e-07, 1.227409e-07, 
    2.920928e-07, 4.38641e-06, 4.144098e-06, 3.884815e-06, 2.497266e-06,
  1.368521e-05, 1.951996e-05, 3.343062e-05, 3.945988e-05, 3.734825e-05, 
    2.381297e-05, 3.41346e-06, 6.309243e-07, 6.228528e-07, 1.720766e-07, 
    9.258977e-07, 5.127358e-06, 4.784124e-06, 6.754755e-06, 3.977434e-06,
  1.492074e-05, 2.179316e-05, 4.268641e-05, 5.011417e-05, 5.773428e-05, 
    4.288991e-05, 7.256131e-06, 1.437733e-06, 7.093695e-07, 9.144026e-07, 
    2.006112e-06, 6.137424e-06, 6.343017e-06, 8.595436e-06, 8.472906e-06,
  1.483766e-05, 2.714774e-05, 4.799396e-05, 6.832034e-05, 7.963824e-05, 
    6.203664e-05, 2.609861e-05, 8.16008e-06, 5.035623e-06, 1.470606e-05, 
    2.020996e-05, 6.487334e-06, 7.191812e-06, 9.797674e-06, 1.212546e-05,
  1.192534e-05, 2.530381e-05, 4.822528e-05, 6.268195e-05, 6.778711e-05, 
    6.354198e-05, 4.083433e-05, 1.911271e-05, 1.73753e-05, 3.213361e-05, 
    3.173972e-05, 1.144127e-05, 1.044275e-05, 1.180327e-05, 1.328066e-05,
  3.472713e-07, 1.159877e-06, 7.81355e-07, 3.761231e-06, 3.316383e-06, 
    1.956326e-06, 2.551845e-06, 3.468517e-06, 3.896267e-06, 1.327e-06, 
    3.07475e-07, 2.83625e-06, 2.158117e-05, 4.949829e-05, 6.396668e-05,
  1.496799e-07, 3.333101e-07, 2.359845e-06, 4.618273e-06, 7.471235e-06, 
    3.022918e-06, 1.816052e-06, 2.600732e-06, 2.449357e-06, 1.589368e-06, 
    3.331382e-07, 7.35161e-06, 3.358743e-05, 7.301837e-05, 7.617828e-05,
  2.532328e-06, 1.65361e-06, 3.787832e-06, 4.096613e-06, 6.146458e-06, 
    1.623433e-05, 2.04173e-06, 1.503026e-06, 1.439246e-06, 9.929064e-07, 
    1.176186e-06, 2.491709e-05, 5.416349e-05, 7.921879e-05, 8.091572e-05,
  2.783071e-06, 2.986276e-06, 4.690554e-06, 6.321613e-06, 9.783455e-06, 
    1.279147e-05, 1.327661e-05, 3.257519e-06, 2.431606e-06, 3.695016e-07, 
    4.760427e-06, 4.736019e-05, 6.784906e-05, 9.270412e-05, 6.997376e-05,
  4.771518e-06, 1.007536e-05, 6.350603e-06, 4.786916e-06, 6.492722e-06, 
    1.59086e-05, 7.585353e-06, 1.227576e-05, 8.496408e-06, 7.447668e-07, 
    1.772965e-05, 6.807232e-05, 7.138098e-05, 5.640325e-05, 2.577782e-05,
  1.684173e-05, 1.731847e-05, 1.302306e-05, 9.070111e-06, 6.129214e-06, 
    9.442996e-06, 7.915005e-06, 9.337988e-07, 2.93471e-07, 1.605929e-07, 
    3.221192e-05, 7.436339e-05, 5.422825e-05, 1.798088e-05, 2.445913e-06,
  1.928926e-05, 2.372843e-05, 1.903972e-05, 1.089759e-05, 5.731958e-06, 
    7.846432e-06, 6.294898e-06, 2.559454e-06, 2.180143e-06, 1.575763e-06, 
    5.225163e-05, 6.141272e-05, 2.08588e-05, 3.868197e-06, 2.207006e-06,
  1.834382e-05, 2.417997e-05, 1.962677e-05, 8.190964e-06, 7.725798e-06, 
    1.095513e-05, 5.936305e-06, 1.41802e-06, 8.222893e-07, 1.935909e-05, 
    5.904615e-05, 2.738099e-05, 5.294511e-06, 3.655412e-06, 4.608925e-06,
  1.537749e-05, 2.355642e-05, 2.623865e-05, 1.765342e-05, 1.639454e-05, 
    1.446516e-05, 6.768009e-06, 6.319514e-07, 5.191992e-06, 3.104529e-05, 
    4.58089e-05, 7.71481e-06, 4.447608e-06, 4.602469e-06, 7.274705e-06,
  1.090825e-05, 1.952959e-05, 3.000567e-05, 2.809484e-05, 2.320253e-05, 
    1.299441e-05, 3.670598e-06, 1.135965e-06, 4.962305e-06, 1.73732e-05, 
    2.369461e-05, 5.823147e-06, 4.98175e-06, 7.493432e-06, 8.751144e-06,
  3.908692e-06, 3.778584e-06, 3.958631e-06, 3.051723e-06, 2.360186e-06, 
    2.089355e-06, 1.455399e-06, 1.633656e-06, 2.40714e-06, 4.932377e-06, 
    4.24995e-06, 3.187641e-06, 3.700365e-06, 2.177717e-06, 4.574229e-06,
  7.589335e-07, 4.138884e-07, 5.077612e-07, 1.206531e-06, 2.266883e-06, 
    1.882712e-06, 1.339251e-06, 2.363679e-06, 3.596122e-06, 3.646161e-06, 
    1.989688e-06, 1.228086e-06, 1.549484e-06, 5.119702e-06, 4.192392e-06,
  1.261664e-07, 3.274246e-08, 8.063184e-07, 1.968847e-06, 2.956954e-06, 
    5.864394e-06, 5.03765e-07, 1.06446e-06, 1.500865e-06, 1.029421e-06, 
    7.993705e-07, 6.635937e-07, 3.256222e-06, 2.184649e-06, 6.092805e-06,
  1.073137e-07, 6.254319e-07, 2.154371e-06, 3.035072e-06, 4.741313e-06, 
    4.64601e-06, 1.1117e-05, 9.096759e-07, 3.66387e-07, 2.530349e-07, 
    3.348684e-07, 2.512429e-06, 1.304443e-05, 8.594911e-06, 1.660594e-05,
  7.109643e-07, 4.041649e-06, 7.534967e-06, 8.916758e-06, 1.084274e-05, 
    1.966459e-05, 1.197095e-05, 3.506378e-05, 5.638339e-06, 7.616785e-07, 
    7.38054e-07, 1.385304e-05, 3.773831e-05, 2.072387e-05, 3.560722e-05,
  4.081059e-06, 1.130967e-05, 1.370579e-05, 1.212152e-05, 8.642119e-06, 
    7.658015e-06, 1.041002e-05, 1.787697e-06, 9.161816e-07, 8.571641e-07, 
    2.340752e-06, 4.197969e-05, 5.470482e-05, 2.622007e-05, 1.994801e-05,
  7.825077e-06, 1.077143e-05, 9.777444e-06, 1.102959e-05, 8.610867e-06, 
    5.45971e-06, 5.50994e-06, 6.194572e-06, 4.841583e-06, 2.014178e-06, 
    2.244983e-05, 7.103716e-05, 4.855235e-05, 1.397276e-05, 1.259776e-05,
  1.068892e-05, 1.109107e-05, 4.726063e-06, 4.18728e-06, 4.942785e-06, 
    4.661038e-06, 3.319984e-06, 4.896723e-06, 3.45338e-06, 8.315069e-06, 
    7.371239e-05, 6.673652e-05, 2.164971e-05, 1.009179e-05, 9.085303e-06,
  1.156579e-05, 5.550651e-06, 4.156227e-06, 3.661475e-06, 4.206776e-06, 
    3.759696e-06, 4.571931e-06, 4.601665e-06, 1.055532e-05, 5.209296e-05, 
    7.992285e-05, 3.466556e-05, 8.042593e-06, 8.160477e-06, 3.079128e-06,
  6.000434e-06, 7.445579e-06, 5.125473e-06, 3.235878e-06, 3.14443e-06, 
    4.389287e-06, 5.970431e-06, 1.126657e-05, 4.585152e-05, 9.094828e-05, 
    4.721541e-05, 9.79133e-06, 7.553771e-06, 4.570599e-06, 3.789345e-07,
  0.0001081594, 7.650707e-05, 5.391962e-05, 3.164092e-05, 2.149284e-05, 
    6.002922e-06, 4.05526e-06, 2.975958e-06, 4.269033e-06, 1.005071e-06, 
    1.429176e-06, 1.793098e-06, 1.431754e-06, 6.103737e-07, 4.350245e-06,
  0.0001555561, 8.088604e-05, 5.561955e-05, 3.776797e-05, 1.737194e-05, 
    4.956497e-06, 1.248297e-06, 2.885675e-06, 3.582628e-06, 1.042864e-06, 
    8.442415e-07, 4.655374e-07, 9.516254e-07, 4.074163e-06, 2.220686e-05,
  0.0002435826, 9.811465e-05, 2.877013e-05, 2.750908e-05, 1.805144e-05, 
    1.992673e-05, 2.866127e-06, 8.391329e-07, 1.072269e-06, 6.516879e-07, 
    9.930444e-07, 3.556431e-08, 2.376008e-06, 5.47039e-06, 6.874976e-05,
  0.0002311492, 0.0001540563, 3.964918e-05, 1.127577e-05, 1.113391e-05, 
    9.380189e-07, 2.20334e-05, 4.29776e-07, 8.620593e-08, 1.750201e-08, 
    2.677238e-09, 4.832201e-09, 3.599806e-06, 6.752647e-06, 9.735669e-05,
  6.465123e-05, 7.827678e-05, 4.148381e-05, 1.001558e-05, 6.528474e-06, 
    7.50089e-06, 2.503431e-06, 1.42165e-05, 2.806888e-06, 1.977354e-08, 
    2.827901e-08, 1.112465e-07, 1.939793e-06, 6.793946e-06, 6.325773e-05,
  6.960008e-07, 4.177937e-06, 5.093906e-06, 3.734901e-06, 3.068282e-06, 
    4.224704e-06, 6.152459e-06, 1.965678e-06, 2.381435e-07, 1.023895e-07, 
    1.316101e-07, 3.27988e-06, 3.089769e-06, 6.488798e-06, 1.630041e-05,
  2.429915e-06, 3.74408e-06, 4.423493e-06, 4.482871e-06, 4.626642e-06, 
    3.894159e-06, 5.145163e-06, 8.660514e-06, 3.876296e-06, 5.143983e-07, 
    2.524543e-07, 9.290566e-07, 3.325821e-06, 8.335894e-06, 1.01929e-05,
  1.013725e-06, 5.015831e-06, 3.463879e-06, 4.627167e-06, 4.277888e-06, 
    4.656695e-06, 4.634829e-06, 4.466349e-06, 3.39724e-06, 6.420412e-07, 
    1.622815e-06, 1.530081e-06, 5.97588e-06, 8.89488e-06, 7.558565e-06,
  2.964614e-06, 8.805739e-06, 1.111722e-05, 1.147567e-05, 1.211668e-05, 
    9.442761e-06, 6.219278e-06, 4.280007e-06, 3.058806e-06, 1.520031e-06, 
    7.998305e-07, 2.867912e-06, 5.535902e-06, 8.395293e-06, 5.632386e-06,
  5.840627e-06, 2.401578e-05, 2.638901e-05, 2.313442e-05, 2.023618e-05, 
    1.58146e-05, 7.28923e-06, 3.980022e-06, 4.866596e-06, 1.761644e-06, 
    8.792509e-07, 3.933916e-06, 5.855939e-06, 1.014388e-05, 2.510395e-06,
  3.340001e-05, 3.226859e-05, 4.847837e-05, 0.00014287, 0.0001312251, 
    9.749053e-05, 7.897235e-05, 5.728327e-05, 2.17409e-05, 6.309074e-06, 
    4.348211e-07, 1.882424e-08, 1.43743e-07, 3.303874e-06, 6.174172e-06,
  7.606853e-05, 3.338964e-05, 5.494629e-05, 9.89523e-05, 8.434065e-05, 
    8.309961e-05, 5.378892e-05, 2.225498e-05, 7.599494e-06, 3.779239e-06, 
    9.285998e-08, 8.235298e-07, 1.773178e-06, 5.973086e-06, 6.379086e-06,
  0.0001437772, 6.610037e-05, 6.981823e-05, 8.38466e-05, 3.726858e-05, 
    5.589697e-05, 1.886732e-05, 7.873966e-06, 4.408619e-06, 1.008208e-06, 
    1.030895e-06, 1.794554e-06, 1.802053e-06, 5.210684e-06, 2.356081e-06,
  0.0001944586, 0.0001593125, 0.0001103443, 7.627908e-05, 4.724378e-05, 
    6.314529e-06, 3.344057e-05, 1.144985e-05, 2.140102e-06, 9.365223e-07, 
    1.850003e-06, 2.097742e-06, 2.850266e-06, 6.037331e-06, 4.979602e-06,
  0.0001435317, 0.0002556331, 0.0001942703, 8.980372e-05, 5.171655e-05, 
    2.505156e-05, 2.743892e-06, 1.129633e-05, 6.23597e-06, 2.396444e-06, 
    1.544003e-06, 3.028772e-06, 4.885042e-06, 5.907547e-06, 6.78019e-06,
  2.51026e-05, 0.0002254853, 0.0002379092, 9.650859e-05, 4.208794e-05, 
    3.493145e-05, 2.309319e-05, 4.233603e-06, 8.482265e-07, 1.201391e-06, 
    1.51049e-06, 2.008898e-06, 4.935785e-06, 7.132558e-06, 6.488201e-06,
  4.1317e-06, 0.0001188884, 0.000234859, 0.0001062806, 2.565285e-05, 
    1.485951e-05, 2.969966e-05, 1.010451e-05, 2.772539e-06, 1.365584e-06, 
    1.68233e-06, 4.107156e-06, 6.214811e-06, 9.315527e-06, 7.828132e-06,
  4.370704e-07, 3.216999e-05, 0.0001939245, 0.0001397285, 2.226021e-05, 
    9.247733e-06, 4.799681e-06, 1.239574e-06, 9.306313e-07, 7.889881e-07, 
    1.99165e-06, 3.009506e-06, 7.531637e-06, 8.776196e-06, 7.215312e-06,
  2.392124e-06, 8.093954e-06, 0.0001213035, 0.0001409431, 3.239936e-05, 
    8.765348e-06, 3.784539e-06, 1.663552e-06, 1.724382e-06, 1.580014e-06, 
    5.648639e-07, 7.60144e-06, 9.532007e-06, 9.076497e-06, 5.391629e-06,
  3.977326e-06, 3.68691e-06, 4.252683e-05, 9.418633e-05, 5.057058e-05, 
    1.609822e-05, 5.669522e-06, 4.571248e-06, 3.663108e-06, 3.283747e-06, 
    8.955937e-07, 8.953618e-06, 9.267427e-06, 8.30625e-06, 6.133222e-06,
  2.709407e-08, 5.707263e-06, 1.996823e-05, 4.304051e-05, 1.581247e-05, 
    6.148317e-06, 1.792555e-05, 7.524552e-05, 0.0001175657, 7.458196e-05, 
    3.626676e-05, 9.09651e-06, 2.668482e-07, 4.194442e-07, 9.577374e-07,
  2.672546e-08, 7.388853e-06, 2.158389e-05, 3.94638e-05, 1.909203e-05, 
    2.608634e-05, 5.631389e-05, 9.750679e-05, 9.739656e-05, 4.461916e-05, 
    4.473131e-06, 2.568505e-07, 3.361181e-07, 2.610563e-06, 2.749923e-06,
  4.456937e-06, 6.488205e-06, 2.101943e-05, 3.895192e-05, 1.905128e-05, 
    6.253172e-05, 5.472432e-05, 8.132857e-05, 5.836913e-05, 4.611938e-06, 
    2.665099e-06, 2.719208e-06, 2.279485e-06, 1.832857e-06, 3.182735e-06,
  3.041193e-05, 6.161588e-06, 2.09732e-05, 1.300168e-05, 1.98526e-05, 
    3.394877e-06, 6.910937e-05, 1.647119e-05, 7.409469e-06, 5.596525e-06, 
    4.891426e-06, 3.260811e-06, 4.157535e-06, 3.975068e-06, 2.278987e-06,
  2.726382e-05, 2.711719e-06, 3.930186e-05, 4.549335e-06, 7.098208e-06, 
    9.903423e-06, 5.286007e-07, 1.0193e-06, 8.339989e-06, 4.339629e-06, 
    6.064787e-06, 4.680501e-06, 4.380373e-06, 2.080521e-06, 1.70863e-06,
  9.539825e-06, 2.176303e-06, 4.548305e-05, 7.467915e-06, 1.147061e-06, 
    4.782435e-06, 1.745004e-06, 1.36864e-06, 3.439388e-07, 4.712746e-06, 
    4.601749e-06, 4.439773e-06, 4.071372e-06, 3.316056e-06, 3.312366e-06,
  3.410795e-06, 1.854827e-06, 5.005777e-05, 1.551557e-05, 2.653333e-06, 
    4.656818e-06, 8.030849e-07, 2.609175e-06, 3.559623e-06, 3.777202e-06, 
    3.559202e-06, 3.556532e-06, 3.686333e-06, 3.284482e-06, 4.713856e-06,
  2.884949e-06, 1.641682e-06, 6.546518e-05, 3.10784e-05, 1.326998e-05, 
    1.060352e-05, 1.860985e-06, 1.751783e-06, 2.725848e-06, 3.587703e-06, 
    2.929371e-06, 4.772606e-06, 5.790781e-06, 5.438678e-06, 5.993681e-06,
  2.377726e-06, 1.704202e-06, 7.466268e-05, 7.051629e-05, 3.358272e-05, 
    2.185132e-05, 4.951018e-06, 3.502187e-06, 3.376852e-06, 4.797446e-06, 
    3.834832e-06, 4.255941e-06, 6.173607e-06, 5.98583e-06, 5.320979e-06,
  2.31764e-06, 3.414581e-06, 7.942537e-05, 0.0001106023, 5.585309e-05, 
    3.464794e-05, 1.268793e-05, 3.516681e-06, 2.928283e-06, 5.200527e-06, 
    7.004304e-06, 5.638472e-06, 5.620592e-06, 6.285713e-06, 6.598602e-06,
  6.173373e-06, 4.783639e-06, 3.440523e-05, 3.610761e-05, 1.320031e-05, 
    6.059841e-06, 6.831408e-06, 9.384058e-06, 5.944439e-06, 3.112352e-06, 
    2.995144e-06, 2.082507e-06, 1.976699e-06, 2.497237e-06, 1.5054e-06,
  2.470741e-05, 2.725163e-05, 5.102103e-05, 4.495131e-05, 1.57972e-05, 
    7.915215e-06, 6.724986e-06, 5.322236e-06, 1.353809e-06, 2.706013e-06, 
    3.294711e-06, 1.604045e-06, 6.37682e-07, 1.039368e-06, 2.255576e-06,
  0.0001047949, 6.132588e-05, 5.034842e-05, 4.112595e-05, 1.694267e-05, 
    2.837889e-05, 1.192108e-05, 5.38664e-06, 4.062617e-06, 2.505079e-06, 
    1.173095e-06, 5.937964e-07, 1.057231e-06, 1.087775e-06, 1.395005e-06,
  0.0001311233, 7.074752e-05, 4.866217e-05, 3.515026e-05, 3.117603e-05, 
    7.168722e-06, 3.41303e-05, 9.676643e-06, 6.962214e-06, 4.4345e-06, 
    2.881885e-06, 2.145651e-06, 1.101977e-06, 1.221791e-06, 2.599689e-06,
  0.0001101728, 8.204015e-05, 6.319572e-05, 4.154263e-05, 3.827765e-05, 
    3.558964e-05, 8.708283e-06, 6.788286e-06, 6.060187e-06, 3.847761e-06, 
    5.937317e-06, 2.549769e-06, 3.863887e-06, 4.980689e-06, 3.949971e-06,
  8.439962e-05, 7.352493e-05, 6.005052e-05, 4.678681e-05, 4.276112e-05, 
    4.661302e-05, 2.934239e-05, 8.302558e-07, 6.631209e-07, 6.550931e-06, 
    4.548865e-06, 4.344083e-06, 3.993498e-06, 4.181179e-06, 5.459651e-06,
  8.239935e-05, 7.791026e-05, 7.254394e-05, 7.205083e-05, 6.876957e-05, 
    5.914621e-05, 4.182504e-05, 1.136193e-05, 4.679386e-06, 7.162048e-06, 
    4.309424e-06, 4.535932e-06, 3.049297e-06, 2.809288e-06, 5.099508e-06,
  0.0001013861, 0.0001090557, 0.0001181682, 0.0001203567, 0.0001038697, 
    7.91382e-05, 3.660339e-05, 9.959997e-06, 6.632161e-06, 7.267229e-06, 
    4.015164e-06, 4.193443e-06, 4.174119e-06, 5.92457e-06, 5.085889e-06,
  9.183311e-05, 0.0001057912, 0.0001512452, 0.0001770577, 0.0001404901, 
    7.414663e-05, 2.701628e-05, 7.992846e-06, 9.044874e-06, 7.279265e-06, 
    4.295306e-06, 3.785088e-06, 5.678671e-06, 5.542453e-06, 4.072953e-06,
  7.738436e-05, 9.58516e-05, 0.0001657027, 0.000198335, 0.0001450121, 
    6.062534e-05, 1.773434e-05, 8.040258e-06, 1.004507e-05, 5.919314e-06, 
    5.182443e-06, 5.548916e-06, 6.262648e-06, 6.344531e-06, 7.938707e-06,
  8.106342e-05, 5.043065e-05, 4.762126e-05, 4.889701e-05, 2.846042e-05, 
    1.698882e-05, 1.079923e-05, 1.159384e-05, 1.398122e-05, 1.090507e-05, 
    6.347475e-06, 5.484216e-06, 7.784164e-06, 8.300276e-06, 5.333437e-06,
  0.0001323275, 0.0001068078, 9.989813e-05, 7.896017e-05, 4.07296e-05, 
    1.110437e-05, 1.371413e-05, 1.137611e-05, 1.32332e-05, 2.079007e-05, 
    1.724176e-05, 7.743224e-06, 5.440074e-06, 2.367651e-06, 3.583237e-06,
  0.0001069144, 7.972173e-05, 5.628862e-05, 3.11604e-05, 1.273031e-05, 
    1.500079e-05, 1.111029e-05, 3.458604e-05, 2.356902e-05, 2.380088e-05, 
    2.022942e-05, 1.410325e-05, 5.348613e-06, 3.59162e-06, 4.022064e-06,
  4.724999e-05, 1.422996e-05, 5.81683e-06, 4.001076e-06, 4.894605e-06, 
    7.297007e-06, 3.035312e-05, 3.862141e-05, 3.204144e-05, 3.261615e-05, 
    3.069348e-05, 2.195755e-05, 1.069742e-05, 5.234617e-06, 3.602605e-06,
  2.037526e-06, 1.656096e-06, 1.39468e-06, 2.123004e-06, 3.508791e-06, 
    1.112393e-05, 1.948985e-05, 4.791009e-05, 2.986778e-05, 3.957266e-05, 
    4.489045e-05, 2.813027e-05, 1.237552e-05, 6.852018e-06, 5.812761e-06,
  3.340918e-07, 2.381915e-07, 1.280915e-07, 3.597199e-07, 1.233044e-06, 
    6.469271e-06, 2.454398e-05, 2.909916e-05, 2.306407e-05, 4.987634e-05, 
    3.63613e-05, 2.824672e-05, 1.654923e-05, 9.312451e-06, 5.160993e-06,
  1.689221e-07, 5.395545e-09, 1.811449e-07, 7.676675e-07, 3.974877e-06, 
    7.866285e-06, 2.578349e-05, 5.946639e-05, 5.49094e-05, 4.170472e-05, 
    3.264385e-05, 3.199396e-05, 1.617818e-05, 8.352903e-06, 5.157142e-06,
  3.193998e-07, 2.281513e-07, 8.374851e-07, 4.564908e-06, 7.520713e-06, 
    1.202709e-05, 3.085612e-05, 4.565046e-05, 3.524598e-05, 3.504802e-05, 
    3.708022e-05, 3.505298e-05, 1.493833e-05, 6.992681e-06, 5.032644e-06,
  1.632532e-06, 8.298836e-07, 5.394475e-06, 7.944098e-06, 1.220594e-05, 
    3.063892e-05, 4.549322e-05, 5.287751e-05, 4.500811e-05, 4.129663e-05, 
    3.706639e-05, 2.693567e-05, 1.1716e-05, 6.350873e-06, 4.365369e-06,
  1.884061e-07, 2.105094e-06, 4.225267e-05, 5.717297e-05, 4.785026e-05, 
    5.49584e-05, 5.49488e-05, 4.993537e-05, 4.047313e-05, 3.477364e-05, 
    2.877654e-05, 1.681646e-05, 6.564568e-06, 2.596992e-06, 1.371531e-06,
  4.946742e-05, 2.748588e-05, 1.891292e-05, 4.088505e-05, 8.894761e-05, 
    0.0001303004, 0.0001605006, 0.0001865876, 0.0001918969, 0.0001737485, 
    0.0001485556, 0.0001281684, 0.0001067343, 6.9815e-05, 1.889831e-05,
  0.0002939305, 0.0002468555, 0.0002007448, 0.000199407, 0.0001882382, 
    0.0001713263, 0.0001091593, 5.560452e-05, 2.90376e-05, 2.966675e-05, 
    2.672828e-05, 3.191287e-05, 3.908796e-05, 3.97701e-05, 1.366501e-05,
  0.0003382408, 0.0002966511, 0.0002558414, 0.0002040488, 0.0001144879, 
    5.244252e-05, 1.403227e-05, 6.608504e-06, 3.926149e-06, 4.063079e-06, 
    4.430528e-06, 8.607247e-06, 1.741773e-05, 2.130755e-05, 1.637181e-05,
  0.0002105539, 0.0001900147, 0.0001446507, 8.237961e-05, 2.372291e-05, 
    2.97477e-06, 2.30912e-06, 2.438522e-06, 8.420415e-07, 3.945929e-06, 
    4.095562e-06, 8.401155e-06, 1.678075e-05, 2.039959e-05, 2.165539e-05,
  2.771424e-05, 2.097184e-05, 1.297812e-05, 6.760443e-06, 4.352262e-06, 
    5.440804e-06, 3.848804e-06, 3.180863e-06, 1.568267e-06, 3.66239e-07, 
    2.972267e-06, 9.260754e-06, 2.034335e-05, 2.047599e-05, 2.284881e-05,
  4.650096e-06, 4.467095e-06, 2.860265e-06, 2.688545e-06, 4.26875e-06, 
    5.584617e-06, 8.420006e-06, 3.370052e-06, 1.870766e-06, 2.701039e-06, 
    4.065597e-06, 8.243637e-06, 1.969788e-05, 2.087834e-05, 1.952924e-05,
  3.57055e-06, 5.032567e-06, 4.577975e-06, 3.041315e-06, 4.087425e-06, 
    4.952666e-06, 5.531354e-06, 8.532677e-06, 1.09883e-05, 6.644395e-06, 
    4.141948e-06, 7.411052e-06, 1.649797e-05, 1.895092e-05, 1.200176e-05,
  4.422766e-06, 5.81235e-06, 6.502257e-06, 5.447669e-06, 2.744794e-06, 
    3.045798e-06, 8.937664e-06, 2.534161e-05, 2.868591e-05, 2.920906e-05, 
    2.074456e-05, 1.069106e-05, 1.925584e-05, 1.988547e-05, 1.105813e-05,
  5.618391e-06, 3.152634e-06, 2.613845e-06, 2.245689e-06, 5.747503e-06, 
    5.847646e-06, 1.835533e-05, 3.09588e-05, 3.663174e-05, 4.171679e-05, 
    3.467384e-05, 2.072148e-05, 2.577609e-05, 2.528816e-05, 1.086984e-05,
  3.765324e-06, 3.762976e-06, 2.103256e-06, 3.669016e-06, 4.913247e-06, 
    4.992665e-06, 9.695449e-06, 1.24199e-05, 1.775689e-05, 2.013382e-05, 
    1.8748e-05, 2.085981e-05, 2.467438e-05, 1.911841e-05, 1.431613e-05,
  4.137768e-07, 8.603013e-07, 6.479875e-07, 2.842469e-06, 2.630467e-06, 
    2.494636e-06, 5.618427e-06, 1.231248e-05, 2.664713e-05, 2.348684e-05, 
    2.159283e-05, 2.035031e-05, 1.875299e-05, 3.340933e-05, 6.477744e-05,
  1.113073e-05, 6.463021e-06, 6.236363e-06, 1.152875e-05, 3.675618e-05, 
    6.250764e-05, 7.996574e-05, 9.458941e-05, 0.0001018119, 9.912252e-05, 
    9.374091e-05, 9.641955e-05, 8.282917e-05, 8.981829e-05, 9.578004e-05,
  9.844197e-05, 8.950161e-05, 6.913004e-05, 8.058715e-05, 0.0001324312, 
    0.0001778564, 0.0001754605, 0.0001615509, 0.000157529, 0.000159734, 
    0.0001478783, 0.0001301626, 0.0001173198, 0.0001018688, 0.0001205608,
  0.0001459567, 0.0001951866, 0.0001909095, 0.0001836673, 0.0001914191, 
    0.0001436942, 0.0001805015, 0.0001676433, 0.00013523, 0.0001156476, 
    9.799752e-05, 7.459956e-05, 6.833801e-05, 7.365737e-05, 8.411792e-05,
  6.549548e-05, 0.0001078801, 0.0001222138, 0.0001003681, 9.47441e-05, 
    0.000104617, 5.898853e-05, 7.02547e-05, 0.0001399298, 0.0001204871, 
    8.83414e-05, 6.334551e-05, 4.012885e-05, 3.370461e-05, 3.893817e-05,
  1.275258e-05, 1.919025e-05, 2.44829e-05, 2.578673e-05, 2.040225e-05, 
    1.930484e-05, 1.928208e-05, 4.127424e-05, 5.066923e-05, 3.635948e-05, 
    2.62764e-05, 1.43103e-05, 8.887157e-06, 9.695143e-06, 1.365529e-05,
  6.569357e-06, 9.221552e-06, 4.806639e-06, 4.967509e-06, 4.702216e-06, 
    4.841904e-06, 4.015899e-06, 6.92914e-06, 1.169126e-05, 1.070982e-05, 
    8.034664e-06, 5.810272e-06, 5.381275e-06, 6.288982e-06, 1.128975e-05,
  6.152326e-06, 5.715471e-06, 3.206276e-06, 3.18522e-06, 2.053019e-06, 
    4.976106e-06, 4.646276e-06, 3.756636e-06, 3.487228e-06, 5.428966e-06, 
    6.919101e-06, 5.48077e-06, 5.077287e-06, 9.093308e-06, 1.023026e-05,
  7.833988e-06, 2.013917e-06, 2.255937e-06, 4.750069e-06, 3.646955e-06, 
    3.434919e-06, 4.63988e-06, 5.654545e-06, 5.117258e-06, 4.497586e-06, 
    5.708629e-06, 7.209864e-06, 5.879091e-06, 1.128349e-05, 7.950074e-06,
  6.786358e-06, 1.536359e-06, 1.198545e-06, 4.406839e-06, 4.703102e-06, 
    3.796576e-06, 5.767257e-06, 8.438149e-06, 7.712628e-06, 4.77482e-06, 
    5.531161e-06, 5.586976e-06, 5.512582e-06, 4.880228e-06, 4.723136e-06,
  0.000384161, 0.0001901183, 6.929762e-05, 3.406258e-05, 1.776729e-05, 
    1.019573e-05, 1.399835e-06, 1.900097e-08, 1.308973e-07, 9.681722e-07, 
    2.520936e-06, 2.728149e-06, 5.863787e-06, 1.886106e-05, 1.229915e-05,
  0.0003003632, 0.0002811599, 0.0001777928, 9.287971e-05, 2.983528e-05, 
    6.899572e-06, 1.62108e-07, 1.28451e-08, 1.153254e-07, 3.119427e-07, 
    1.211596e-06, 4.279444e-06, 1.098475e-05, 3.655463e-05, 2.010872e-05,
  0.0001262678, 0.000141637, 9.957921e-05, 4.86391e-05, 1.154197e-05, 
    5.994822e-06, 7.602474e-07, 7.666343e-08, 5.104543e-07, 7.957319e-07, 
    1.75128e-06, 6.795833e-06, 1.253357e-05, 2.071067e-05, 2.483386e-05,
  6.82537e-06, 9.864296e-06, 9.450957e-06, 4.849647e-06, 1.4395e-06, 
    1.831993e-06, 1.549016e-05, 4.465361e-07, 7.968052e-07, 3.306748e-06, 
    6.057935e-06, 7.421292e-06, 8.161213e-06, 1.1893e-05, 2.055197e-05,
  2.576198e-06, 3.353693e-06, 3.661235e-06, 2.636621e-06, 2.661968e-06, 
    1.782414e-06, 2.43734e-06, 8.692353e-06, 1.472236e-05, 9.136469e-06, 
    1.731411e-05, 1.724035e-05, 1.335489e-05, 1.613071e-05, 3.25145e-05,
  3.805676e-06, 3.247841e-06, 3.713739e-06, 2.117585e-06, 1.551752e-06, 
    2.051031e-06, 3.609546e-06, 4.549301e-06, 5.479133e-06, 7.405362e-06, 
    2.006565e-05, 3.382065e-05, 4.397351e-05, 5.186226e-05, 6.175668e-05,
  5.527605e-06, 3.710242e-06, 2.586114e-06, 2.85858e-06, 4.194448e-06, 
    4.462929e-06, 5.780243e-06, 4.704702e-06, 5.295444e-06, 8.391251e-06, 
    1.640815e-05, 2.156228e-05, 4.204553e-05, 5.391487e-05, 3.800068e-05,
  6.34721e-06, 2.863738e-06, 2.211409e-06, 5.369318e-06, 4.816938e-06, 
    4.95099e-06, 3.495485e-06, 4.033541e-06, 6.494188e-06, 8.726352e-06, 
    1.611563e-05, 1.404014e-05, 2.238565e-05, 2.351768e-05, 1.736638e-05,
  6.080586e-06, 1.747996e-06, 2.117109e-06, 7.026777e-06, 4.537689e-06, 
    6.014006e-06, 3.918153e-06, 2.768318e-06, 3.099628e-06, 4.148657e-06, 
    1.146003e-05, 1.391573e-05, 1.233312e-05, 1.280622e-05, 7.653259e-06,
  2.300719e-06, 2.434293e-06, 3.74928e-06, 3.279286e-06, 3.233303e-06, 
    3.03204e-06, 3.158003e-06, 2.307919e-06, 3.501487e-06, 1.447525e-06, 
    9.054722e-06, 1.154502e-05, 5.964357e-06, 6.118541e-06, 5.991289e-06,
  1.18644e-05, 4.500873e-06, 2.115623e-06, 5.630082e-06, 9.209676e-07, 
    3.38927e-06, 1.239014e-05, 1.024726e-05, 6.752086e-06, 5.091524e-06, 
    5.514629e-06, 5.080251e-06, 5.249619e-06, 3.013818e-06, 3.958578e-06,
  9.541825e-05, 8.549583e-05, 6.264204e-05, 5.441114e-05, 3.680338e-05, 
    3.4434e-05, 2.834329e-05, 2.306508e-05, 2.142669e-05, 2.267187e-05, 
    1.904234e-05, 1.364263e-05, 5.415781e-06, 5.842224e-06, 5.800077e-06,
  0.0001752641, 0.0001970042, 0.0002001279, 0.0001888102, 0.0001288289, 
    0.0001392783, 9.410972e-05, 5.654791e-05, 4.051752e-05, 3.434722e-05, 
    2.213718e-05, 1.253016e-05, 3.928658e-06, 4.341863e-06, 5.466675e-06,
  0.0001052766, 0.0001752743, 0.0001966651, 0.0001883942, 0.0001725992, 
    9.804912e-05, 0.0001377881, 0.000106635, 7.420794e-05, 4.721642e-05, 
    3.601947e-05, 1.529277e-05, 7.233553e-06, 3.023192e-06, 5.952856e-06,
  2.138256e-05, 5.332571e-05, 8.498751e-05, 8.84553e-05, 0.0001039815, 
    0.0001169445, 4.857585e-05, 8.674481e-05, 9.254582e-05, 4.249943e-05, 
    3.414778e-05, 8.379499e-06, 4.85093e-06, 3.960371e-06, 9.287319e-06,
  4.916831e-06, 9.943153e-06, 2.265314e-05, 3.637608e-05, 3.984183e-05, 
    5.578074e-05, 6.009778e-05, 1.81637e-05, 1.036329e-05, 1.553456e-05, 
    8.131494e-06, 2.45567e-06, 2.804434e-06, 9.160167e-06, 1.661879e-05,
  6.019722e-06, 3.073661e-06, 4.340307e-06, 9.103918e-06, 1.386751e-05, 
    1.686234e-05, 2.493563e-05, 3.19419e-05, 1.944754e-05, 8.76488e-06, 
    5.364449e-06, 4.097878e-07, 1.60991e-06, 1.192919e-05, 1.828211e-05,
  5.063775e-06, 3.45053e-06, 1.226641e-06, 2.932715e-06, 4.916266e-06, 
    5.961322e-06, 5.790323e-06, 6.055016e-06, 5.895786e-06, 4.461036e-06, 
    3.177753e-06, 2.114682e-06, 1.383295e-06, 1.092883e-05, 1.37237e-05,
  7.977015e-06, 1.713918e-06, 1.764497e-06, 2.872031e-06, 2.381674e-06, 
    2.639339e-06, 3.558544e-06, 4.355642e-06, 3.865506e-06, 4.147666e-06, 
    3.555106e-06, 3.167919e-06, 1.637408e-06, 1.020444e-05, 1.376132e-05,
  1.973403e-06, 2.024517e-06, 2.373569e-06, 1.623738e-06, 2.144936e-06, 
    1.59362e-06, 4.500351e-06, 3.460634e-06, 3.308527e-07, 4.296347e-06, 
    3.84631e-06, 4.420938e-06, 6.859859e-06, 1.328109e-05, 1.110465e-05,
  2.752676e-06, 1.917036e-06, 1.506785e-05, 7.631961e-05, 1.61785e-05, 
    2.885268e-07, 7.065025e-06, 3.366434e-06, 8.688731e-06, 8.600147e-08, 
    5.165208e-08, 1.101368e-07, 2.118275e-07, 1.240865e-06, 9.677915e-07,
  5.275477e-06, 4.872217e-06, 2.587371e-06, 1.582906e-05, 2.627115e-05, 
    1.302849e-06, 2.606661e-06, 3.075169e-06, 2.808893e-06, 7.070432e-06, 
    1.333611e-07, 7.847387e-07, 1.683622e-06, 3.551018e-06, 1.042632e-06,
  5.297663e-06, 5.2241e-06, 3.960506e-06, 4.457403e-06, 4.291802e-06, 
    7.301289e-06, 2.901123e-06, 9.852087e-07, 3.252471e-06, 6.49703e-06, 
    9.164423e-06, 2.532432e-06, 8.049217e-06, 1.891574e-06, 5.696456e-06,
  4.377638e-06, 6.726222e-06, 7.338283e-06, 4.816916e-06, 8.95845e-06, 
    2.978046e-06, 9.049431e-06, 4.76029e-06, 2.627898e-06, 2.388377e-06, 
    5.218104e-06, 9.300384e-06, 9.731486e-06, 3.253531e-06, 1.457612e-05,
  6.136221e-06, 8.13306e-06, 9.86964e-06, 1.438785e-05, 1.121553e-05, 
    6.913699e-06, 5.0876e-06, 2.639229e-05, 2.710314e-05, 1.076152e-05, 
    2.439907e-05, 1.723778e-05, 1.328058e-05, 1.884859e-05, 4.646628e-05,
  6.70829e-06, 5.427326e-06, 9.168781e-06, 1.779031e-05, 1.81136e-05, 
    2.183073e-05, 3.581342e-05, 7.987302e-06, 6.410161e-06, 6.783618e-05, 
    6.572807e-05, 4.295797e-05, 6.420945e-05, 7.404913e-05, 8.637822e-05,
  9.410211e-06, 4.816217e-06, 3.695424e-06, 1.999555e-05, 1.97123e-05, 
    2.168477e-05, 3.716182e-05, 9.265346e-05, 0.0001439404, 0.0001222752, 
    9.450957e-05, 9.362733e-05, 0.000105168, 0.0001014653, 6.460346e-05,
  8.527129e-06, 4.711717e-06, 3.497023e-06, 6.231729e-06, 1.468894e-05, 
    2.019077e-05, 2.406631e-05, 4.432288e-05, 9.046667e-05, 9.787574e-05, 
    8.942954e-05, 8.081026e-05, 7.993801e-05, 6.536092e-05, 2.083464e-05,
  2.830758e-06, 2.9612e-06, 3.677819e-06, 3.842774e-06, 1.250806e-05, 
    2.505797e-05, 5.080365e-05, 8.305164e-05, 0.0001056214, 0.0001019166, 
    7.643614e-05, 5.929258e-05, 5.039621e-05, 2.692704e-05, 5.136287e-06,
  2.14831e-06, 2.231518e-06, 4.330397e-06, 4.228681e-06, 1.304368e-05, 
    3.836955e-05, 6.440593e-05, 8.91584e-05, 9.022309e-05, 7.287315e-05, 
    6.034249e-05, 4.731334e-05, 3.119857e-05, 1.212358e-05, 5.012777e-06,
  5.918642e-05, 8.614919e-05, 9.851828e-05, 6.610613e-05, 7.146527e-06, 
    1.737335e-06, 7.460935e-06, 8.957199e-06, 1.15206e-05, 1.422903e-07, 
    2.802864e-07, 4.959377e-09, 1.741172e-08, 9.210027e-08, 5.160717e-07,
  2.878695e-05, 2.075289e-05, 2.278368e-05, 7.003683e-05, 5.767717e-05, 
    1.372465e-06, 3.191523e-06, 5.020219e-06, 6.405707e-06, 1.020191e-05, 
    4.566939e-07, 1.170736e-06, 1.49224e-06, 9.069252e-08, 1.749162e-06,
  6.398904e-06, 8.096235e-06, 4.363558e-06, 9.780828e-06, 5.328346e-05, 
    5.936528e-05, 6.598023e-07, 5.5015e-06, 6.22895e-06, 1.076447e-05, 
    1.279941e-05, 8.361322e-06, 8.516244e-06, 1.002128e-06, 1.061028e-07,
  4.308263e-06, 4.682963e-06, 2.379824e-06, 2.963473e-06, 2.481427e-06, 
    3.02626e-05, 3.688321e-05, 1.759583e-06, 2.928952e-06, 8.395467e-06, 
    1.20118e-05, 1.337296e-05, 5.966037e-06, 3.699069e-06, 9.797969e-08,
  1.700078e-06, 5.318815e-06, 2.732038e-06, 1.581243e-06, 2.857618e-06, 
    1.887031e-06, 1.459132e-05, 1.911064e-05, 1.106923e-05, 3.380178e-06, 
    6.311506e-06, 9.736894e-06, 1.187874e-05, 4.049289e-06, 1.315153e-06,
  1.174463e-06, 5.423818e-06, 3.104041e-06, 1.403106e-06, 3.338268e-06, 
    2.7401e-06, 2.363208e-06, 2.891863e-06, 1.627768e-06, 8.178349e-07, 
    3.047774e-06, 7.124852e-06, 7.174e-06, 6.541105e-06, 4.564696e-06,
  2.033298e-06, 3.992001e-06, 4.232915e-06, 1.155657e-06, 2.507601e-06, 
    3.661428e-06, 2.310895e-06, 1.406115e-06, 2.951982e-06, 2.29098e-06, 
    1.560806e-06, 1.303401e-06, 2.830177e-06, 4.164892e-06, 2.106685e-05,
  1.678019e-06, 2.569211e-06, 4.624319e-06, 1.532989e-06, 3.048266e-06, 
    3.639355e-06, 2.079136e-06, 2.048776e-06, 1.498535e-06, 1.234602e-06, 
    2.254108e-06, 2.764638e-06, 3.569952e-06, 1.195628e-05, 4.436642e-05,
  2.623695e-06, 2.362427e-06, 5.4351e-06, 9.540685e-07, 2.848915e-06, 
    3.866e-06, 2.783515e-06, 3.863993e-06, 7.318364e-06, 3.932028e-06, 
    3.614686e-06, 4.500136e-06, 1.383594e-05, 4.079557e-05, 4.997733e-05,
  2.11246e-06, 2.184241e-06, 3.201791e-06, 2.239081e-06, 2.956437e-06, 
    3.262216e-06, 6.042126e-06, 8.276013e-06, 1.160978e-05, 8.011248e-06, 
    9.663162e-06, 1.736636e-05, 3.627808e-05, 5.494072e-05, 5.372731e-05,
  0.0005030062, 0.0001558666, 5.775887e-05, 6.341383e-06, 5.583871e-06, 
    4.38295e-06, 6.374818e-06, 4.484948e-06, 5.57471e-06, 1.547525e-07, 
    2.630606e-08, 2.747471e-09, 3.700864e-07, 1.894648e-08, 2.665784e-07,
  0.0004493719, 0.00025492, 0.0001351986, 7.365417e-05, 1.000751e-05, 
    3.18993e-06, 3.799345e-06, 3.348254e-06, 9.396372e-06, 1.604937e-05, 
    1.481096e-06, 1.420596e-05, 1.483858e-05, 5.879825e-07, 1.982397e-07,
  0.0002491354, 0.0003036468, 0.0001753387, 0.000133376, 3.976267e-05, 
    1.974126e-05, 5.917193e-06, 8.364481e-06, 7.003922e-06, 1.239781e-05, 
    1.4027e-05, 1.080457e-05, 1.317407e-05, 9.714905e-06, 2.932764e-07,
  7.047668e-05, 0.0001709874, 0.0002070343, 0.0001429371, 0.0001091089, 
    2.248178e-05, 3.305396e-05, 6.61881e-06, 5.348347e-06, 9.172345e-06, 
    6.634879e-06, 9.672035e-06, 9.818003e-06, 1.36906e-05, 1.321491e-05,
  8.353342e-06, 4.539646e-05, 0.0001201523, 0.0001429017, 0.0001271873, 
    0.000117857, 1.185888e-05, 1.776133e-05, 1.972553e-05, 4.659362e-06, 
    4.835405e-06, 5.761331e-06, 8.051049e-06, 9.992542e-06, 1.626352e-05,
  8.055529e-07, 6.446124e-06, 2.824721e-05, 7.930391e-05, 0.0001163647, 
    0.0001216886, 0.0001158023, 3.694814e-06, 9.695235e-07, 1.038541e-06, 
    1.432517e-06, 2.049062e-06, 4.635258e-06, 6.905907e-06, 1.028011e-05,
  1.022065e-07, 8.119676e-07, 4.326796e-06, 1.60264e-05, 5.325566e-05, 
    8.76809e-05, 0.0001068124, 0.0001109356, 4.167564e-05, 4.378237e-06, 
    1.680563e-06, 4.535127e-07, 7.748412e-07, 4.268693e-06, 5.766542e-06,
  3.376393e-07, 6.828632e-08, 4.871071e-07, 4.433698e-06, 1.253026e-05, 
    4.281037e-05, 7.014209e-05, 5.848556e-05, 3.93087e-05, 2.40214e-05, 
    9.709534e-06, 1.01229e-06, 1.914175e-07, 2.766826e-07, 1.11813e-06,
  1.862482e-06, 2.118187e-08, 2.778557e-06, 3.037838e-06, 4.317501e-06, 
    7.581244e-06, 1.911152e-05, 4.287743e-05, 4.814212e-05, 3.213134e-05, 
    1.097476e-05, 1.215158e-06, 7.406776e-07, 4.237284e-07, 4.72889e-07,
  2.279471e-07, 8.902628e-08, 2.292859e-07, 3.238455e-06, 2.732606e-06, 
    4.144564e-06, 4.583095e-06, 5.953108e-06, 1.24029e-05, 1.513995e-05, 
    9.794424e-06, 3.800723e-06, 1.701842e-06, 1.23723e-06, 1.098469e-06,
  5.315629e-05, 1.778166e-05, 1.324532e-06, 1.179163e-08, 6.36063e-09, 
    1.635117e-05, 4.699533e-05, 1.100923e-05, 1.165822e-05, 1.787551e-07, 
    5.648144e-08, 7.116004e-11, 3.420546e-08, 1.240077e-08, 3.890361e-10,
  8.622507e-05, 2.014183e-05, 3.177331e-06, 2.624371e-08, 5.578366e-08, 
    1.295059e-05, 4.805432e-05, 1.80147e-05, 3.717415e-06, 2.073072e-05, 
    2.167061e-07, 1.016231e-05, 2.047964e-06, 1.913458e-08, 8.355717e-09,
  0.0001685021, 6.546926e-05, 7.914487e-06, 1.923991e-07, 1.002157e-07, 
    3.054795e-05, 5.475919e-05, 3.640288e-05, 2.678906e-06, 7.765671e-06, 
    1.565345e-05, 2.35146e-06, 2.72435e-06, 8.976797e-06, 1.660945e-08,
  0.0001896875, 0.0001524061, 5.028877e-05, 1.687033e-06, 2.732199e-07, 
    9.276078e-06, 6.957883e-05, 5.769591e-05, 3.533307e-06, 1.025557e-05, 
    5.951209e-06, 6.229978e-06, 5.902653e-06, 7.470656e-06, 1.402716e-05,
  8.116505e-05, 0.0001750793, 0.0001377715, 4.924429e-05, 1.272972e-05, 
    4.665556e-05, 1.033753e-05, 7.252801e-05, 2.05009e-05, 5.65872e-06, 
    1.311672e-05, 8.840202e-06, 6.221465e-06, 1.173791e-05, 1.605813e-05,
  2.342481e-05, 0.0001016399, 0.0001505653, 0.0001275743, 9.64938e-05, 
    5.405631e-05, 2.437443e-05, 2.000268e-05, 1.896261e-06, 4.661332e-06, 
    6.753272e-06, 6.264058e-06, 6.320614e-06, 6.255615e-06, 1.007467e-05,
  5.057602e-07, 2.184147e-05, 8.199342e-05, 0.0001445798, 0.0001565742, 
    8.962808e-05, 2.716684e-05, 6.36297e-05, 1.839108e-05, 4.79889e-06, 
    6.126572e-06, 5.11755e-06, 4.263494e-06, 5.268809e-06, 5.94133e-06,
  1.216105e-06, 5.777878e-06, 2.045435e-05, 7.869246e-05, 0.0001439636, 
    0.0001525985, 6.221713e-05, 2.239099e-05, 1.519092e-05, 5.917581e-06, 
    4.037255e-06, 4.553749e-06, 3.455888e-06, 4.475103e-06, 5.124519e-06,
  1.631368e-06, 9.947665e-07, 5.432198e-06, 1.973142e-05, 7.635118e-05, 
    0.0001446078, 0.0001624199, 0.0001102682, 5.798394e-05, 2.474498e-05, 
    1.785689e-05, 9.093082e-06, 4.017948e-06, 3.232326e-06, 4.59913e-06,
  7.578137e-07, 2.19984e-07, 1.600646e-06, 4.513123e-06, 1.693958e-05, 
    7.812857e-05, 0.0001318391, 0.0001398519, 0.0001123476, 7.780647e-05, 
    4.195979e-05, 1.4858e-05, 6.406699e-06, 3.874874e-06, 2.855839e-06,
  8.068814e-05, 2.963968e-05, 1.820964e-06, 5.70356e-07, 2.045339e-08, 
    8.76278e-08, 1.229898e-05, 0.0001326726, 2.002453e-05, 6.19449e-06, 
    1.092543e-08, 2.052598e-25, 3.010437e-12, 1.507175e-11, 7.119658e-11,
  8.162703e-05, 3.0103e-05, 7.165615e-06, 1.037402e-06, 2.323887e-07, 
    4.030123e-08, 1.5166e-05, 0.0001191901, 8.294125e-06, 1.287781e-05, 
    1.708833e-08, 2.766468e-10, 1.03674e-13, 6.998988e-12, 3.205724e-11,
  7.883955e-05, 3.80027e-05, 1.294483e-05, 2.342473e-06, 6.228877e-07, 
    2.474731e-07, 2.236015e-05, 0.0001248187, 5.313088e-06, 1.227313e-05, 
    1.972305e-06, 8.778837e-09, 9.282866e-07, 1.341207e-05, 9.66413e-11,
  5.04971e-05, 5.122949e-05, 1.452738e-05, 5.788771e-06, 3.582131e-07, 
    3.680166e-08, 3.989632e-05, 8.215888e-05, 5.845768e-06, 7.975137e-06, 
    2.333134e-06, 1.502779e-06, 4.964587e-06, 8.244678e-06, 4.879592e-06,
  3.182319e-05, 7.35093e-05, 2.741939e-05, 7.632856e-06, 1.326191e-06, 
    8.487547e-07, 2.538579e-05, 6.642153e-05, 1.755342e-05, 5.814923e-06, 
    5.185285e-06, 2.095352e-06, 3.853183e-06, 9.281107e-06, 1.343942e-05,
  1.830383e-05, 4.978305e-05, 4.872248e-05, 1.883002e-05, 2.050396e-05, 
    6.151563e-06, 1.133316e-05, 2.220876e-05, 8.828348e-07, 5.99643e-06, 
    7.000584e-06, 2.047917e-06, 5.36843e-06, 2.780647e-06, 5.299942e-06,
  2.882669e-06, 2.407962e-05, 4.559908e-05, 4.365638e-05, 8.079599e-05, 
    5.08943e-05, 1.211001e-05, 1.350057e-05, 2.373962e-06, 5.897387e-06, 
    9.509585e-06, 1.371807e-06, 3.307807e-06, 1.744955e-06, 3.090053e-06,
  6.587253e-07, 1.125467e-05, 1.483797e-05, 4.902978e-05, 0.0001250223, 
    0.0001283348, 2.77338e-05, 3.672043e-06, 2.302375e-06, 2.098782e-06, 
    5.761357e-06, 2.029296e-06, 2.11799e-06, 3.253412e-06, 2.920803e-06,
  9.37107e-07, 1.912092e-06, 4.949651e-06, 1.255686e-05, 0.0001015194, 
    0.0001558507, 8.439616e-05, 4.383929e-06, 3.863826e-06, 2.859053e-06, 
    1.864213e-06, 4.669436e-06, 5.926095e-06, 2.833095e-06, 1.341465e-06,
  1.219691e-06, 6.473096e-07, 7.813104e-07, 3.598291e-06, 4.246258e-05, 
    0.0001639377, 0.0001240859, 5.409143e-05, 1.305388e-05, 4.919177e-06, 
    2.462655e-06, 3.495879e-06, 4.910356e-06, 3.308768e-06, 2.832701e-06,
  7.947369e-06, 4.405259e-06, 6.423565e-06, 4.526877e-06, 4.411527e-06, 
    2.724794e-06, 1.065876e-06, 3.223993e-06, 2.342774e-05, 4.507113e-06, 
    3.442319e-06, 1.179401e-07, 3.88072e-09, 3.250308e-09, 1.675692e-09,
  3.273921e-06, 3.509487e-06, 3.882529e-06, 5.166414e-06, 6.345642e-06, 
    4.100568e-06, 1.227776e-06, 8.535409e-06, 1.410916e-05, 7.139808e-06, 
    3.031824e-06, 1.481075e-07, 4.434132e-08, 1.354031e-06, 1.009753e-06,
  5.702151e-06, 6.142648e-06, 3.977022e-06, 4.934268e-06, 4.074514e-06, 
    8.007838e-06, 1.055482e-06, 2.418185e-05, 1.48488e-05, 9.110924e-06, 
    1.388936e-06, 2.157836e-07, 1.468243e-06, 1.265424e-05, 1.243068e-07,
  8.191632e-06, 1.156613e-05, 8.413035e-06, 8.623075e-06, 3.730313e-06, 
    2.272983e-06, 1.806548e-05, 3.841209e-05, 1.35112e-05, 6.599854e-06, 
    5.589148e-06, 1.527636e-06, 8.488384e-06, 1.18255e-05, 7.660522e-08,
  8.580339e-06, 1.780142e-05, 1.262389e-05, 6.893963e-06, 5.309301e-06, 
    4.612375e-06, 3.976746e-05, 5.190476e-05, 1.565012e-05, 7.515059e-06, 
    9.652387e-06, 4.139248e-06, 6.012268e-06, 1.150448e-05, 1.296629e-05,
  6.738239e-06, 1.622464e-05, 2.083663e-05, 7.129526e-06, 6.44651e-06, 
    9.293573e-06, 6.714836e-05, 4.862268e-05, 1.595576e-06, 9.814918e-06, 
    8.139425e-06, 6.003373e-06, 8.483759e-06, 8.463433e-06, 8.802011e-06,
  5.042069e-06, 1.066963e-05, 2.637637e-05, 1.406313e-05, 8.117722e-06, 
    9.590418e-06, 6.864582e-05, 9.69582e-05, 9.301815e-06, 1.514316e-05, 
    9.206085e-06, 6.85917e-06, 1.073191e-05, 9.867138e-06, 9.94261e-06,
  3.04571e-06, 1.121406e-05, 2.553615e-05, 2.792297e-05, 7.652616e-06, 
    1.238162e-05, 6.588375e-05, 6.108329e-05, 6.444955e-06, 1.375494e-05, 
    6.99149e-06, 5.333548e-06, 1.051123e-05, 8.087361e-06, 9.100104e-06,
  1.479104e-06, 1.039318e-05, 2.265863e-05, 4.15268e-05, 2.005401e-05, 
    2.494932e-05, 5.914433e-05, 6.015715e-05, 9.455612e-06, 1.213074e-05, 
    8.025627e-06, 8.192392e-06, 9.001926e-06, 9.710556e-06, 7.572178e-06,
  1.482705e-06, 4.9099e-06, 1.606293e-05, 5.049585e-05, 5.247984e-05, 
    5.327123e-05, 6.071269e-05, 5.376215e-05, 1.056967e-05, 8.913834e-06, 
    4.666862e-06, 8.125743e-06, 7.035312e-06, 6.050684e-06, 5.780911e-06,
  5.132506e-07, 2.047324e-07, 1.900865e-06, 2.621426e-06, 3.496478e-06, 
    3.415145e-06, 4.100834e-06, 3.600638e-06, 2.428525e-07, 3.620529e-07, 
    7.880131e-06, 5.551718e-06, 1.207358e-05, 3.623887e-06, 5.536934e-07,
  4.49316e-09, 1.751149e-07, 5.905045e-07, 2.96311e-06, 5.637949e-06, 
    1.735262e-06, 1.361547e-06, 9.281378e-07, 1.000309e-07, 1.029857e-06, 
    2.520606e-06, 6.83809e-06, 2.238723e-06, 6.874802e-06, 1.23216e-06,
  1.960552e-07, 1.569406e-07, 1.302025e-06, 3.735731e-06, 7.963295e-06, 
    9.733858e-06, 3.60275e-07, 1.208467e-06, 8.375141e-08, 3.814941e-06, 
    5.489115e-06, 4.626103e-06, 2.219782e-06, 2.200762e-06, 2.429799e-07,
  2.277577e-08, 5.328938e-07, 3.628842e-06, 4.668108e-06, 4.138758e-06, 
    9.67055e-06, 8.210268e-06, 1.210342e-07, 9.02286e-08, 7.215547e-06, 
    1.329602e-05, 1.093197e-05, 4.026867e-06, 2.132093e-06, 3.592665e-08,
  7.808097e-08, 5.985646e-07, 3.434517e-06, 5.121937e-06, 4.815425e-06, 
    5.313701e-06, 5.969575e-06, 1.054464e-05, 2.344109e-06, 3.51703e-06, 
    1.738971e-05, 1.634729e-05, 4.541886e-06, 3.73595e-06, 2.589311e-06,
  7.371389e-07, 4.352218e-07, 2.3752e-06, 2.502064e-06, 2.820359e-06, 
    3.636486e-06, 4.460229e-06, 3.313147e-06, 6.417713e-06, 3.757165e-06, 
    1.130701e-05, 1.881647e-05, 7.204673e-06, 1.466913e-06, 2.238158e-06,
  2.289828e-06, 2.359888e-06, 4.195808e-06, 2.123959e-06, 1.586173e-06, 
    1.748687e-06, 4.458313e-06, 4.563777e-06, 4.595629e-06, 3.733014e-06, 
    7.176203e-06, 1.560568e-05, 1.101439e-05, 1.963749e-06, 2.863261e-06,
  4.106101e-06, 5.12097e-06, 9.528677e-06, 9.730598e-06, 4.541092e-06, 
    2.440082e-06, 3.305631e-06, 2.176491e-06, 3.182518e-06, 5.04321e-06, 
    5.937639e-06, 1.168603e-05, 1.69531e-05, 3.869014e-06, 2.747339e-06,
  8.759085e-06, 9.409358e-06, 1.5124e-05, 1.516767e-05, 5.098119e-06, 
    2.755855e-06, 4.689511e-06, 1.406426e-06, 2.450965e-06, 4.265859e-06, 
    5.006654e-06, 9.862553e-06, 2.06763e-05, 8.494744e-06, 7.596824e-06,
  8.291918e-06, 8.729433e-06, 1.546256e-05, 2.330941e-05, 1.512681e-05, 
    5.9212e-06, 5.012377e-06, 2.990155e-06, 4.304609e-06, 4.302113e-06, 
    4.535686e-06, 6.726454e-06, 1.755487e-05, 9.045098e-06, 7.838393e-06,
  4.31121e-09, 3.516037e-08, 4.952718e-07, 1.883714e-06, 3.765735e-06, 
    2.766744e-06, 2.369893e-06, 4.637514e-06, 3.713476e-06, 6.332411e-06, 
    3.439291e-06, 1.870285e-06, 4.48181e-07, 6.652729e-08, 7.361859e-08,
  2.164003e-08, 3.085102e-08, 1.879883e-08, 4.179065e-07, 4.000275e-06, 
    6.107191e-07, 6.466792e-07, 1.257575e-06, 3.881923e-06, 1.065642e-05, 
    4.60424e-06, 2.014811e-06, 1.639836e-06, 2.676942e-06, 5.311339e-06,
  1.783442e-07, 2.274084e-08, 9.389782e-08, 3.157288e-07, 9.11025e-07, 
    7.063614e-06, 1.985206e-07, 1.690855e-06, 1.311166e-06, 1.931627e-05, 
    5.716719e-06, 9.51559e-07, 5.067443e-06, 7.922281e-06, 4.563819e-07,
  6.320097e-07, 2.423662e-07, 1.117632e-06, 2.815509e-07, 1.191767e-06, 
    1.870248e-06, 5.198242e-06, 5.437837e-08, 1.480592e-07, 8.71796e-06, 
    9.503712e-06, 2.838931e-06, 7.554742e-06, 1.087679e-05, 1.281537e-07,
  9.060742e-09, 1.972817e-08, 7.068929e-07, 1.265563e-06, 1.169998e-06, 
    1.115628e-06, 3.464067e-06, 2.479568e-06, 3.795855e-06, 1.145582e-06, 
    8.100205e-06, 1.176885e-05, 6.114071e-06, 8.011136e-06, 3.813829e-06,
  3.51737e-07, 5.067248e-07, 1.292138e-06, 8.703175e-07, 1.083539e-07, 
    9.585376e-07, 1.060566e-06, 2.353572e-06, 5.935485e-06, 1.257698e-06, 
    5.953702e-07, 1.204511e-05, 5.141228e-06, 8.695578e-06, 4.652111e-06,
  3.017029e-06, 3.582433e-06, 3.940171e-06, 4.815094e-06, 4.717233e-06, 
    1.944431e-06, 1.236397e-06, 1.613786e-06, 2.1069e-06, 1.911864e-06, 
    1.341584e-06, 2.364174e-06, 9.312658e-06, 8.525692e-06, 3.59332e-06,
  4.987256e-06, 3.565184e-06, 4.530831e-06, 6.387419e-06, 4.498636e-06, 
    4.616617e-06, 3.40939e-06, 3.128582e-06, 1.613143e-06, 1.806191e-06, 
    1.746757e-06, 1.040848e-06, 6.796685e-06, 7.251197e-06, 4.336337e-06,
  9.114415e-06, 6.036812e-06, 5.219517e-06, 3.903279e-06, 5.001434e-06, 
    2.886504e-06, 3.825489e-06, 3.620652e-06, 2.336184e-06, 1.894108e-06, 
    2.062875e-06, 1.091066e-06, 4.376878e-06, 8.398772e-06, 8.507018e-06,
  7.697294e-06, 7.683064e-06, 5.335255e-06, 4.780029e-06, 3.518667e-06, 
    3.438246e-06, 4.61609e-06, 4.266741e-06, 4.424621e-06, 3.04527e-06, 
    2.498964e-06, 2.668529e-06, 3.7478e-06, 3.356839e-06, 1.112358e-05 ;

 scalar_axis = 0 ;


 time = 0.5, 1.5, 2.5, 3.5, 4.5, 5.5, 6.5, 7.5, 8.5, 9.5, 10.5, 11.5, 12.5, 
    13.5, 14.5, 15.5, 16.5, 17.5, 18.5, 19.5, 20.5, 21.5, 22.5, 23.5, 24.5, 
    25.5, 26.5, 27.5, 28.5, 29.5, 30.5, 31.5, 32.5, 33.5, 34.5, 35.5, 36.5, 
    37.5, 38.5, 39.5, 40.5, 41.5, 42.5, 43.5, 44.5, 45.5, 46.5, 47.5, 48.5, 
    49.5, 50.5, 51.5, 52.5, 53.5, 54.5, 55.5, 56.5, 57.5, 58.5, 59.5, 60.5, 
    61.5, 62.5, 63.5, 64.5, 65.5, 66.5, 67.5, 68.5, 69.5, 70.5, 71.5, 72.5, 
    73.5, 74.5, 75.5, 76.5, 77.5, 78.5, 79.5, 80.5, 81.5, 82.5, 83.5, 84.5, 
    85.5, 86.5, 87.5, 88.5, 89.5, 90.5, 91.5, 92.5, 93.5, 94.5, 95.5, 96.5, 
    97.5, 98.5, 99.5, 100.5, 101.5, 102.5, 103.5, 104.5, 105.5, 106.5, 107.5, 
    108.5, 109.5, 110.5, 111.5, 112.5, 113.5, 114.5, 115.5, 116.5, 117.5, 
    118.5, 119.5, 120.5, 121.5, 122.5, 123.5, 124.5, 125.5, 126.5, 127.5, 
    128.5, 129.5, 130.5, 131.5, 132.5, 133.5, 134.5, 135.5, 136.5, 137.5, 
    138.5, 139.5, 140.5, 141.5, 142.5, 143.5, 144.5, 145.5, 146.5, 147.5, 
    148.5, 149.5, 150.5, 151.5, 152.5, 153.5, 154.5, 155.5, 156.5, 157.5, 
    158.5, 159.5, 160.5, 161.5, 162.5, 163.5, 164.5, 165.5, 166.5, 167.5, 
    168.5, 169.5, 170.5, 171.5, 172.5, 173.5, 174.5, 175.5, 176.5, 177.5, 
    178.5, 179.5, 180.5, 181.5 ;

 time_bnds =
  0, 1,
  1, 2,
  2, 3,
  3, 4,
  4, 5,
  5, 6,
  6, 7,
  7, 8,
  8, 9,
  9, 10,
  10, 11,
  11, 12,
  12, 13,
  13, 14,
  14, 15,
  15, 16,
  16, 17,
  17, 18,
  18, 19,
  19, 20,
  20, 21,
  21, 22,
  22, 23,
  23, 24,
  24, 25,
  25, 26,
  26, 27,
  27, 28,
  28, 29,
  29, 30,
  30, 31,
  31, 32,
  32, 33,
  33, 34,
  34, 35,
  35, 36,
  36, 37,
  37, 38,
  38, 39,
  39, 40,
  40, 41,
  41, 42,
  42, 43,
  43, 44,
  44, 45,
  45, 46,
  46, 47,
  47, 48,
  48, 49,
  49, 50,
  50, 51,
  51, 52,
  52, 53,
  53, 54,
  54, 55,
  55, 56,
  56, 57,
  57, 58,
  58, 59,
  59, 60,
  60, 61,
  61, 62,
  62, 63,
  63, 64,
  64, 65,
  65, 66,
  66, 67,
  67, 68,
  68, 69,
  69, 70,
  70, 71,
  71, 72,
  72, 73,
  73, 74,
  74, 75,
  75, 76,
  76, 77,
  77, 78,
  78, 79,
  79, 80,
  80, 81,
  81, 82,
  82, 83,
  83, 84,
  84, 85,
  85, 86,
  86, 87,
  87, 88,
  88, 89,
  89, 90,
  90, 91,
  91, 92,
  92, 93,
  93, 94,
  94, 95,
  95, 96,
  96, 97,
  97, 98,
  98, 99,
  99, 100,
  100, 101,
  101, 102,
  102, 103,
  103, 104,
  104, 105,
  105, 106,
  106, 107,
  107, 108,
  108, 109,
  109, 110,
  110, 111,
  111, 112,
  112, 113,
  113, 114,
  114, 115,
  115, 116,
  116, 117,
  117, 118,
  118, 119,
  119, 120,
  120, 121,
  121, 122,
  122, 123,
  123, 124,
  124, 125,
  125, 126,
  126, 127,
  127, 128,
  128, 129,
  129, 130,
  130, 131,
  131, 132,
  132, 133,
  133, 134,
  134, 135,
  135, 136,
  136, 137,
  137, 138,
  138, 139,
  139, 140,
  140, 141,
  141, 142,
  142, 143,
  143, 144,
  144, 145,
  145, 146,
  146, 147,
  147, 148,
  148, 149,
  149, 150,
  150, 151,
  151, 152,
  152, 153,
  153, 154,
  154, 155,
  155, 156,
  156, 157,
  157, 158,
  158, 159,
  159, 160,
  160, 161,
  161, 162,
  162, 163,
  163, 164,
  164, 165,
  165, 166,
  166, 167,
  167, 168,
  168, 169,
  169, 170,
  170, 171,
  171, 172,
  172, 173,
  173, 174,
  174, 175,
  175, 176,
  176, 177,
  177, 178,
  178, 179,
  179, 180,
  180, 181,
  181, 182 ;

}
