netcdf atmos.1980-1981.alb_sfc.05 {
dimensions:
	time = UNLIMITED ; // (1 currently)
	lat = 18 ;
	lon = 29 ;
	bnds = 2 ;
variables:
	float alb_sfc(time, lat, lon) ;
		alb_sfc:long_name = "Surface Albedo for  Flux" ;
		alb_sfc:units = "percent" ;
		alb_sfc:_FillValue = 1.e+20f ;
		alb_sfc:missing_value = 1.e+20f ;
		alb_sfc:cell_measures = "area: area" ;
		alb_sfc:interp_method = "conserve_order1" ;
		alb_sfc:cell_methods = "time: mean within months time: mean over years" ;
		alb_sfc:time_avg_info = "average_T1,average_T2,average_DT" ;
	double average_DT(time) ;
		average_DT:long_name = "Length of average period" ;
		average_DT:units = "days" ;
	double average_T1(time) ;
		average_T1:long_name = "Start time for average period" ;
		average_T1:units = "days since 1979-01-01 00:00:00" ;
	double average_T2(time) ;
		average_T2:long_name = "End time for average period" ;
		average_T2:units = "days since 1979-01-01 00:00:00" ;
	double climatology_bounds(time, bnds) ;
	double lat(lat) ;
		lat:standard_name = "latitude" ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_N" ;
		lat:axis = "Y" ;
		lat:bounds = "lat_bnds" ;
	double lat_bnds(lat, bnds) ;
	double lon(lon) ;
		lon:standard_name = "longitude" ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_E" ;
		lon:axis = "X" ;
		lon:bounds = "lon_bnds" ;
	double lon_bnds(lon, bnds) ;
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:climatology = "climatology_bounds" ;
		time:units = "days since 1979-01-01 00:00:00" ;
		time:calendar = "standard" ;
		time:axis = "T" ;

// global attributes:
		:CDI = "Climate Data Interface version 2.4.4 (https://mpimet.mpg.de/cdi)" ;
		:Conventions = "CF-1.6" ;
		:title = "c96L65_am5f9d8r0_amip" ;
		:associated_files = "area: 19800101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:code_release_version = "2024.05" ;
		:git_hash = "5d306c05d9fe755cab04eedc8fd3de0d3c8355a0" ;
		:creationtime = "Mon Aug 25 14:09:46 2025" ;
		:hostname = "pp050" ;
		:history = "Mon Aug 25 13:32:18 2025: ncks -d lat,,,10 -d lon,,,10 atmos.1980-1981.alb_sfc.05.nc reduced/atmos.1980-1981.alb_sfc.05.nc\n",
			"Mon Aug 25 14:40:05 2025: cdo -O -s -select,month=5 merged_output.nc monthly_nc_files/all_years.5.nc\n",
			"Mon Aug 25 14:40:01 2025: cdo -O -s -mergetime /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/shards/ts/regrid-xy/180_288.conserve_order2/atmos_month/P1M/P1Y/atmos_month.198001-198012.alb_sfc.nc /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/shards/ts/regrid-xy/180_288.conserve_order2/atmos_month/P1M/P1Y/atmos_month.198101-198112.alb_sfc.nc merged_output.nc\n",
			"Mon Aug 25 14:12:17 2025: cdo --history splitname 19800101.atmos_month.nc /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/split/regrid-xy/180_288.conserve_order2/19800101.atmos_month.\n",
			"fregrid --debug --standard_dimension --input_mosaic C96_mosaic.nc --input_dir /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/history/native --input_file 19800101.atmos_month --associated_file_dir /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/history/native --interp_method conserve_order2 --remap_file fregrid_remap_file_288_by_180.nc --nlon 288 --nlat 180 --scalar_field (**please see the field list in this file**) --output_file 19800101.atmos_month.nc" ;
		:CDO = "Climate Data Operators version 2.4.4 (https://mpimet.mpg.de/cdo)" ;
		:comment = "FMS time averaging, version 3.0, precision=double" ;
		:NCO = "netCDF Operators version 5.2.4 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 alb_sfc =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  9.315227, 10.34629, 9.541336, 8.956, 9.375626, 9.345503, 10.41593, 
    9.410661, 9.590737, 9.664564, 9.523396, 9.391825, 9.373642, 8.994425, 
    6.691735, 5.967158, 5.755425, 4.86621, 3.144291, 5.907794, 8.391279, 
    7.376364, 9.095936, 9.128046, 10.93114, 11.12055, 10.37096, 10.67018, 
    10.98792,
  3.227689, 3.376851, 3.51312, 3.495361, 3.086202, 3.171341, 2.922724, 
    3.284616, 3.191985, 3.166385, 3.08326, 2.975619, 2.769753, 2.860591, 
    3.074463, 2.901403, 3.092146, 3.27263, 3.289683, 3.523782, 3.329674, 
    3.330898, 3.159152, 2.784958, 2.616785, 6.229997, 8.645849, 2.842087, 
    3.00063,
  3.467694, 3.263082, 3.544885, 3.356402, 3.427048, 3.357849, 3.338865, 
    3.482047, 3.538132, 3.706975, 3.665656, 3.41745, 3.497999, 3.400967, 
    3.460522, 3.623785, 3.674454, 3.731247, 3.993306, 3.781584, 3.817134, 
    3.8564, 3.312707, 6.187984, 3.822006, 3.295657, 3.185718, 3.42124, 
    3.366722,
  3.399229, 3.902489, 3.921805, 3.69517, 3.703316, 3.801198, 3.639075, 
    3.711672, 3.813079, 3.896279, 4.025496, 3.992018, 4.03173, 3.867468, 
    7.388952, 3.880878, 3.695259, 3.759204, 3.625407, 3.607922, 3.529266, 
    3.68997, 3.738098, 7.541125, 4.102207, 3.821036, 4.034548, 3.758322, 
    3.60208,
  3.822296, 4.145777, 11.2161, 4.008784, 3.98181, 3.994334, 3.972641, 
    4.023785, 3.854388, 4.05711, 9.098351, 13.14781, 9.457155, 4.083877, 
    3.891454, 3.661244, 3.744233, 3.71077, 3.456757, 3.618692, 3.734815, 
    3.824527, 3.870749, 4.239537, 8.318481, 3.930769, 3.916754, 3.956764, 
    3.867814,
  3.728884, 9.36224, 10.85146, 3.900688, 3.718375, 3.777515, 3.74753, 
    3.950277, 3.563082, 4.068318, 11.38541, 11.64131, 3.961482, 3.655666, 
    3.707916, 3.682545, 3.791664, 3.564642, 3.876626, 3.747868, 4.022102, 
    3.895439, 3.573172, 3.847096, 8.700519, 8.818244, 3.660357, 4.138689, 
    3.586023,
  3.443919, 6.277357, 9.026695, 8.858206, 3.38299, 3.373006, 3.365948, 
    3.475805, 3.283594, 3.418563, 4.439122, 3.541595, 4.194944, 3.275928, 
    3.577508, 3.516071, 3.795824, 3.755558, 3.902683, 3.752987, 3.931529, 
    3.614608, 3.221654, 8.602573, 8.545502, 8.715535, 3.827954, 3.808989, 
    3.438847,
  3.24108, 8.356108, 8.129475, 9.875414, 3.517595, 3.433336, 3.418583, 
    3.375093, 8.605091, 8.270144, 3.396075, 3.435077, 3.628129, 3.57872, 
    3.482556, 3.565988, 3.585059, 3.696088, 3.645716, 3.75978, 3.656106, 
    3.657391, 3.179319, 8.223961, 8.435246, 3.385286, 3.464901, 3.372029, 
    3.293659,
  9.891521, 10.34822, 10.62297, 9.8488, 15.33679, 3.316631, 5.124622, 
    3.235157, 3.620952, 3.269718, 4.502257, 3.314658, 3.358404, 3.290248, 
    3.318104, 3.328341, 3.280668, 3.563137, 3.346688, 3.514529, 3.31153, 
    3.370025, 8.996595, 7.43478, 3.573122, 3.345837, 3.397923, 3.142288, 
    8.965476,
  18.81184, 21.49005, 23.61653, 3.467838, 23.86943, 3.587384, 11.24572, 
    3.309018, 9.448616, 3.366932, 3.722297, 3.599894, 3.5844, 3.68028, 
    3.749297, 3.787791, 3.681931, 3.84277, 3.45777, 3.682419, 3.944757, 
    6.776785, 3.683537, 4.175476, 3.568425, 3.621579, 3.852234, 3.624187, 
    24.57278,
  25.31693, 21.36546, 22.21407, 20.43048, 13.37598, 15.21047, 13.18178, 
    17.65078, 9.58258, 10.82275, 3.642455, 3.580141, 3.553987, 3.658432, 
    3.783865, 3.667621, 3.799699, 3.757928, 3.669127, 3.943927, 11.31887, 
    12.33128, 9.874399, 3.769473, 3.704233, 3.730701, 3.733134, 3.748908, 
    11.79719,
  8.354622, 4.059175, 6.423914, 10.93807, 2.25141, 15.88468, 10.39898, 
    16.63562, 14.34889, 11.68631, 8.162962, 4.050352, 3.914348, 3.793821, 
    3.73597, 3.7701, 3.830188, 3.737904, 3.796819, 13.06235, 11.99576, 
    14.76489, 13.81985, 4.797532, 3.870162, 3.955023, 3.936255, 4.245406, 
    5.293092,
  6.530665, 13.59773, 15.2687, 15.96566, 14.77654, 12.95619, 9.126854, 
    23.7811, 9.980349, 8.342518, 8.152871, 8.61923, 4.229256, 4.303335, 
    4.195891, 4.160845, 4.11981, 4.276142, 4.309749, 11.01408, 11.55526, 
    10.97829, 7.785349, 12.36461, 5.717352, 4.066529, 4.320925, 4.325253, 
    4.387384,
  5.241005, 8.822186, 11.77337, 8.656593, 9.910458, 9.702132, 17.775, 
    20.59941, 12.30763, 11.89044, 9.891288, 43.69605, 48.05891, 31.75549, 
    5.757899, 5.540265, 19.71458, 20.75815, 34.78181, 8.597003, 8.571713, 
    35.6644, 48.38116, 40.42075, 4.960068, 10.2443, 4.543864, 4.779098, 
    5.016929,
  6.337687, 7.263758, 27.98028, 7.009218, 40.57874, 72.92844, 65.12985, 
    64.16106, 64.35599, 64.1152, 38.14975, 31.93423, 63.0641, 71.83592, 
    71.42769, 66.80812, 59.8702, 53.21343, 61.02293, 60.48425, 59.92126, 
    64.99384, 58.21626, 64.01723, 63.75109, 69.48351, 70.51353, 62.67989, 
    6.240237,
  74.39044, 74.32516, 77.64673, 83.58186, 78.16887, 82.96732, 84.51709, 
    81.78259, 81.45703, 81.22802, 81.60091, 80.98, 80.228, 78.40942, 
    78.05727, 77.77582, 76.10445, 75.11678, 75.61371, 75.78523, 75.4718, 
    72.25565, 71.98791, 75.28175, 73.8129, 76.3017, 76.48036, 72.58675, 
    76.27917 ;

 average_DT = 730 ;

 average_T1 = 136.5 ;

 average_T2 = 866.5 ;

 climatology_bounds =
  136.5, 866.5 ;

 lat = -89.5, -79.5, -69.5, -59.5, -49.5, -39.5, -29.5, -19.5, -9.5, 0.5, 
    10.5, 20.5, 30.5, 40.5, 50.5, 60.5, 70.5, 80.5 ;

 lat_bnds =
  -90, -89,
  -80, -79,
  -70, -69,
  -60, -59,
  -50, -49,
  -40, -39,
  -30, -29,
  -20, -19,
  -10, -9,
  0, 1,
  10, 11,
  20, 21,
  30, 31,
  40, 41,
  50, 51,
  60, 61,
  70, 71,
  80, 81 ;

 lon = 0.625, 13.125, 25.625, 38.125, 50.625, 63.125, 75.625, 88.125, 
    100.625, 113.125, 125.625, 138.125, 150.625, 163.125, 175.625, 188.125, 
    200.625, 213.125, 225.625, 238.125, 250.625, 263.125, 275.625, 288.125, 
    300.625, 313.125, 325.625, 338.125, 350.625 ;

 lon_bnds =
  0, 1.25,
  12.5, 13.75,
  25, 26.25,
  37.5, 38.75,
  50, 51.25,
  62.5, 63.75,
  75, 76.25,
  87.5, 88.75,
  100, 101.25,
  112.5, 113.75,
  125, 126.25,
  137.5, 138.75,
  150, 151.25,
  162.5, 163.75,
  175, 176.25,
  187.5, 188.75,
  200, 201.25,
  212.5, 213.75,
  225, 226.25,
  237.5, 238.75,
  250, 251.25,
  262.5, 263.75,
  275, 276.25,
  287.5, 288.75,
  300, 301.25,
  312.5, 313.75,
  325, 326.25,
  337.5, 338.75,
  350, 351.25 ;

 time = 0 ;
}
