netcdf atmos_4xdaily.0001010100-0005123118.slp.tile1 {
dimensions:
	grid_xt = 1 ;
	grid_yt = 1 ;
	time = UNLIMITED ; // (7300 currently)
variables:
	double grid_xt(grid_xt) ;
		grid_xt:standard_name = "longitude" ;
		grid_xt:long_name = "T-cell longitude" ;
		grid_xt:units = "degrees_E" ;
		grid_xt:axis = "X" ;
	double grid_yt(grid_yt) ;
		grid_yt:standard_name = "latitude" ;
		grid_yt:long_name = "T-cell latitude" ;
		grid_yt:units = "degrees_N" ;
		grid_yt:axis = "Y" ;
	float slp(time, grid_yt, grid_xt) ;
		slp:long_name = "sea level pressure" ;
		slp:units = "pa" ;
		slp:_FillValue = 1.e+20f ;
		slp:missing_value = 1.e+20f ;
		slp:cell_methods = "time: point" ;
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:units = "days since 0001-01-01 00:00:00" ;
		time:calendar = "365_day" ;
		time:axis = "T" ;

// global attributes:
		:CDI = "Climate Data Interface version 2.4.4 (https://mpimet.mpg.de/cdi)" ;
		:Conventions = "CF-1.6" ;
		:title = "proto4_c48l33o1degSPEAR" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:history = "Wed Jan 28 16:56:37 2026: ncks -d grid_xt,0,0 -d grid_yt,0,0 /home/Dana.Singh/PT6H/P10Y/atmos_4xdaily.0001010100-0005123118.slp.tile1.nc fre/tests/test_files/ascii_files/atmos_4xdaily.0001010100-0005123118.slp.tile1.nc\nTue Jan 27 16:11:07 2026: cdo --history -O mergetime atmos_4xdaily.0001010100-0001123118.slp.tile1.nc atmos_4xdaily.0002010100-0002123118.slp.tile1.nc atmos_4xdaily.0003010100-0003123118.slp.tile1.nc atmos_4xdaily.0004010100-0004123018.slp.tile1.nc atmos_4xdaily.0005010100-0005123118.slp.tile1.nc /home/Niki.Zadeh/cylc-run/proto4_c48l33o1degSPEAR__gfdl.ncrc5-intel23__prod-openmp/share/shards/ts/native/atmos_4xdaily/PT6H/P10Y/atmos_4xdaily.0001010100-0005123118.slp.tile1.nc" ;
		:CDO = "Climate Data Operators version 2.4.4 (https://mpimet.mpg.de/cdo)" ;
		:NCO = "netCDF Operators version 5.2.4 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 grid_xt = 1 ;

 grid_yt = 1 ;

 slp =
  101330.1,
  101555.5,
  101604.3,
  101604.7,
  101638.4,
  101750.6,
  101664.9,
  101729.3,
  101610.5,
  101520,
  101348.8,
  101223.5,
  100981.1,
  100716.4,
  100433.6,
  100349.6,
  100280.6,
  100389.5,
  100900.2,
  101138.7,
  101416,
  101705.5,
  101849,
  101927.3,
  101863,
  101928.8,
  101838.1,
  101584,
  101358.1,
  101336.3,
  101171.3,
  100897.7,
  100784.8,
  100631.6,
  100262.2,
  100027.3,
  99788.7,
  99792.68,
  99815.77,
  99890.49,
  99994.74,
  100110.3,
  100071.9,
  100037.7,
  100097.2,
  100243.9,
  100174.4,
  100082.9,
  100081.9,
  100272.6,
  100220.6,
  100270.4,
  100316.5,
  100524.2,
  100557.8,
  100673.4,
  100799.7,
  101017.5,
  101026.6,
  101222.4,
  101452.2,
  101718,
  101827.6,
  101792.5,
  101805.5,
  101745.8,
  101604.5,
  101501.9,
  101433.5,
  101505.1,
  101303.8,
  101167.9,
  101127.6,
  101116.9,
  100991.5,
  100977.8,
  101007.8,
  101152.6,
  101139.4,
  100965.6,
  100963.6,
  101040.2,
  100880.2,
  100746.7,
  100661.6,
  100694.6,
  100514.5,
  100388.5,
  100250.7,
  100293.3,
  100314.5,
  100258.7,
  100354.4,
  100640.3,
  101000,
  101371.6,
  101542.9,
  101847.1,
  101888.5,
  101882.2,
  101926.8,
  101975.6,
  101906.2,
  101894.3,
  101860.5,
  101956.9,
  101981.7,
  101864.8,
  101796.2,
  102042.4,
  101932.2,
  101813.1,
  101750.2,
  101717.6,
  101551.6,
  101360.2,
  101315.3,
  101320.1,
  101188.1,
  101187.5,
  101268.2,
  101365.7,
  101261.7,
  101302.4,
  101361.8,
  101513.9,
  101517.4,
  101499.4,
  101475.6,
  101606.3,
  101540.1,
  101468,
  101542.6,
  101642.3,
  101476,
  101242.1,
  101332,
  101381.6,
  101197,
  101183.2,
  101182.2,
  101342.3,
  101322.1,
  101342.2,
  101449.2,
  101666.2,
  101649.7,
  101698,
  101765.9,
  101933.1,
  101807.4,
  101773.4,
  101822.8,
  101967.8,
  101831,
  101671.6,
  101637.9,
  101712.5,
  101379.7,
  101300.5,
  101124.8,
  101190.2,
  101036.4,
  100932.7,
  100849.7,
  100934.9,
  100827.5,
  100821.7,
  100849.2,
  100990.9,
  100932.2,
  101025.9,
  101095,
  101251.8,
  101157.2,
  101105.2,
  101144.9,
  101254.2,
  101109.8,
  101208.3,
  101294,
  101448.9,
  101499.1,
  101626.3,
  101685.9,
  101791.4,
  101627.1,
  101337.5,
  101310.8,
  101225.7,
  100855.8,
  100704.9,
  100716.9,
  100741.4,
  100713.5,
  100923,
  101184.2,
  101360.1,
  101429.5,
  101457.5,
  101525.5,
  101689.5,
  101529.3,
  101378.3,
  101239,
  101188.3,
  100812.2,
  100996.6,
  101104.4,
  101203.3,
  101102.6,
  101096.4,
  101023.8,
  101111.5,
  101014.9,
  100964.3,
  101036.6,
  101201.1,
  101148.1,
  101073.4,
  101155.7,
  101327.9,
  101202.5,
  101181.7,
  101211.5,
  101214,
  100915.2,
  100846.2,
  100803.3,
  100896.1,
  100696.2,
  100584.4,
  100638.8,
  100622.4,
  100750.5,
  100952.7,
  101246,
  101481,
  101444.5,
  101418.6,
  101388.7,
  101395.7,
  101240.8,
  101261.2,
  101339.3,
  101512.9,
  101324.8,
  101225.9,
  101226.7,
  101277.8,
  101043,
  101056.2,
  101155.3,
  101361.1,
  101508.6,
  101742.6,
  101719.7,
  101835.4,
  101746.1,
  101454.3,
  101092.1,
  100790.2,
  100552.6,
  100622.4,
  100750.7,
  100837.7,
  100763.5,
  100663.7,
  100450.6,
  100313.9,
  100033.1,
  99814.49,
  99826.03,
  100035.9,
  100266.1,
  100679.9,
  101007.5,
  101265.1,
  101420,
  101750.5,
  101909.3,
  102102.8,
  102254,
  102279.3,
  102411.8,
  102564.8,
  102421.5,
  102255.8,
  102197.3,
  102317.2,
  102100.4,
  101926,
  101839.1,
  101896.5,
  101595.8,
  101356.2,
  101351.2,
  101341,
  101071,
  100894,
  100936.1,
  101000.4,
  100799.6,
  100790.2,
  100656.9,
  100542.5,
  100164.5,
  100108.1,
  99872.85,
  100488.4,
  100908.1,
  101130,
  101295,
  101608.3,
  101703.2,
  101766.1,
  101863.6,
  101990.4,
  101773.4,
  101672.9,
  101805.4,
  101793.7,
  101583.6,
  101547.4,
  101642.7,
  101791.5,
  101734.5,
  101857,
  101961.9,
  102118.9,
  102124.3,
  102152.9,
  102118.6,
  102242.4,
  102161.4,
  102073.7,
  102000.9,
  102060,
  101936.4,
  101827.4,
  101754.1,
  101770.8,
  101600.4,
  101495.8,
  101438,
  101456.4,
  101251.4,
  101094.5,
  101049.5,
  101078.8,
  100954.1,
  101096.6,
  101097.3,
  101308.2,
  101191.3,
  101387,
  101360.1,
  101559.2,
  101535.3,
  101782.8,
  101685.5,
  101899.5,
  101835.7,
  101791.1,
  101702.3,
  101746.8,
  101589.8,
  101513.9,
  101455.9,
  101626.2,
  101766.4,
  101848.8,
  101794.7,
  102103.6,
  102012,
  101988,
  101869.9,
  101853.6,
  101567.4,
  101451.8,
  101311.8,
  101121.6,
  100572.6,
  101031,
  101156.3,
  101456.1,
  101669.9,
  101898.6,
  102014.1,
  102124.1,
  101981.8,
  101828.2,
  101632.5,
  101515.4,
  101309.4,
  101364.1,
  101361.9,
  101491.3,
  101381.7,
  101345.5,
  101346.3,
  101412.8,
  101252,
  101363.8,
  101450.8,
  101633.9,
  101636.8,
  101817.6,
  101850.4,
  101968.9,
  101839,
  101827.4,
  101741,
  101641.7,
  101360.8,
  101328.2,
  101326.8,
  101348.9,
  101185.7,
  101005.1,
  100954.8,
  100928.4,
  100947.8,
  101160.2,
  101345.7,
  101401.7,
  101372.3,
  101473.5,
  101424.6,
  101423.3,
  101273.6,
  101208.8,
  101223.4,
  101305.3,
  101218.6,
  101248,
  101276.3,
  101381.8,
  101268.4,
  101293.9,
  101311.5,
  101416.5,
  101463.2,
  101698.8,
  101704.4,
  101645.2,
  101950.2,
  101657.5,
  101831.7,
  101914.9,
  101727.3,
  101647,
  101693.1,
  101688.2,
  101552.4,
  101675.7,
  101603.1,
  101599.3,
  101476.4,
  101589.2,
  101668.2,
  101910.5,
  102157.2,
  102377.5,
  102387.2,
  102496.8,
  102464.8,
  102355.8,
  102313.6,
  102359.2,
  102194.1,
  102325.1,
  102339.6,
  102420.1,
  102401.8,
  102452.1,
  102468.8,
  102529.7,
  102353.7,
  102322.7,
  102242,
  102255.4,
  102038.4,
  102009.7,
  101941,
  101965.4,
  101767.8,
  101740.4,
  101708.4,
  101744.2,
  101682.6,
  101744.7,
  101783.8,
  101955.6,
  101902.1,
  101809.2,
  101639.5,
  101489.9,
  101169.4,
  101065.7,
  100987.1,
  101122,
  101039.7,
  101181.6,
  101301.7,
  101380.8,
  101218.6,
  101185.9,
  101188.5,
  101308.3,
  101524.5,
  101732.3,
  101965.8,
  102173.6,
  102159,
  102170,
  102220,
  102197.7,
  101667.1,
  101373.5,
  101446.8,
  101535.5,
  101649.6,
  101791.3,
  101763.7,
  101831.3,
  101628.4,
  101499.3,
  101204.9,
  100715.2,
  100595.1,
  100297.1,
  100897.5,
  101336.5,
  101610.3,
  101885.4,
  101963.1,
  102007.7,
  101907.3,
  102027.9,
  101954.5,
  101958.9,
  101856.8,
  101695,
  101648.6,
  101730.1,
  101616.4,
  101576.2,
  101423.4,
  101246.5,
  101015.9,
  101083.1,
  101123.8,
  101186,
  101066.4,
  101060.6,
  101013.9,
  101100.9,
  101090.3,
  101062,
  100885.8,
  100723.5,
  100396.9,
  100731.1,
  101087.7,
  101482,
  101730.2,
  102093.3,
  102276.7,
  102476,
  102550.1,
  102675.9,
  102680.2,
  102640.2,
  102481.8,
  102489.2,
  102402,
  102426,
  102253.2,
  102199.9,
  102145.1,
  102195.2,
  102045.1,
  101985.5,
  101874,
  101889.7,
  101720.5,
  101693,
  101661.1,
  101723.7,
  101570.8,
  101615.8,
  101609.2,
  101651.5,
  101532,
  101468.2,
  101342.1,
  101288.9,
  101114.4,
  101353.5,
  101620.3,
  101772.2,
  101583.8,
  101554.4,
  101019.3,
  100695.9,
  101079.9,
  101328.8,
  101385.6,
  101492.3,
  101308.3,
  101453.2,
  101504.7,
  101718.6,
  101905.1,
  101960.1,
  101889.4,
  101836.7,
  101668.4,
  101669.3,
  101439.9,
  101253.7,
  100911.6,
  100978.4,
  101107.6,
  101291.4,
  101427.2,
  101553.4,
  101431.9,
  101312.4,
  100844.9,
  100543.6,
  100377.5,
  100708.1,
  101244.7,
  101806.1,
  102171,
  102482,
  102500.4,
  102481.7,
  102376.2,
  102325.1,
  102332.8,
  102480.5,
  102545.3,
  102693.1,
  102711.7,
  102768.8,
  102775.2,
  102785.6,
  102634.5,
  102609.7,
  102565.9,
  102581.5,
  102488.3,
  102564.4,
  102469.3,
  102525.3,
  102488,
  102515.2,
  102544.8,
  102633.8,
  102567.2,
  102623.6,
  102574.3,
  102687.1,
  102710.8,
  102834.7,
  102940.5,
  103109.9,
  103234.6,
  103362.3,
  103353.2,
  103455,
  103361.6,
  103315.6,
  103136.9,
  103024.7,
  102669.2,
  102517.8,
  102276.6,
  102268.2,
  102206.8,
  102295.7,
  102350.8,
  102393.6,
  102228.9,
  102143.8,
  101955.4,
  101754.6,
  101353.6,
  101155,
  101107.6,
  101161.3,
  101258.4,
  101752.4,
  102304.7,
  102830,
  102925,
  103066.6,
  103097.9,
  103070.5,
  102683.4,
  102471,
  102309.4,
  102262.8,
  102086.8,
  102042.3,
  102068.1,
  102181.3,
  102150.5,
  102322.1,
  102456.7,
  102596.3,
  102518.6,
  102509,
  102364.2,
  102238.6,
  101958.2,
  102043.7,
  102140.9,
  102346.1,
  102285.4,
  102518.6,
  102464.8,
  102577.1,
  102382.6,
  102323.9,
  102194.1,
  102096.7,
  101905.3,
  101782.9,
  101407.2,
  101240,
  101368,
  101556.2,
  101471.9,
  101441.8,
  101375.5,
  101506.3,
  101576,
  101816.2,
  101866.5,
  101951.4,
  101815.5,
  101774.7,
  101513,
  101500.8,
  101544.5,
  101682.6,
  101636.6,
  101886.7,
  102111.4,
  102277.2,
  102268.5,
  102326.4,
  102214.9,
  102182.6,
  102014.6,
  101981.9,
  101990.2,
  101929.7,
  101765.2,
  101740.1,
  101614.3,
  101727.8,
  102004.2,
  102253.2,
  102218,
  102199.3,
  101940.6,
  101812.8,
  101794.9,
  102075.8,
  102190.5,
  102382.3,
  102425.2,
  102516.7,
  102289.4,
  102035,
  101772.7,
  101531.9,
  101279.8,
  101491.2,
  101991.7,
  102283.8,
  102643,
  103021.2,
  103180.2,
  103355,
  103390.6,
  103446.3,
  103250.2,
  103191.7,
  103005.8,
  102963.1,
  102869.1,
  102841.8,
  102641.9,
  102589.5,
  102440.8,
  102347.1,
  101963.1,
  101853.7,
  101759.7,
  101735,
  101567.4,
  101592.8,
  101638.2,
  101710.3,
  101817,
  102097.4,
  102238.5,
  102506.4,
  102613.5,
  102741.1,
  102712.9,
  102724.8,
  102554.1,
  102496.2,
  102429.4,
  102490.9,
  102378.5,
  102379.9,
  102332.6,
  102654.6,
  102577.7,
  102674.5,
  102662.6,
  102774.9,
  102690.6,
  102746.3,
  102731,
  102778.7,
  102599.8,
  102595.5,
  102495,
  102413.9,
  102253.2,
  102193.3,
  102187.3,
  102224.7,
  101975.4,
  101898.2,
  101832,
  101918.1,
  101835.5,
  102227.1,
  102556.6,
  102782.7,
  102729.7,
  102820.5,
  102799.8,
  102897.7,
  102955.5,
  103310.4,
  103460,
  103593.8,
  103649.1,
  103846.9,
  103733.4,
  103738.7,
  103465.6,
  103296.4,
  102902.4,
  102911.2,
  102692.7,
  102762.8,
  102786.1,
  102893.2,
  102851.1,
  103042.6,
  102990.7,
  102958,
  102587.2,
  102213.9,
  101859.6,
  101706.5,
  101270.9,
  101180.4,
  101232.2,
  101439.3,
  101451.9,
  101527.6,
  101521.6,
  101552.4,
  101432.6,
  101643.4,
  101868.4,
  102093.6,
  102171.5,
  102370.7,
  102434.2,
  102523,
  102542,
  102716,
  102739.9,
  102854.6,
  102810.4,
  102905.9,
  102936.4,
  103122.6,
  103014.4,
  102959.9,
  102802,
  102651.5,
  102038.6,
  101804.6,
  101626.1,
  101681.5,
  101592.9,
  101964.9,
  102610.1,
  103075.7,
  103203.9,
  103338.8,
  103342.7,
  103380.6,
  103088.9,
  103015.2,
  102764.1,
  102573.9,
  102175.9,
  102212.7,
  102156.3,
  102304.2,
  102164.7,
  102028,
  101862.9,
  101784.3,
  101527,
  101600,
  101742.4,
  102098.7,
  102363.8,
  102644.6,
  102760.1,
  102930.5,
  102671,
  102405.2,
  102132.5,
  101981.2,
  101876.4,
  102127.1,
  102361.6,
  102531.3,
  102406.9,
  102212.3,
  101875.4,
  101720.4,
  101462.6,
  101604.7,
  102008.2,
  102608.7,
  102910.2,
  103232.7,
  103135,
  103139.2,
  102762.4,
  102442.6,
  102097.4,
  101898.7,
  101648.7,
  101610.4,
  101636.9,
  101698.2,
  101498.1,
  101686.1,
  101833.9,
  102080.8,
  102145,
  102351,
  102471,
  102685.5,
  102788.3,
  102857.9,
  102706.3,
  102539.9,
  102206.4,
  102018.8,
  101879,
  101791.6,
  101431.2,
  101313.8,
  101215,
  101270.3,
  101305.1,
  101667.5,
  101950.4,
  102109.7,
  101856.7,
  101889.7,
  101909.7,
  101905.8,
  101836,
  102092.7,
  102199.7,
  102372.5,
  102471.3,
  102639,
  102598.3,
  102684.8,
  102515.5,
  102397,
  102379.1,
  102350,
  102034.7,
  101850,
  101734.4,
  101789.9,
  101755.2,
  101978.4,
  102204.9,
  102395.5,
  102300,
  102303.8,
  102357.9,
  102469.6,
  102343.6,
  102365.4,
  102204.5,
  102188,
  101869.2,
  101680.5,
  101532.5,
  101351.7,
  101112.3,
  101196.5,
  101236.6,
  101496.7,
  101660.4,
  101799.5,
  101961.8,
  102178.9,
  102108,
  102027.6,
  101893.6,
  101968.9,
  101717.5,
  101662.6,
  101615.8,
  101829.8,
  101767.2,
  102007.8,
  102242.9,
  101945.8,
  102140.2,
  102082.2,
  101775.4,
  101737,
  101430.6,
  101347.8,
  101356.3,
  101674.4,
  101933.7,
  102291,
  102474.5,
  102693.3,
  102654.3,
  102579.7,
  102310.7,
  102292,
  101871.1,
  101511.5,
  101382,
  101492.9,
  101353.3,
  101466.6,
  101472.1,
  101731.7,
  101818.8,
  101887.4,
  101700.9,
  101763.4,
  101531.1,
  101476,
  101553.2,
  101727.6,
  101775.1,
  102000.9,
  102091.1,
  102376.8,
  102371.5,
  102657.5,
  102864.6,
  103017.5,
  103199.2,
  103326.8,
  103301.3,
  103344.5,
  103223.1,
  102956.6,
  102888.4,
  102686.3,
  102414.2,
  102163.6,
  101959,
  101885,
  101590.4,
  101646.6,
  101750.7,
  101891.1,
  101882.9,
  102045.9,
  102190.1,
  102455.5,
  102530,
  102730,
  102851.5,
  102918.4,
  102905.1,
  102853.3,
  102814.6,
  102872,
  102615.2,
  102570.8,
  102358.1,
  102343.1,
  102121.3,
  102031.3,
  101934.4,
  102048.4,
  101918.4,
  101868.9,
  101787.6,
  101850.7,
  101666.6,
  101678.8,
  101732.6,
  101984.5,
  101887.6,
  101848.3,
  101933.6,
  102035.4,
  101864.7,
  101973,
  102063.5,
  102201.1,
  102121.6,
  102151.2,
  102102.5,
  102037.8,
  101758.7,
  101411.2,
  101184.9,
  101083.4,
  100836,
  100675.3,
  100708.8,
  100773.4,
  100582.1,
  100589.6,
  100584.9,
  100479.1,
  100636.3,
  101056.7,
  101316.3,
  101380.7,
  101249.2,
  101323.6,
  101397.8,
  101522.6,
  101630.8,
  101904.8,
  102098.6,
  102237.8,
  102022.3,
  101792.5,
  101619.8,
  101539,
  101335,
  101461.8,
  101773.1,
  102254.4,
  102194,
  102602.8,
  102528.1,
  102724.7,
  102744.9,
  102779,
  102714,
  102812,
  102677.5,
  102431.9,
  102208,
  102208.8,
  101728.1,
  101461.4,
  101519.6,
  101800.6,
  102018.9,
  102333.6,
  102445.4,
  102510.5,
  102232.5,
  102175.2,
  102010.9,
  101691.4,
  101383.9,
  101052.1,
  100965.5,
  101012.9,
  101077.5,
  101471,
  101748.6,
  102049.2,
  102346.9,
  102618.2,
  102795.7,
  102839.4,
  102861.8,
  102727.8,
  102735.2,
  102721.7,
  102429.9,
  102370.3,
  102289.7,
  102304.3,
  102110.5,
  102052.6,
  101978.9,
  102003.9,
  101807.3,
  101729.2,
  101361.8,
  101025.1,
  100958.1,
  101055.7,
  101149.8,
  101296.5,
  101344.4,
  101371.2,
  101369.5,
  101530.2,
  101513,
  101521.8,
  101561.8,
  101789.6,
  101833,
  101892.6,
  102015.5,
  102210.9,
  102243.7,
  102243.9,
  102274.2,
  102432.1,
  102257.8,
  102091.5,
  102032.2,
  102025,
  101705.5,
  101497.3,
  101470.8,
  101461.6,
  101006.2,
  100920.9,
  100892.6,
  101106.1,
  100924.4,
  101195.3,
  101397.7,
  101695.8,
  101662,
  101597.3,
  101681.3,
  101704.3,
  101695.1,
  101766.4,
  101749.8,
  101895.4,
  101716.7,
  101622.7,
  101648.6,
  101777.5,
  101617.9,
  101527.1,
  101523.7,
  101615.9,
  101429.9,
  101350.4,
  101416.8,
  101574.4,
  101473.3,
  101498.4,
  101475.5,
  101381.4,
  101043.1,
  100801.3,
  100687.7,
  100671,
  100480.5,
  100657.1,
  100725.9,
  101026.1,
  101251.5,
  101569.5,
  101578.2,
  101645.4,
  101462.4,
  101412.2,
  101346.2,
  101410.8,
  101057.7,
  100930.7,
  100849.6,
  100890.8,
  100998.2,
  101292.6,
  101429.9,
  101528.4,
  101447.6,
  101376.8,
  101241.3,
  101145.4,
  100870.3,
  100983.6,
  101393.1,
  101839.1,
  102005.2,
  102096.6,
  102102.3,
  102280.4,
  102071,
  101970.8,
  102032.9,
  102207,
  102019.9,
  101926.7,
  101919.5,
  102004.8,
  101860.5,
  101721.5,
  101679.8,
  101707.2,
  101109.5,
  101130,
  101044.1,
  101021.3,
  100566.8,
  100626,
  100676.4,
  100800.1,
  100560.5,
  100476.6,
  100597.4,
  100797.5,
  100877.5,
  101074.3,
  101213.3,
  101350.9,
  101664.5,
  101662.2,
  101747.1,
  101921.5,
  101875,
  101804.9,
  101839.4,
  101961.9,
  101689.3,
  101580.1,
  101393.1,
  101419.4,
  101124.6,
  101068.7,
  101037.1,
  101216,
  101192.8,
  101301.7,
  101293.8,
  101285.6,
  101033,
  100921.4,
  101079.5,
  101275.9,
  100943.9,
  100782.6,
  100865.1,
  100941.2,
  100814.2,
  101175.9,
  101436.3,
  101616.9,
  101379.6,
  101049.9,
  100919.8,
  100990.6,
  101104.5,
  101505.3,
  101619.7,
  101702.7,
  101457.1,
  101214,
  101182,
  101241.5,
  101008.9,
  100952.3,
  101184.7,
  101500.3,
  101405.4,
  101368.6,
  101418.7,
  101432.5,
  101038.7,
  100849.3,
  100803.5,
  100827.2,
  100575,
  100289.7,
  100357.5,
  100454,
  101008.8,
  101290.5,
  101209,
  101046.7,
  100741.8,
  100542.9,
  100645.7,
  101015.2,
  101192.1,
  101375.8,
  101536.4,
  101641.6,
  101640.3,
  101508.6,
  101450.9,
  101458.9,
  101210.4,
  101072.5,
  101111.3,
  101177.6,
  100910.4,
  100757.8,
  100861.8,
  101127.1,
  101281.7,
  101360,
  101361.6,
  101527.9,
  101525.8,
  101558.6,
  101670.1,
  101777.3,
  101652.2,
  101570.5,
  101637,
  101733.6,
  101571.3,
  101271.6,
  101272.3,
  101343.8,
  101028.9,
  100908.4,
  101010.8,
  101090.8,
  101006.4,
  100968.7,
  101034.5,
  101179.3,
  100897.8,
  100799.4,
  100852.9,
  100860.6,
  100498.2,
  100487.6,
  100704,
  100941.8,
  100974.3,
  101181.1,
  101346.2,
  101539.9,
  101615.3,
  101532.1,
  101591.3,
  101686.2,
  101593.5,
  101519,
  101449.2,
  101529.1,
  101423.5,
  101316.8,
  101381,
  101365.2,
  101004.1,
  100798.8,
  100690.6,
  100640.9,
  100604.4,
  100714.7,
  100794.4,
  100910.5,
  100718.5,
  100583.7,
  100476.7,
  100383.3,
  99963.34,
  99750.79,
  99851.88,
  100221.2,
  100385.4,
  100419.5,
  100349.9,
  100407,
  100027.2,
  99874.99,
  99744.36,
  99623.48,
  100175.7,
  100902.7,
  101360.8,
  101670.2,
  101805.1,
  101706.9,
  101743.2,
  101724.9,
  101390.2,
  101154.2,
  101096.4,
  101176.8,
  101034.5,
  100973.9,
  101114.2,
  101286.5,
  101238.5,
  101201.2,
  101147.1,
  101167.9,
  100943.3,
  100799.3,
  100731.3,
  100730.6,
  100450.4,
  100509.3,
  100688.2,
  100864.2,
  100708.2,
  100869.4,
  100687.2,
  100737.6,
  100289.1,
  100285.5,
  100280.3,
  100414.1,
  100374.5,
  100465.2,
  100572.4,
  100845.3,
  100905.4,
  100901.2,
  100799,
  100733.1,
  100515.8,
  100433.2,
  100418.4,
  100602.8,
  100553,
  100733.4,
  100856.7,
  101075.9,
  101146.2,
  101223.7,
  101320,
  101481.1,
  101276.4,
  101203.7,
  101172.7,
  101327,
  101098.2,
  100973,
  101018,
  101119.1,
  100822.9,
  100821.8,
  101022,
  101223.8,
  101124.1,
  101149.3,
  101211.4,
  101388.3,
  101039.9,
  101049.5,
  100974.1,
  100944.2,
  100681.3,
  100723.8,
  100847.1,
  101187.3,
  101315.8,
  101410.5,
  101483.6,
  101660.9,
  101613.2,
  101537.3,
  101599.4,
  101681.8,
  101469.6,
  101349.8,
  101414.1,
  101458,
  101158.6,
  101080,
  101059.4,
  101035,
  100845.4,
  100898.1,
  100964.8,
  101208.1,
  101216.2,
  101345.5,
  101368.6,
  101620.3,
  101550.2,
  101562,
  101625.7,
  101772.7,
  101721.3,
  101508.4,
  101472.9,
  101611.4,
  101058.1,
  101057.3,
  100840.2,
  100985.3,
  100925,
  101151,
  101255,
  101426.7,
  101400.9,
  101345.2,
  101348.8,
  101453.4,
  101278.1,
  101201.6,
  101224.7,
  101380.3,
  101199.3,
  101230,
  101378.3,
  101568.4,
  101468.3,
  101456.1,
  101605.4,
  101599.5,
  101285.3,
  101162.3,
  101192.4,
  101169.1,
  100781.2,
  100726.3,
  100688.3,
  100680.4,
  100500.3,
  100362.9,
  100266.3,
  100356.1,
  100330.3,
  100341.3,
  100511.9,
  100705,
  100701.7,
  100842.7,
  100959.8,
  101026.5,
  100863.6,
  100815.3,
  100858.8,
  100928.6,
  100888.4,
  100931.4,
  101071.8,
  101038.3,
  100646.9,
  100353.2,
  100345.2,
  100637.6,
  100642.5,
  101011.2,
  101330.8,
  101515.7,
  101461,
  101506.9,
  101556.4,
  101655.6,
  101674.2,
  101836.5,
  101883.2,
  102041.8,
  101941.4,
  101863.8,
  101835.8,
  101938.6,
  101710.3,
  101652.5,
  101776.2,
  101792.7,
  101677.3,
  101679.1,
  101779,
  101921.9,
  101689,
  101512.1,
  101530,
  101563.5,
  101314.6,
  101166.6,
  101225.8,
  101310.2,
  101065.2,
  100906.8,
  101014.7,
  100982.3,
  100525.1,
  100266.9,
  100169.1,
  100149.6,
  99895.59,
  100012.6,
  100168.8,
  100491,
  100801.3,
  101085.5,
  101255.6,
  101422.6,
  101670.1,
  101800.7,
  102014.7,
  102145,
  102092.3,
  102080.4,
  102073.1,
  102224.7,
  101990.4,
  101821.8,
  101810.6,
  101882.9,
  101666.1,
  101512.9,
  101591.9,
  101716.9,
  101483.4,
  101431.2,
  101440,
  101524.7,
  101342.4,
  101259,
  101180.1,
  101217.4,
  101022.2,
  100918.2,
  100896.7,
  100993.5,
  100836.3,
  100943.3,
  100949.3,
  100986.1,
  100814.1,
  100736,
  100713.1,
  100761.1,
  100713.7,
  101235.6,
  101378.1,
  101582.4,
  101384.3,
  101325.7,
  101321,
  101269.5,
  100914.3,
  100686.3,
  100564.6,
  100754.8,
  101286.1,
  101774.3,
  101917.1,
  102206.6,
  102310.2,
  102276.4,
  102249.7,
  102450.4,
  102348.7,
  102340.9,
  102330.4,
  102538.7,
  102349,
  102243.1,
  102304,
  102511.3,
  102263.6,
  102195.6,
  102207.8,
  102375.1,
  102246.2,
  102236.3,
  102331.2,
  102539.9,
  102420.8,
  102380.8,
  102451.7,
  102469.6,
  102295,
  102148.3,
  102049.4,
  102026.2,
  101707.4,
  101572.4,
  101515.7,
  101588.7,
  101495.4,
  101461.4,
  101538.6,
  101716.6,
  101517.4,
  101583.3,
  101734.1,
  101851.6,
  101582.1,
  101787.7,
  101701.2,
  101784.3,
  101604.6,
  101646.9,
  101637.4,
  101648.8,
  101590.1,
  101590.1,
  101711.2,
  101713.2,
  101634.4,
  101701.9,
  101678.2,
  101852.3,
  101795.1,
  101766.2,
  101746.9,
  101840.2,
  101604.7,
  101490.5,
  101469.1,
  101508.3,
  101420.3,
  101561.9,
  101757.7,
  102104.4,
  102163.9,
  102425.6,
  102647.5,
  102843.9,
  102890.2,
  102871.2,
  102908.8,
  102995.5,
  102834.1,
  102683.4,
  102629.4,
  102704.1,
  102531.8,
  102517.8,
  102514,
  102671.5,
  102540.8,
  102542.3,
  102557.4,
  102644.6,
  102492.1,
  102463,
  102411.5,
  102494,
  102285.2,
  102243.1,
  102217.3,
  102346.4,
  102139.1,
  102101.3,
  102015,
  102035.6,
  101854.9,
  101827.1,
  102094.4,
  102191.4,
  102341.1,
  102495.7,
  102509.2,
  102622.2,
  102446.2,
  102332.8,
  102242.2,
  102266.9,
  102018,
  101986.4,
  101925.3,
  101867.2,
  101570.1,
  101472,
  101359.6,
  101461.1,
  101279.4,
  101305.3,
  101323.6,
  101492.2,
  101381.5,
  101393.4,
  101391.4,
  101422.4,
  101292.8,
  101434.9,
  101495.7,
  101684.8,
  101695.4,
  101697,
  101631.6,
  101635.2,
  101234.4,
  101263.2,
  101343.9,
  101305.6,
  101262.6,
  101370.8,
  101221.5,
  101457.7,
  101187.2,
  101313.6,
  101263.7,
  101161.1,
  101076.2,
  101518.1,
  101815.3,
  102071.9,
  102305.6,
  102401.6,
  102615.8,
  102832.1,
  102672.4,
  102678.8,
  102559,
  102629.2,
  102488,
  102400.7,
  102267.7,
  102173.5,
  101804,
  101641.5,
  101381.1,
  100945,
  100658.5,
  101027.9,
  101300.1,
  101605.8,
  101856.6,
  102122.2,
  102193.1,
  102223.5,
  102087,
  101946.6,
  101888,
  101819.8,
  101652.5,
  101710.6,
  101860.5,
  101971.9,
  101801.7,
  101820.6,
  101644.6,
  101537.9,
  101327.2,
  101322.7,
  101230.3,
  100976.8,
  100558.3,
  100283,
  100310.7,
  100777.7,
  100843.6,
  100826.9,
  100770.2,
  100932.2,
  101127.4,
  101363.1,
  101494.3,
  101713.6,
  101862.3,
  102122.4,
  102094.5,
  102142.2,
  102057,
  101909.6,
  101893.1,
  101884.9,
  101794.3,
  101925.6,
  102032.4,
  102222.5,
  102153.1,
  102231.4,
  102245.3,
  102273.8,
  102128.1,
  101991.2,
  101934.9,
  101959.4,
  101781.2,
  101768.5,
  101660.7,
  101592,
  101309.3,
  101196.2,
  101122.3,
  101657.2,
  101618.5,
  101948.2,
  102127,
  102385.2,
  102425.2,
  102592.8,
  102591.8,
  102815.9,
  102888.4,
  103052.4,
  103067.1,
  103096.7,
  103094.3,
  103081.9,
  102986.7,
  102956.2,
  102776.9,
  102692.1,
  102616.1,
  102675.9,
  102659.2,
  102809.9,
  102810.9,
  102897.1,
  102675.8,
  102654.2,
  102553.7,
  102538.2,
  102265.4,
  102188.7,
  102051.5,
  101864.3,
  101636.2,
  101671,
  101598,
  101590.4,
  101315.6,
  101154,
  100976.4,
  100830.5,
  100332.2,
  100060.5,
  99970.45,
  100327.4,
  100452.1,
  100901.5,
  101261,
  101531,
  101574.7,
  101502,
  101251.4,
  101001.8,
  100593.2,
  100500.9,
  100349,
  100112,
  99622.17,
  99683.95,
  99249.06,
  99319.91,
  100947.3,
  101932.3,
  102295.2,
  102615,
  102879.4,
  103147.8,
  103245.3,
  103391.1,
  103408.4,
  103386.9,
  103199.5,
  103018.3,
  102601.2,
  102546,
  102430.8,
  102454.2,
  102408.6,
  102521.3,
  102487.2,
  102516.6,
  102376,
  102343.3,
  102239.4,
  102191.6,
  101990.4,
  102020.4,
  102011.5,
  102075.8,
  101975.3,
  101971.4,
  101900.8,
  101853.7,
  101586.4,
  101632.3,
  101697,
  101721.8,
  101646.5,
  101830.4,
  102018.4,
  102135.5,
  102074.8,
  102092.2,
  101933,
  101977,
  101829.9,
  101880.7,
  101811,
  101890.2,
  101622.5,
  101575.8,
  101561.4,
  101583.6,
  101293.5,
  101344.4,
  101418.5,
  101484.2,
  101093.5,
  101391.2,
  101743.3,
  102174.6,
  102393.5,
  102797.6,
  102977.8,
  103182.1,
  103181.6,
  103195.8,
  103087.7,
  102931.5,
  102632,
  102549,
  102427.8,
  102460,
  102134.9,
  102113.1,
  101875.7,
  101615.4,
  101079.8,
  100774.3,
  100394.9,
  100146.8,
  99902.63,
  100039,
  100090.2,
  100178.7,
  99946.8,
  99913.74,
  99743.57,
  100034.6,
  99946.65,
  100438.7,
  100686.7,
  101060.9,
  101411.6,
  101548.4,
  101377.8,
  101047.1,
  100694.4,
  100739.8,
  101059.2,
  101169.6,
  100728.2,
  100618.2,
  100541.9,
  100719.7,
  101280.7,
  101759,
  101914.6,
  102128.9,
  102152.1,
  102126.8,
  101957.9,
  101878.9,
  101597.1,
  101555.2,
  101521.1,
  101503.3,
  101309.8,
  101337.4,
  101159.3,
  101361.8,
  101625.4,
  102051.3,
  102232.4,
  102327.7,
  102265.8,
  102289.4,
  102128,
  102063.2,
  101537.7,
  100841.6,
  100153.9,
  100073,
  100798.5,
  101680.2,
  101896.2,
  101992.5,
  101823,
  101942.7,
  101968.3,
  101989.6,
  102045,
  102134.8,
  102104.5,
  102104,
  101939.1,
  101988.6,
  102057.8,
  102134.3,
  101974,
  101863.3,
  101705.3,
  101664.1,
  101555,
  101746.7,
  101786.1,
  101849.3,
  101866,
  101992.7,
  101998.9,
  102033.8,
  101987.5,
  101959,
  101840.2,
  101919.3,
  101871.3,
  102120.4,
  102328,
  102485.7,
  102380.5,
  102380.9,
  102313,
  102344.3,
  102304.7,
  102597.2,
  102730.7,
  102828.7,
  102863.6,
  102855.5,
  102680.8,
  102673,
  102385.5,
  102334.1,
  102270.2,
  102308.7,
  101985.8,
  101836.2,
  101686.2,
  101597.1,
  101427.1,
  101656,
  101769.5,
  102067.8,
  102518.8,
  102996.4,
  103155,
  103365.5,
  103374.7,
  103467.1,
  103407.7,
  103473.6,
  103357.4,
  103321,
  103244.6,
  103198.3,
  103047.8,
  103021,
  102995.7,
  103016,
  102787.8,
  102751.4,
  102668.1,
  102417.6,
  102118,
  102115.2,
  102092.5,
  102152,
  102070.5,
  102177.2,
  102176.8,
  102084.5,
  101822.2,
  101696.7,
  101576.8,
  101467.5,
  101232.2,
  101233.4,
  101172.2,
  100852,
  100197.8,
  100554.3,
  101390.9,
  101713.6,
  101775.3,
  102037.3,
  102145.8,
  102197,
  102010,
  102003.6,
  102060.4,
  102314,
  102576.8,
  103143.1,
  103521.7,
  103935.9,
  104132.4,
  104327.9,
  104267,
  104339,
  104224.5,
  104113.5,
  103891.6,
  103894,
  103574.6,
  103409.2,
  103208.6,
  103132.6,
  102768.3,
  102621.9,
  102592.9,
  102629.1,
  102424.4,
  102559,
  102651.9,
  102797.6,
  102871.4,
  103102.2,
  103203.7,
  103268.9,
  103158.9,
  103041.3,
  102791,
  102582.6,
  102193.1,
  102024.3,
  102041.6,
  102195.3,
  102100.3,
  102076.7,
  101802.8,
  101672.3,
  101995,
  102636.4,
  102785.6,
  103027.1,
  103001.4,
  102865,
  102546.5,
  102352.4,
  101761.8,
  101448.6,
  101357.7,
  101511.8,
  101644.7,
  102003.3,
  102171.3,
  102337.1,
  102312.5,
  102339.1,
  102289.2,
  102259.7,
  102030,
  101845.1,
  101639.6,
  101523.1,
  101317.5,
  101520.5,
  101795.1,
  102243,
  102451.4,
  102679.7,
  102697.6,
  102757.2,
  102628.1,
  102697,
  102713.3,
  102829.1,
  102683.5,
  102673.2,
  102461.2,
  102287.2,
  101865.9,
  101753.8,
  101674.1,
  101904.6,
  101952.5,
  102208.5,
  102263.4,
  102485,
  102528.4,
  102662.5,
  102668.4,
  102825.5,
  102809.6,
  102825.1,
  102775.4,
  102810.6,
  102534.1,
  102378.3,
  102188.5,
  101999.4,
  101653.1,
  101639.4,
  101965.3,
  102676.3,
  102906.3,
  103115.9,
  102997.3,
  103054.4,
  102748.6,
  102523.9,
  102345,
  102209,
  101923.2,
  101845.4,
  101939,
  102311.5,
  102536.9,
  102749.2,
  102690.6,
  102711.3,
  102132.2,
  101851.2,
  101683.6,
  101549.3,
  101101,
  101049.5,
  101676.3,
  102282.6,
  102371.4,
  102879,
  103124.4,
  103375.6,
  103426.3,
  103492.7,
  103424,
  103503.2,
  103205,
  103019.8,
  102923.6,
  102994.9,
  102784.2,
  102735.8,
  102622.6,
  102609.8,
  102322.6,
  102202.4,
  102066,
  102039.1,
  101867.8,
  101917,
  101857.3,
  101842.9,
  101575.2,
  101377.4,
  101334.2,
  101335.4,
  101228.6,
  101521.8,
  101775.9,
  101864.3,
  101511.1,
  101323.3,
  101255.7,
  101416.2,
  101294.2,
  101538.5,
  101748.5,
  101862.2,
  101831.5,
  101870,
  101806.2,
  101765.1,
  101624.5,
  101814.8,
  102061.7,
  102400.6,
  102487.6,
  102716.6,
  102558.7,
  102423.4,
  102268.9,
  102289.4,
  102229.8,
  102286.8,
  102150.9,
  102109.8,
  101879.8,
  101751.6,
  101678.8,
  101666.3,
  101643.5,
  101749.5,
  101555.9,
  101507.1,
  101436.5,
  101641.2,
  101415.8,
  102116.5,
  102262.2,
  102831.6,
  102927.9,
  103134.3,
  103026.7,
  103084.8,
  102974.6,
  102948.9,
  102848.2,
  102798.3,
  102500.8,
  102383.1,
  102164.2,
  102101.7,
  101726.1,
  101601.2,
  101378.4,
  101632.6,
  101441.7,
  101642,
  101985.3,
  102336.4,
  102342.5,
  102388.2,
  102382.1,
  102340.5,
  101970.4,
  101742.7,
  101705.2,
  101882.6,
  101970.8,
  102316.7,
  102334.1,
  102140.3,
  102019.1,
  101467,
  101146.6,
  101025.6,
  101138.2,
  101543.8,
  101766.4,
  101894.6,
  101793,
  101676.7,
  101546.1,
  101150.2,
  101116,
  101112.5,
  101135,
  101306.4,
  101367.5,
  101594.2,
  101728.1,
  101807.8,
  102105.1,
  102208.1,
  102198.7,
  102387.2,
  102301,
  102255.8,
  102245.2,
  102394.6,
  102279.9,
  102302.1,
  102239.6,
  102253.8,
  101942.5,
  101815.4,
  101639.7,
  101832.7,
  101719.3,
  102092.8,
  102330.5,
  102468.8,
  102477.7,
  102186.5,
  101864.2,
  101487.5,
  101248.8,
  101341.8,
  101540.2,
  101677.5,
  101752.8,
  101777.2,
  101779.7,
  101894.4,
  101625.7,
  101636.4,
  101582.9,
  101856.9,
  101966.3,
  102160.3,
  102201.3,
  102304.5,
  102111.8,
  101974.8,
  101697.7,
  101642.3,
  101332.4,
  101146.3,
  101044.9,
  101335.7,
  101846.9,
  102339.9,
  102390.8,
  102595.6,
  102559.9,
  102533.5,
  102414.1,
  102466,
  102175.3,
  101959.5,
  101837.6,
  101616,
  101086.5,
  100914.4,
  101196,
  101483.3,
  101578.7,
  101478.9,
  101473,
  101444.8,
  100924.1,
  100701.1,
  100782,
  100986,
  101405.4,
  101175.7,
  101666.3,
  101773.9,
  101828.1,
  101869.3,
  101964.5,
  102138.6,
  102103.6,
  102159.8,
  102262.4,
  102414.6,
  102431.6,
  102397.3,
  102367.7,
  102486.7,
  102322.5,
  102230.6,
  102302.6,
  102428.4,
  102324.6,
  102328.9,
  102345,
  102421.1,
  102173,
  102143.2,
  101899,
  101818.4,
  101382.3,
  101122.8,
  100952.1,
  100942.3,
  100713.8,
  100819.7,
  100844.1,
  101088,
  101015.8,
  101182.6,
  101329.1,
  101424.5,
  101474.3,
  101690,
  101976,
  102258.5,
  102158.7,
  101992.9,
  101904.4,
  101854.9,
  101521.7,
  101328.9,
  101308.8,
  101320.8,
  101041,
  101052.8,
  101186.4,
  101314.1,
  101279.5,
  101325.3,
  101465.2,
  101715.9,
  101605.6,
  101586.3,
  101560.6,
  101608.7,
  101343.2,
  101268.6,
  101211.6,
  101265.3,
  101059.6,
  101078.3,
  101176.3,
  101286,
  101468,
  101436,
  101465.2,
  101655.2,
  101449.9,
  101299.9,
  101186.3,
  101197.9,
  100968.5,
  101093.3,
  101175.9,
  101271.7,
  101297.4,
  101305.7,
  101287.6,
  101386.2,
  101248.1,
  101265.5,
  101295.8,
  101348.1,
  101281.7,
  101220.6,
  101288.4,
  101465.8,
  101457,
  101474.9,
  101614.5,
  102003.9,
  102021.9,
  102211.5,
  102185,
  102435.7,
  102291.9,
  102081.2,
  102018.5,
  101978.7,
  101621.8,
  101405.3,
  101152.7,
  101145.5,
  100951.8,
  101125.5,
  101507.1,
  101847,
  101884.6,
  101796.8,
  101805.1,
  101811.9,
  101398.3,
  101391.3,
  101123.7,
  100993.9,
  100478.7,
  100269.7,
  100388.5,
  100624.4,
  100576.7,
  100631.4,
  100657,
  100810.2,
  100883.2,
  101182.4,
  101365.8,
  101368.3,
  101056.9,
  100915.1,
  100750.6,
  100880.4,
  100890.2,
  101149.9,
  101426,
  101859.2,
  102199.1,
  102317.5,
  102352.7,
  102539.5,
  102460.1,
  102343.9,
  102357.5,
  102444,
  102074.5,
  101780.8,
  101648,
  101610.7,
  101280.8,
  101089.2,
  100997.5,
  100952,
  100605.6,
  100300.2,
  100492.4,
  101079.9,
  101370.1,
  101509,
  101703.4,
  101868.1,
  101704.4,
  101521,
  101445.3,
  101161,
  100652.4,
  100438.3,
  100406.1,
  100923.8,
  101297.4,
  101292.7,
  101316.2,
  101471.5,
  101327.3,
  101471.5,
  101491.8,
  101626,
  101567.3,
  101559.7,
  101498.7,
  101599.7,
  101529.1,
  101510.7,
  101489.8,
  101495.6,
  101115.1,
  100862.1,
  100662.9,
  100523.9,
  100303.1,
  100492.7,
  100883.6,
  101167.2,
  101020.3,
  100809.1,
  100697.5,
  100701.8,
  100567.1,
  100475.6,
  100596.8,
  100713.4,
  100474.2,
  100170.3,
  99958.43,
  99965.56,
  99886.99,
  100313.3,
  100574.1,
  100609.6,
  100256.6,
  99843.55,
  99794.81,
  99883.15,
  99952.8,
  100308.7,
  100481.8,
  100941.1,
  101158.3,
  101264.5,
  101458.7,
  101456.7,
  100999.8,
  100681.7,
  100752.1,
  101140.1,
  101511.3,
  101593.3,
  101447.5,
  101311.1,
  100906.6,
  100410.6,
  100425.7,
  101101.1,
  101349.1,
  101529.7,
  101775.3,
  101979.3,
  101898.7,
  101955.1,
  101961.2,
  102005.9,
  101910.2,
  101858.1,
  101850.1,
  101923.1,
  101662.9,
  101404.7,
  101428.5,
  101376.7,
  100939.8,
  100793,
  100812.7,
  100907.5,
  100590.4,
  101034.2,
  101060.2,
  101187.3,
  101049.6,
  100982.4,
  101112.7,
  101382,
  101330.8,
  101277.2,
  101433.2,
  101511.7,
  101305.4,
  101139.3,
  101013,
  100637,
  100218,
  100613.9,
  101000.4,
  101297.6,
  101461.9,
  101508.4,
  101532.3,
  101618,
  101305.5,
  101174.7,
  101322.1,
  101499.5,
  101416.9,
  101512.3,
  101539.5,
  101634.3,
  101823.4,
  101999.4,
  102142.8,
  102245.8,
  102207.1,
  101993.5,
  101902.6,
  101826.2,
  101449.4,
  101154.8,
  101216.7,
  101294.5,
  101115.1,
  101070.3,
  101108.1,
  101282.2,
  101471.1,
  101469.7,
  101525.4,
  101629.3,
  101586.9,
  101527.3,
  101497.3,
  101482.2,
  101257.2,
  101046.5,
  100957.7,
  100880.9,
  100841.3,
  100969.1,
  101024.2,
  100847.4,
  100921.7,
  101053.4,
  101163.6,
  101519.3,
  101600.4,
  101776.8,
  101608.6,
  101715.9,
  101460.3,
  101227,
  100862,
  100481.1,
  100317.4,
  100580.6,
  100846.6,
  101224.1,
  101611.3,
  101826.4,
  101987.2,
  102279.4,
  102557.5,
  102562.6,
  102544.8,
  102651.5,
  102432.8,
  102185.1,
  101957.9,
  101997.6,
  101636.3,
  101409.4,
  101463.6,
  101522.6,
  101441.5,
  101402.7,
  101467.4,
  101657,
  101565,
  101451.9,
  101440.8,
  101489.2,
  101372.7,
  101282.8,
  101230.6,
  101329.9,
  101039.8,
  101051.4,
  100967.1,
  101134.6,
  101052,
  101166.5,
  101152.8,
  101310.5,
  101183.5,
  101237.1,
  101134.5,
  101199.3,
  101031.4,
  100995.6,
  101031.9,
  101158.8,
  101083,
  100851.2,
  100878,
  100814.1,
  100681.7,
  100699.5,
  100959.6,
  100910.1,
  100948.5,
  100964.4,
  101103.5,
  101293.6,
  101473.4,
  101454.2,
  101580.1,
  101798.1,
  101842.6,
  101758.4,
  101829.4,
  101967.3,
  101745.1,
  101621.9,
  101724.4,
  101805.7,
  101541.1,
  101543.1,
  101589.1,
  101651.4,
  101490.7,
  101374.4,
  101435.9,
  101508.3,
  101365.3,
  101290.5,
  101321.8,
  101483.8,
  101419.2,
  101419.9,
  101424.3,
  101602.6,
  101564.5,
  101453,
  101417.2,
  101544.2,
  101457,
  101439.4,
  101456.9,
  101623.2,
  101509.3,
  101473,
  101467,
  101501.1,
  101301.1,
  101185.2,
  101172.2,
  101162.4,
  100971.4,
  100951.1,
  100985.7,
  101067.2,
  101024.4,
  101039.3,
  101067,
  101141.9,
  101006.2,
  101076.4,
  101030.6,
  101076.4,
  100878.2,
  100861,
  100771.7,
  100829.9,
  100778.1,
  100907.9,
  100995.3,
  101214.4,
  101360.2,
  101599.5,
  101642.5,
  101730,
  101741.9,
  101690.2,
  101717.8,
  101831.2,
  101679.1,
  101611.2,
  101715.1,
  101881.6,
  101850.3,
  101886.1,
  101926.2,
  102136.4,
  102095.5,
  102059.2,
  101996,
  102070.9,
  101875.4,
  101671.1,
  101566,
  101563.5,
  101290.7,
  101194.1,
  101146.3,
  101217.5,
  101040.9,
  101012.1,
  101033.8,
  100978.5,
  100606.3,
  100485,
  100665.3,
  101140.4,
  101292.3,
  101402.2,
  101383.1,
  101396.4,
  101515.7,
  101928.3,
  101858.9,
  101984.5,
  101978.2,
  101822.7,
  101773.6,
  101873.3,
  101532.4,
  101554.4,
  101555,
  101585.9,
  101392.6,
  101371,
  101343.2,
  101368.7,
  101412.4,
  101397.4,
  101295.4,
  101374.8,
  101394.4,
  101559.8,
  101638.5,
  101774.7,
  101868,
  101877.1,
  101836.6,
  101985.2,
  101930.2,
  101837.5,
  101844.4,
  101878,
  101726.6,
  101560.3,
  101523.6,
  101555.8,
  101372.6,
  101469.5,
  101488.9,
  101659.4,
  101544.2,
  101498.1,
  101441.6,
  101461.8,
  101213.6,
  101158.9,
  101128.7,
  101133.4,
  100939,
  100872.1,
  100948.4,
  101200.7,
  101257.1,
  101260.6,
  101205.9,
  101384.2,
  101081.8,
  100768.9,
  100721.7,
  100679.2,
  100656.4,
  100883.2,
  101005.3,
  101083.8,
  100925,
  100726.9,
  100498.3,
  100343.8,
  100124.5,
  100133.3,
  100335.9,
  100772.1,
  100808.5,
  101268.1,
  101354.6,
  101623.7,
  101637.1,
  101546.3,
  101443.6,
  101326.9,
  100844.7,
  100919.3,
  101130.6,
  101275.5,
  100982.7,
  101038.4,
  100971.5,
  100995,
  100612.4,
  100514.1,
  100535.7,
  101250.1,
  101326,
  101672.6,
  101821.7,
  102023.2,
  102039.4,
  102063.5,
  102108.9,
  102199.4,
  102096.5,
  101982.5,
  101894.7,
  102063.2,
  101804.6,
  101624.7,
  101628.2,
  101695.9,
  101412.7,
  101404.6,
  101503.8,
  101680.6,
  101586.4,
  101660.9,
  101564.6,
  101788.3,
  101481.8,
  101536,
  101412.1,
  101500.2,
  101331.2,
  101108.9,
  101058.4,
  101159.9,
  100995.4,
  101217.6,
  101389.8,
  101736.2,
  101884.7,
  102061.5,
  101996.7,
  102024.1,
  101874.1,
  101817.9,
  101659.6,
  101801.5,
  101810.5,
  101903.5,
  101985.3,
  102050.6,
  101961.9,
  101966.8,
  101872.4,
  101805.1,
  101520.3,
  101444.1,
  101391.1,
  101417.5,
  101194.5,
  101198.5,
  101114.6,
  101188.2,
  101029.8,
  101022.4,
  101091.2,
  101274.6,
  101336.3,
  101710.9,
  101938.5,
  102114.2,
  102130.5,
  102106.9,
  101990.3,
  102077.8,
  101942.1,
  101815.1,
  101651.2,
  101724.8,
  101413.1,
  101256.1,
  101059.3,
  101061.5,
  100837.1,
  100860,
  101067.1,
  101338.4,
  101424.1,
  101506.5,
  101511.9,
  101733.7,
  101711.1,
  101853,
  101821.7,
  101934.2,
  101953.2,
  102077.3,
  102013.1,
  102095.3,
  102090.3,
  102159.8,
  102189.9,
  102282.1,
  102149,
  102116.9,
  102078.7,
  102181.3,
  101963.3,
  101880.9,
  101813.8,
  101765.1,
  101613.6,
  101593.6,
  101596.3,
  101754.7,
  101702.7,
  101833,
  101816.8,
  102002,
  101842.3,
  101759.2,
  101653.6,
  101696.5,
  101787.8,
  101920.9,
  101997.8,
  102181.5,
  102327.7,
  102552.1,
  102656.1,
  102860.8,
  102911.5,
  102950.1,
  102946,
  103116.9,
  103012.4,
  102928.7,
  102849.8,
  102945.4,
  102686.9,
  102595.2,
  102554,
  102611.3,
  102349.8,
  102283.5,
  102248.9,
  102310.7,
  102142.5,
  102105.5,
  102134.1,
  102186.8,
  102073.7,
  102074.6,
  102125.5,
  102203.8,
  102081,
  102120.6,
  102168.7,
  102291.2,
  102210.1,
  102236.8,
  102271.1,
  102324.1,
  102192.7,
  102104.6,
  102080.2,
  102141.5,
  101960.8,
  101740.3,
  101625.9,
  101781.9,
  101747.8,
  101875.8,
  101867,
  101958.6,
  101848.4,
  101805.5,
  101564.2,
  101314.9,
  101192.1,
  101506.6,
  101971.7,
  102249.6,
  102462.1,
  102761.8,
  102743.7,
  102914,
  102945.7,
  102981.2,
  102950.1,
  102986,
  102924.7,
  102857.3,
  102623.3,
  102545.5,
  102215.5,
  102003.3,
  101890.6,
  101870.4,
  101712.5,
  101769.3,
  101769.6,
  101808.4,
  101706.1,
  101738.3,
  101673.4,
  101640.8,
  101410.4,
  100889.2,
  100824.8,
  101132.9,
  101149.6,
  101167.3,
  101410.6,
  101592.8,
  101606.2,
  101870.1,
  101947.2,
  102128,
  101986.4,
  102042,
  101907.9,
  102009.6,
  101776.9,
  101636.2,
  101468.1,
  101355.9,
  100982.9,
  101033.7,
  101148.9,
  101637.6,
  101865.4,
  102148.6,
  102232.9,
  102367,
  102273.1,
  102248.3,
  102072.1,
  102082.6,
  101998.2,
  102223.2,
  102348.4,
  102584,
  102593.3,
  102654.4,
  102585.3,
  102558,
  102637.8,
  102659.7,
  102593.2,
  102638.5,
  102408.9,
  102241,
  102103,
  102034.4,
  101738.6,
  101601.8,
  101473.4,
  101391.9,
  101483,
  101847.6,
  102235.9,
  102435.9,
  102543.7,
  102657.3,
  102594.3,
  102578.6,
  102346.7,
  102337.8,
  102118.7,
  102038.1,
  101700.6,
  101614.3,
  101421.3,
  101472.4,
  101211.8,
  101230.1,
  101296.5,
  101698.3,
  102167.3,
  102559.9,
  102662,
  102789,
  102777,
  102767.6,
  102625.2,
  102552,
  102262,
  102207.7,
  102036.7,
  102011.4,
  101754.9,
  101792.9,
  101801.6,
  101795.6,
  101629,
  101655.2,
  101574,
  101439.5,
  101410.1,
  101496.8,
  101414.9,
  101377.8,
  101391.6,
  101708,
  101854.4,
  102048.9,
  102025.3,
  102159.5,
  102032.2,
  102138.5,
  101935.6,
  101984,
  101915.4,
  101966.6,
  101806.4,
  101827.4,
  101729,
  101733.2,
  101534.8,
  101471.2,
  101357.5,
  101596.8,
  101616.5,
  101663.6,
  101665.8,
  101754.3,
  101700,
  101583,
  101418.2,
  101256.5,
  101124.6,
  101103.7,
  101102.1,
  101229.3,
  101106,
  100928.3,
  100576.1,
  100515.6,
  100493.2,
  100705.4,
  100601.7,
  100891.2,
  101035.2,
  101355.1,
  101442.9,
  101605.8,
  101577.7,
  101759.9,
  101610.5,
  101782.8,
  101886.2,
  102187.9,
  102576,
  102850.5,
  103080.5,
  103302.9,
  103302.5,
  103397.6,
  103406.8,
  103458.9,
  103279.6,
  103301.9,
  103103.2,
  103182.9,
  103049.6,
  103083.8,
  102991.5,
  103033.3,
  102927.5,
  102919.8,
  102755,
  102728.1,
  102549.5,
  102540.7,
  102417.8,
  102483.6,
  102489.8,
  102444.7,
  102368.6,
  102234.7,
  101866,
  101550.6,
  101046.7,
  100989,
  101113.3,
  101409.1,
  101496.2,
  101589,
  101539.9,
  101504.5,
  101341.6,
  101445.9,
  101571.7,
  101651.1,
  101495.4,
  101450.6,
  101340.8,
  101446.2,
  101419.4,
  101452.1,
  101300.3,
  101137.1,
  100928.2,
  100613.3,
  100199.3,
  100695.5,
  100655.1,
  100513.7,
  100304.6,
  100774.2,
  100648.1,
  100789.8,
  100700,
  101066.4,
  101282.9,
  101605.1,
  101645.8,
  101750.4,
  101763.8,
  102052,
  102114.2,
  102135.2,
  102061,
  102051.6,
  101738.8,
  101519.3,
  101576.2,
  101636.2,
  101601.1,
  101676.2,
  101574,
  101603.5,
  101527.7,
  101501.2,
  101494.2,
  101687.5,
  101807.1,
  101875.3,
  101868.8,
  101997.1,
  102139.5,
  102059.5,
  101889.1,
  102099.6,
  102074,
  102113.9,
  102080.7,
  102202.5,
  102215.6,
  102287.3,
  102363.8,
  102625.7,
  102723.5,
  102886.1,
  102950.6,
  103066.3,
  102899.4,
  102796.2,
  102488,
  102263.4,
  102009.1,
  101863.4,
  101574.4,
  101713.3,
  101822.4,
  102032.1,
  102225.4,
  102562.5,
  102729,
  103084.9,
  103143.5,
  103189,
  102959.3,
  102987.5,
  102746.6,
  102326.6,
  101917.6,
  101618,
  101372,
  101328.8,
  101228.7,
  101255.2,
  101077.2,
  101209.7,
  101172.1,
  101101,
  101784.2,
  102399.3,
  102507.4,
  102628,
  102455.9,
  102391.7,
  102057.2,
  101911.4,
  101669.6,
  101900.7,
  102041.7,
  102255.3,
  102278.3,
  102332.3,
  102140.5,
  101861.1,
  101505.6,
  101587.9,
  101787.8,
  102008.7,
  102015.6,
  102177.7,
  102179.4,
  102291.3,
  102269.4,
  102284.7,
  102199.8,
  101782.6,
  101400.2,
  101709.1,
  102191.6,
  102558.7,
  102681.5,
  102835.9,
  102928.2,
  102943.2,
  102716.4,
  102493.4,
  102202.2,
  101966.5,
  101762.8,
  101826,
  101933.8,
  102123.7,
  102151,
  102366.2,
  102484.6,
  102593.2,
  102603.6,
  102738.9,
  102717,
  102753,
  102631.3,
  102699.2,
  102653.7,
  102788.3,
  102767.7,
  102992.1,
  103114.4,
  103350.9,
  103407,
  103594.1,
  103592.4,
  103607.8,
  103446.4,
  103375.2,
  103162.5,
  102972.8,
  102632.5,
  102576.7,
  102294.1,
  102333.4,
  102288,
  102463.4,
  102512.3,
  102525.2,
  102257.9,
  102044,
  101943.2,
  102058.8,
  101914,
  102018.3,
  101966.2,
  101971.4,
  101919.4,
  102248.6,
  102453.5,
  102506.5,
  102287.2,
  102076.4,
  101886.9,
  102066.9,
  102282.4,
  102632.1,
  102716.1,
  102779,
  102529.3,
  102329.1,
  101960.1,
  101769.6,
  101453,
  101663.1,
  102026.1,
  102418.2,
  102541,
  102798.8,
  102809.7,
  102904,
  102681.4,
  102502.8,
  102327.7,
  102058.7,
  101479.4,
  101014.5,
  100957.9,
  101556.9,
  101991.5,
  102080.6,
  102311.8,
  102490.3,
  102344.2,
  102366.7,
  102241.9,
  102175,
  101935.1,
  101974.1,
  102191.5,
  102512.5,
  102594.9,
  102723.7,
  102741,
  102858.8,
  102743.9,
  102752,
  102689.6,
  102756.2,
  102537.2,
  102360.5,
  102179.5,
  102214.2,
  102161.8,
  102251.4,
  102296.3,
  102410.5,
  102352.6,
  102461.5,
  102640.6,
  103106.7,
  103338.3,
  103481.1,
  103434,
  103480.3,
  103237.3,
  103116.6,
  102955,
  102933.6,
  102733,
  102720.3,
  102735.5,
  102881.1,
  102679.6,
  102646.6,
  102671.1,
  102682.8,
  102366.1,
  102318.4,
  102301.6,
  102325.8,
  102170.8,
  102127,
  101997.5,
  102000.3,
  101708,
  101667.3,
  101646.3,
  101814.7,
  101607.6,
  101602.6,
  101674.4,
  101959,
  101809.1,
  101645.2,
  101579,
  101677.9,
  101558.8,
  101595.2,
  101437.1,
  101718.8,
  101867,
  102112.1,
  102118.5,
  102390.6,
  102368.3,
  102394.1,
  102391.8,
  102366.1,
  102091.8,
  102053,
  101935.2,
  102139.1,
  102082,
  101718.5,
  101876,
  102184.7,
  102005.3,
  102253.7,
  102259.3,
  102255.3,
  102214.9,
  102100.5,
  102021,
  102187.9,
  102192.2,
  102318.8,
  102175.7,
  102189,
  102475.7,
  102539.6,
  102538.2,
  102701.1,
  102527.3,
  102364.9,
  102149.8,
  102059.2,
  101828.5,
  101931.4,
  101989.6,
  102062.9,
  102009.2,
  102293.3,
  102279.3,
  102525.4,
  102650.2,
  102759,
  102652.1,
  102641.5,
  102273.9,
  102047.1,
  101820.6,
  101644.1,
  101769.5,
  102186,
  102305.6,
  102422.1,
  102310.6,
  102234.1,
  102190.6,
  102236.1,
  102076.8,
  102189.6,
  102424.6,
  102753.6,
  102767.3,
  102694.1,
  102552.4,
  102497.5,
  102166.7,
  101984,
  101792.4,
  101658.5,
  101278.9,
  101125.1,
  101002.2,
  100967.7,
  100739.9,
  100852.9,
  101341,
  101783.4,
  101792.1,
  101990.7,
  101990,
  102092.9,
  102158.4,
  102332.3,
  102271.5,
  102301.2,
  102135.7,
  101962.9,
  101820.7,
  101852.9,
  101632,
  101564.4,
  101561.8,
  101734.5,
  101682.9,
  102007,
  102210.6,
  102371.3,
  102245.1,
  102163,
  101901.1,
  101758.6,
  101279.5,
  101180.5,
  101114.8,
  101167.6,
  101018,
  101141.4,
  101445.4,
  101779.7,
  101821.9,
  101906.6,
  101985.2,
  102127.3,
  101960.4,
  101854.6,
  101784.2,
  101828.8,
  101482.1,
  101271.7,
  101149.1,
  101346.1,
  101209.3,
  101309.7,
  101531.7,
  101689.5,
  101553.6,
  101432.4,
  101107.6,
  100794.2,
  100238.6,
  100374.1,
  100795.6,
  101443.4,
  101717,
  102003.6,
  102269.3,
  102674.6,
  102649.4,
  102665.8,
  102495.2,
  102248.2,
  101489.1,
  100877.6,
  100599,
  100873.8,
  101179.1,
  101623.2,
  101721.5,
  102078.5,
  101940.2,
  101728.3,
  101490.4,
  101290,
  100898.7,
  101075.4,
  101386.8,
  101510.8,
  101302.1,
  101321.2,
  101389.5,
  101670,
  101980.3,
  102549.3,
  102700.6,
  102911.4,
  102873.8,
  102752.6,
  102708.2,
  102703.9,
  102472.9,
  102342,
  102237.2,
  102212.7,
  101913.8,
  101867.2,
  101671.2,
  101749.8,
  101523.2,
  101379.6,
  101243.2,
  101114.2,
  100754.4,
  100801.5,
  100955.3,
  101154.5,
  101245.3,
  101375.9,
  101598.4,
  101827.3,
  101874.2,
  101917.6,
  102017.2,
  102204.5,
  102043.9,
  101996.8,
  101866.5,
  101915.1,
  101641.1,
  101426.6,
  101284.6,
  101161.9,
  101000.5,
  101410.8,
  101476.6,
  102005,
  102310.7,
  102380.1,
  102504,
  102646.4,
  102495.8,
  102344.8,
  102206,
  102268.4,
  102074.6,
  101904,
  101959.7,
  102120.8,
  102197,
  102275,
  102341.9,
  102447.7,
  102324.9,
  102174.4,
  102120.4,
  102085.5,
  101742.9,
  101605.3,
  101606.4,
  101576.6,
  101226.2,
  101204.6,
  101186.8,
  101236,
  101039.8,
  100875.8,
  100987.8,
  101224.8,
  101438,
  101690.5,
  102025.2,
  102257.6,
  102264.3,
  102193.9,
  102159.1,
  102189.9,
  101888.7,
  101625.6,
  101533.4,
  101475.5,
  101081,
  100947.8,
  100973.4,
  100807,
  101065.6,
  101288.3,
  101387.9,
  101498,
  101913.6,
  101658.6,
  101690.1,
  101745.9,
  101687.6,
  101623,
  101675.5,
  101856.3,
  101843.2,
  101776.5,
  101813.9,
  101911,
  101788.7,
  101698.9,
  101583.7,
  101643.9,
  101357.6,
  101209,
  101141.6,
  101039.1,
  100726.7,
  100672.7,
  100524.5,
  100590.3,
  100137.5,
  100066.4,
  99852.38,
  100105.5,
  100118.6,
  100556.1,
  100918.1,
  101308.3,
  101127.6,
  101795,
  101815.5,
  102154.8,
  102054.5,
  101955,
  101987.3,
  101953.3,
  101883.1,
  101847.9,
  101779.7,
  101811.1,
  101642.4,
  101477,
  101482.6,
  101613.5,
  101361.6,
  101138.1,
  101117.7,
  100963.9,
  100963.1,
  101101,
  101217.8,
  101371.7,
  101251,
  101314.5,
  101259.1,
  101324.6,
  101531.7,
  101864.1,
  102165,
  102475.6,
  102691.7,
  102626.5,
  102573.8,
  102587.8,
  102413.9,
  102247,
  102129.7,
  102268.8,
  102084.3,
  101857.1,
  101826.9,
  101873.2,
  101722.8,
  101652.9,
  101559.5,
  101685.4,
  101655.2,
  101578.6,
  101548.8,
  101702.1,
  101477.4,
  101508.5,
  101497.8,
  101504.8,
  101271.4,
  101237.1,
  101261,
  101516,
  101674.6,
  101762.1,
  101750.3,
  101781,
  101755.2,
  101618,
  101591.6,
  101540.1,
  101492.1,
  101369.3,
  101393.5,
  101428.7,
  101173.4,
  101189.3,
  101254.5,
  101441.7,
  101367,
  101465.3,
  101513.1,
  101805.8,
  101929.2,
  102013.7,
  102052.7,
  102199,
  102159,
  102036.5,
  102058.1,
  102144.6,
  102267.3,
  102153.2,
  102163.5,
  102290.6,
  102249.1,
  102081.2,
  101997.5,
  101962.3,
  101686.1,
  101388.4,
  101319.5,
  101273.8,
  101042.8,
  101090.1,
  101143.5,
  101430.7,
  101511.8,
  101695.2,
  101652.4,
  101765.3,
  101684.2,
  101429.6,
  101383,
  101368.4,
  101103.4,
  100988.5,
  101086.5,
  101208.8,
  101377.7,
  101822.6,
  101991,
  102162.1,
  102228.6,
  102265.6,
  102227.5,
  102286.5,
  102233.7,
  102042.6,
  101886.5,
  101936.8,
  101649.2,
  101239.1,
  101193.8,
  101062.1,
  100593.8,
  100356,
  100322.9,
  100643.1,
  100882.6,
  101189.7,
  101045.1,
  100988.5,
  100828.5,
  100801.4,
  100823.6,
  101015.4,
  101113.4,
  101132.4,
  101007,
  101099.3,
  100899.7,
  100718.4,
  100600.5,
  100406.3,
  99906.87,
  100345.2,
  100976.5,
  101383.4,
  101477,
  101425.2,
  101283.2,
  101205.1,
  101011.7,
  101020,
  100928.7,
  101014.2,
  100905.5,
  101126.7,
  100875.7,
  100966.7,
  100936.1,
  101370.8,
  101738.2,
  102028.2,
  102079,
  102013.4,
  102291.2,
  102242,
  102054.1,
  101845.9,
  101653.4,
  101688.1,
  101485.6,
  101424.8,
  101529.5,
  101770,
  101985.6,
  102136.5,
  102178.7,
  102340.5,
  102279.5,
  102107.2,
  102011.4,
  102022.1,
  101825,
  101717,
  101725.5,
  101887.4,
  101717.4,
  101551.8,
  101595.7,
  101590.8,
  101227.2,
  101064.3,
  101134.3,
  101168.5,
  100909.1,
  101011.6,
  101026.8,
  101165,
  101002,
  101096,
  101163.5,
  101252.7,
  101059.5,
  101162.7,
  101127.8,
  101187.6,
  100933.4,
  101055.7,
  100992.8,
  101189.1,
  101016.1,
  101011.2,
  101109,
  101197.9,
  101040.9,
  100993.4,
  101027.3,
  101112.9,
  100875.1,
  100886.6,
  100896.3,
  100986,
  100704.8,
  100590.7,
  100548.6,
  100552.5,
  100426.8,
  100635.2,
  100780.8,
  101004.4,
  101054.3,
  101194.5,
  101207.5,
  101345.7,
  101195.9,
  101166.3,
  101268,
  101357,
  101136.7,
  101090.8,
  101141.7,
  101209.2,
  101049.3,
  101008,
  101064.5,
  101039.6,
  100681.1,
  100668,
  100794.8,
  101015.3,
  101092.4,
  101225.6,
  101409.1,
  101576,
  101432.7,
  101248.9,
  101262.1,
  101227,
  100936.3,
  100816.6,
  100879.6,
  100935.8,
  100745.5,
  100729.5,
  100667.6,
  100490.6,
  99902.05,
  100170.3,
  100707,
  101000.2,
  101224.8,
  101300.7,
  101087.1,
  101126.2,
  101001.9,
  100767.8,
  100715.4,
  100558.1,
  100087.9,
  100018.1,
  100256.1,
  100619.5,
  100655.2,
  100835.8,
  100821.9,
  101090.4,
  101191.6,
  101723.1,
  102009.8,
  102296.2,
  102182.1,
  102147.5,
  102019.6,
  102041.4,
  101617.8,
  101513.7,
  101426.2,
  101435.1,
  101152.9,
  101084.9,
  101092.2,
  101119.5,
  100920.7,
  100965.2,
  100910.6,
  101118.6,
  101056.7,
  101195.7,
  101251,
  101388.3,
  101405.2,
  101457,
  101524.7,
  101699,
  101640.5,
  101624.4,
  101679.4,
  101859.4,
  101529.2,
  101383.4,
  101296.8,
  101353.8,
  101045,
  100940.9,
  101057.3,
  101208.3,
  100967.3,
  100904.1,
  101045.2,
  101115.6,
  100816.9,
  100726.1,
  100839,
  100869.5,
  100711.2,
  100879.8,
  100995.8,
  101219,
  101030.5,
  101143.5,
  100921.2,
  100894.3,
  100438,
  100386.8,
  100387.1,
  100832.5,
  101146.7,
  101316.7,
  101420.3,
  101570.2,
  101595.5,
  101578.7,
  101577,
  101649,
  101537.7,
  101431.2,
  101419.1,
  101437.4,
  101455.5,
  101390.8,
  101548.2,
  101691.7,
  101630.2,
  101554.6,
  101704.4,
  101817,
  101610.3,
  101546.8,
  101586.4,
  101647.5,
  101365,
  101221.3,
  101198.5,
  101184.2,
  100868.9,
  100779.1,
  100635.9,
  100580.6,
  100388.2,
  100388.9,
  100434.9,
  100798.4,
  100899.1,
  101148.8,
  101192.2,
  101284.6,
  101216.7,
  101214.6,
  101214.9,
  101316.2,
  101227.8,
  101279.9,
  101387.8,
  101520.7,
  101429.4,
  101530.1,
  101623.9,
  101845.6,
  101732.4,
  101709.5,
  101754.3,
  101928.8,
  101758.5,
  101757.4,
  101750.1,
  101877.1,
  101724.3,
  101764.6,
  101807.7,
  101931.3,
  101747.2,
  101643.2,
  101669.5,
  101667.9,
  101352.9,
  101186.2,
  101209,
  101146,
  100762.7,
  100737.5,
  100780.7,
  100983.2,
  100957.7,
  101103.4,
  101199.7,
  101392.9,
  101195.1,
  101158.1,
  100966.7,
  100978.5,
  100553.9,
  100623.3,
  100532.1,
  100866.1,
  100770.3,
  101025.9,
  101047.9,
  101202.4,
  100957.8,
  101161.2,
  100961.1,
  101064.6,
  101091.6,
  101283.8,
  101498.4,
  101596.9,
  101554.2,
  101500.7,
  101555.2,
  101633.3,
  101266.2,
  101143.2,
  101134.6,
  101186,
  100921.9,
  101019.6,
  101099.8,
  101430.6,
  101686.9,
  101937.3,
  101959.6,
  102165.1,
  101940.1,
  101807.1,
  101802.2,
  101671.2,
  101141.3,
  101097,
  101122.9,
  101276.5,
  101133,
  101454.6,
  101531.2,
  101867.6,
  102042.8,
  101955.1,
  101877.2,
  101868.2,
  101499.6,
  101085.9,
  100976.4,
  100927.1,
  100540.8,
  100431.9,
  99834.67,
  99955.52,
  100184.1,
  100835.7,
  101436.7,
  101927.1,
  102083.7,
  102260.1,
  102281.1,
  102448.1,
  102335.1,
  102181.7,
  102131.6,
  102112.8,
  101898.4,
  101788.4,
  101713.6,
  101801.2,
  101669.2,
  101634.7,
  101622.1,
  101784.8,
  101704.3,
  101745.7,
  101741.4,
  101929.1,
  101857.3,
  101880.5,
  101902.1,
  102044.8,
  101943.4,
  101933.6,
  101926.8,
  102054,
  102076.6,
  102039.5,
  102127.6,
  102264.7,
  102235.1,
  102143.3,
  102081.7,
  102216,
  102125.6,
  102029.5,
  101985.4,
  102126.5,
  102020.8,
  101937.7,
  101861.6,
  101998.6,
  101695.1,
  101454.3,
  101358.3,
  101302.9,
  100767.8,
  100484.3,
  100532.8,
  100591.8,
  100624.7,
  100870,
  100940.8,
  100969.9,
  100664.5,
  100551.6,
  100451.9,
  100465.7,
  100912.8,
  101030,
  101259.9,
  101629.4,
  101776.2,
  101905.4,
  102122.4,
  102315.8,
  102254.4,
  102085,
  101998.1,
  101960.8,
  101596.4,
  101455.9,
  101439,
  101542.7,
  101497.9,
  101840,
  102087.1,
  102285.6,
  102145,
  102506.1,
  102252.6,
  102267.6,
  102101.6,
  102054.5,
  101951.4,
  101896,
  101680.1,
  101724.7,
  101623.4,
  101642.3,
  101511.9,
  101544.3,
  101485.2,
  101538.1,
  101434.9,
  101419,
  101377.9,
  101466.2,
  101384.2,
  101517.4,
  101842.7,
  102264,
  102406.1,
  102572.9,
  102687.6,
  102798.7,
  102686.2,
  102669.3,
  102573,
  102682.8,
  102440,
  102351.8,
  102411.3,
  102401.8,
  102259.4,
  102233.5,
  102070.6,
  102001.2,
  101803.6,
  101569.8,
  101484.3,
  101504.8,
  101477.3,
  102157.4,
  102582.3,
  102773.3,
  102806.7,
  102782.7,
  102622,
  102564.2,
  102227.7,
  101962.2,
  101754.7,
  101689.9,
  101370,
  101227.1,
  101380,
  101601.4,
  101507.3,
  101550.8,
  101562.9,
  101747,
  101566.4,
  101527.3,
  101540,
  101604.4,
  101445.2,
  101433.7,
  101393.6,
  101337.2,
  101187.6,
  101193.6,
  101194.2,
  101193.4,
  100960.9,
  100983.3,
  100998.8,
  101058.1,
  100727.7,
  100861.3,
  100886.2,
  100819.4,
  100684.6,
  101516.3,
  101751.3,
  102208.1,
  102182,
  102267.6,
  102367.3,
  102329.6,
  102322.5,
  102384.7,
  102443.6,
  102502.6,
  102473.9,
  102528.6,
  102388.9,
  102196,
  101828,
  101650.3,
  101252.2,
  101145,
  101110.8,
  101285.4,
  101230.2,
  101187,
  100836.1,
  100718.7,
  100671.9,
  100594.5,
  100773.2,
  101096.3,
  101013.3,
  101001.6,
  100838.5,
  101109.5,
  101149.2,
  101747,
  102206,
  102622.2,
  102885.4,
  103145.5,
  103125.1,
  103170,
  103151.4,
  103193.5,
  103007.6,
  102858,
  102606.9,
  102378.6,
  102078.9,
  101879.5,
  101572.8,
  101537,
  101288.5,
  101192.1,
  101287.4,
  101662,
  101749.8,
  101870.8,
  101817.4,
  101401,
  100711.6,
  100729.8,
  101647.5,
  102060.8,
  102215.4,
  102370.3,
  102414.1,
  102546.2,
  102515.7,
  102617.1,
  102525.9,
  102504.2,
  102249.5,
  102063.4,
  101791.3,
  101618.3,
  101319.7,
  101380.5,
  101635.4,
  102073.2,
  102323.9,
  102548.3,
  102569.4,
  102725.5,
  102695.4,
  102780.5,
  102800,
  102854.9,
  102706.7,
  102588.7,
  102402.2,
  102276.3,
  101985.8,
  101943.2,
  101847,
  101972.9,
  101754.5,
  101797.5,
  101775.8,
  101863.3,
  101840,
  101830.4,
  101846.7,
  101775.6,
  101538.2,
  101422.8,
  101326.1,
  101252.4,
  100731,
  100946.8,
  101208.6,
  101575.6,
  101755.5,
  101819.9,
  101863.6,
  101743.8,
  101307.9,
  101306,
  101183.2,
  101168.1,
  100559.1,
  100580.1,
  100906.4,
  101214.2,
  101382.3,
  101651.9,
  101688.8,
  101695.1,
  101462,
  101463.5,
  101322.5,
  101190.5,
  100991.6,
  101216.2,
  101323.1,
  101425.4,
  101372,
  101180.1,
  100987.7,
  100187.6,
  99324.68,
  99189.9,
  99779.72,
  100134.4,
  100450.4,
  100986.5,
  101412.2,
  101751.3,
  101967.1,
  102217.1,
  102411.4,
  102434.4,
  102219,
  102238.9,
  102320.8,
  102534,
  102559,
  102589.1,
  102515.4,
  102380,
  102281.3,
  102356.2,
  102458.7,
  102544.9,
  102509.6,
  102572.3,
  102558.3,
  102542.2,
  102358.6,
  102295.1,
  102207.2,
  102143.1,
  101853.6,
  101804.5,
  101712.3,
  101653.2,
  101715.8,
  102026.1,
  102231.1,
  102554.2,
  102697.7,
  102799.4,
  102799.7,
  102701.3,
  102474.3,
  102317.6,
  102178,
  102138,
  101979.9,
  101974.6,
  102061.7,
  102132.7,
  102099.2,
  102188.7,
  102252.9,
  102365.2,
  102236.9,
  102200.3,
  102073,
  102115.8,
  101869.5,
  101933,
  101981.9,
  102059,
  101974,
  101922.2,
  101673.4,
  101620.2,
  101758.9,
  102328.9,
  102544.4,
  102669.1,
  102427.7,
  102384.9,
  102162.4,
  101908.3,
  101642.4,
  101697.5,
  101834.1,
  101958.5,
  101930.3,
  101923,
  101767.5,
  101666.7,
  101774.7,
  102255.3,
  102509.2,
  102704.1,
  102626.1,
  102645,
  102446.5,
  102400.5,
  102206.9,
  102183.6,
  102073.2,
  102063.6,
  101817.5,
  101755,
  101775.2,
  101831.7,
  101745.6,
  101840.5,
  101783.5,
  101647,
  101334,
  101113.8,
  100533.1,
  100650.8,
  100834.5,
  101016.2,
  101014.5,
  101025.7,
  101366.9,
  101517.5,
  101601.7,
  101748.5,
  101712.6,
  101695.1,
  101596.4,
  101502.5,
  101369.8,
  101588,
  101559.2,
  101432.4,
  101370.2,
  101515.9,
  101522.3,
  101605.5,
  101641,
  101961.7,
  102146,
  102460.6,
  102811.4,
  103071.2,
  103176.6,
  103178.2,
  103098.8,
  102851.2,
  102506.9,
  101992.5,
  101587.5,
  101468.1,
  101461.8,
  101809.6,
  101826,
  101746.4,
  101417.3,
  101029.6,
  100790.4,
  100941.6,
  100814.4,
  100626.9,
  100347.9,
  100446.8,
  100882.7,
  101387.8,
  101789.4,
  102187.1,
  102386.5,
  102606.8,
  102564.4,
  102469.1,
  102352.5,
  102290.8,
  102128.8,
  102328.5,
  102489.9,
  102697.4,
  102766.3,
  102783,
  102715.5,
  102655.2,
  102299.7,
  102061.6,
  101709.9,
  101501.2,
  101254.4,
  101527.3,
  101746.9,
  102086.5,
  102391.9,
  102791.9,
  103034.5,
  103420.1,
  103620.2,
  103834.5,
  103853.8,
  103806.2,
  103677.6,
  103574,
  103447,
  103347,
  103080,
  102897.8,
  102652,
  102669.5,
  102360.1,
  102219.6,
  102163.8,
  102120.4,
  101870.2,
  101564.5,
  101854.6,
  101953.5,
  101907.6,
  101854.2,
  101672.3,
  101428.7,
  101136.4,
  101067.2,
  100895.5,
  101137.2,
  101293.3,
  101274.9,
  100831.8,
  100933.3,
  101058.3,
  101100,
  101228.7,
  101628.7,
  102050.8,
  102323.3,
  102559.2,
  102708.3,
  102818.1,
  103010.1,
  103094.3,
  103177.6,
  103036.5,
  102820.5,
  102547.6,
  102339.4,
  102024.2,
  101902.6,
  101944.5,
  101985.6,
  101999,
  102211.2,
  102280,
  102401.5,
  102337.8,
  102309.2,
  102263.1,
  102292.2,
  102287.7,
  102611.5,
  102599.8,
  102728.2,
  102757,
  102935.4,
  102869.4,
  102955.9,
  102835.7,
  102824.3,
  102750.4,
  102778.9,
  102565.4,
  102519,
  102345.9,
  102275.7,
  102015.5,
  101997,
  102013.1,
  102199.8,
  101852.8,
  101939.6,
  101677.9,
  101785.9,
  101694.9,
  101782.5,
  101660.1,
  101741.2,
  101666.4,
  101565,
  101364.9,
  101234.6,
  101109.4,
  101145.3,
  101199.9,
  101351.6,
  101224.4,
  101402.8,
  101585.2,
  101973.6,
  102095.4,
  102251.1,
  102134.9,
  101810.2,
  101169.4,
  100925.9,
  101221.5,
  101693.3,
  101792.1,
  101858.1,
  101890.5,
  102017.1,
  102012.4,
  102143.6,
  102150.8,
  102215.1,
  102218.6,
  102480.5,
  102711.1,
  103008.4,
  103153.7,
  103443.1,
  103650.7,
  103923.9,
  104000.8,
  104103.1,
  104065.1,
  104104.9,
  104006.1,
  104029.4,
  103942.8,
  104029.4,
  103902.4,
  103830.8,
  103615.4,
  103347.7,
  102975.8,
  102716.7,
  102487.9,
  102413.1,
  102066,
  102023.1,
  102005.8,
  101921.1,
  101452.5,
  101241.8,
  101362.6,
  101662.2,
  101679.8,
  101838.6,
  101933.8,
  102063.2,
  101965,
  101962.4,
  101839.9,
  101719.2,
  101375.9,
  101231.8,
  101004.5,
  100892,
  100554.7,
  100667,
  100772.4,
  101047.7,
  101294.4,
  101385.1,
  101499.2,
  101698.3,
  101417.8,
  101168.6,
  100699.5,
  100872.2,
  100987.7,
  101154.7,
  101363.6,
  101616.2,
  101515.8,
  101846.5,
  102050.8,
  102318.1,
  102456,
  102848.4,
  103055.7,
  103229.9,
  103197.7,
  103353.3,
  103338.1,
  103370.8,
  103231.7,
  103242.7,
  103118.2,
  103089.5,
  102912.5,
  102956,
  102849,
  102956.5,
  102835.9,
  102920.5,
  102948.1,
  103071,
  102931.3,
  102942.9,
  102845.9,
  102966.4,
  102708.4,
  102670,
  102611.9,
  102697.4,
  102377,
  102290.5,
  102166.3,
  102084.5,
  101703.9,
  101637.1,
  101651.1,
  101951.7,
  102039.5,
  102435.6,
  102437.7,
  102514,
  102181.4,
  102102.6,
  102059.9,
  102393.7,
  102647,
  102853.5,
  102708.7,
  102599.5,
  102124.4,
  101854,
  101715.6,
  101864.4,
  101675.3,
  101738.3,
  101868.5,
  102115.3,
  102107.3,
  102132.1,
  102096.6,
  102320.3,
  102083.5,
  101743.1,
  101607.6,
  101869.1,
  101926,
  102191.1,
  102227.8,
  102519.7,
  102429.7,
  102420.4,
  102221.6,
  102348,
  102129.8,
  102129.4,
  102203.2,
  102422.9,
  102317.7,
  102337.1,
  102177.8,
  102219.6,
  102070.6,
  102105.5,
  102088.3,
  102289.5,
  102262.9,
  102200.9,
  102114.3,
  102212.8,
  102091.7,
  102048.1,
  101888.5,
  101847.2,
  101568.3,
  101393.7,
  101172.3,
  101324.9,
  101243.2,
  101481.2,
  101701.7,
  101808.8,
  101665,
  101784.2,
  101575.2,
  101567.1,
  101508.1,
  101248.7,
  101354.8,
  101013,
  100590.3,
  100730.4,
  101040.9,
  101474.2,
  101806.7,
  102044.1,
  102199.2,
  102273.8,
  102371.2,
  102549,
  102928.5,
  103217.2,
  103342.4,
  103421.7,
  103399.9,
  103274.9,
  102853.9,
  102541.3,
  102254.5,
  102067.7,
  101830.8,
  101819.5,
  101996.7,
  102255.8,
  102367.7,
  102386.5,
  102376.8,
  102317.9,
  102280.9,
  102199.4,
  102130.7,
  102109.4,
  101928.9,
  101837.6,
  101670.1,
  101734.5,
  101554.9,
  101676.9,
  101770.5,
  101982,
  101813,
  101578.3,
  101405.2,
  101514.1,
  101749.1,
  102013.7,
  102191.1,
  102365.4,
  102106.9,
  101907.3,
  101788.7,
  101781.5,
  101534.2,
  101747.7,
  101883.5,
  102026.1,
  102141,
  102268.8,
  102256.5,
  102478.5,
  102447.3,
  102439.3,
  102421.6,
  102589.3,
  102410.6,
  102254.3,
  102193.5,
  102279.5,
  101908.8,
  101826.9,
  101873.1,
  101898.7,
  101733.4,
  101877.4,
  101895.6,
  102076.2,
  102142,
  102107.5,
  102158,
  102273.1,
  102197.2,
  102158.2,
  102061.5,
  102221,
  102083.2,
  101906.5,
  101859.4,
  101992.2,
  101742.3,
  101987.3,
  101962.4,
  102195.9,
  102394.4,
  102558.1,
  102639.3,
  102721.8,
  102530.2,
  102326.8,
  101980.5,
  101738.5,
  101156.4,
  100697.2,
  100461.6,
  100462.7,
  100534.3,
  101206.8,
  101798.4,
  102195.8,
  102265.9,
  102283,
  102280.5,
  102377.4,
  102143.5,
  101929.3,
  101897.7,
  101845,
  101517.4,
  101277.4,
  101137.5,
  101235.4,
  101082.8,
  101085,
  101161.4,
  100841.4,
  100809,
  100273.6,
  100464.4,
  100673.8,
  100606,
  101003.9,
  101158.2,
  101548.2,
  101623.3,
  101772.7,
  101703.3,
  101731.5,
  101464.1,
  101223.5,
  101136.1,
  101264.6,
  101191.9,
  101550.3,
  101791,
  102054.3,
  102057.2,
  102002.5,
  102172.6,
  102265.8,
  102303.5,
  102297.1,
  102440.7,
  102564.1,
  102508.7,
  102344,
  102247.9,
  102353.5,
  102187,
  101991,
  101937.6,
  101896.3,
  101592.4,
  101316.8,
  101359.3,
  101369.9,
  101107.9,
  100964.3,
  100908.6,
  100931.7,
  100659.2,
  100564.6,
  100524.4,
  100707.5,
  100630.3,
  100631.5,
  100661.4,
  100723.3,
  100750.2,
  100418.1,
  100642.7,
  100827.6,
  100887.2,
  101118.2,
  101714.1,
  102160.2,
  102403,
  102473.7,
  102481.6,
  102488.1,
  102211.1,
  102026.1,
  101915.5,
  101866.8,
  101436.6,
  101225.9,
  101004.4,
  100688.6,
  99926.23,
  99654.42,
  100258.2,
  100708.4,
  100711.7,
  101029,
  101256.9,
  101669.9,
  102061.4,
  102049.1,
  102083.2,
  102317.9,
  102022.6,
  101829.4,
  101627.5,
  101605.4,
  101196.9,
  101142.1,
  100943.1,
  101182.8,
  101462.3,
  101680.2,
  101850.6,
  102073.6,
  102074.1,
  102057.8,
  102112.7,
  102228,
  101997.5,
  101826.1,
  101807.4,
  101753.7,
  101446,
  101274.7,
  101184.4,
  101053.2,
  100783.7,
  100709,
  100887.4,
  101126.2,
  101120.2,
  101180.2,
  101340.2,
  101576.3,
  101431.3,
  101501.7,
  101547.8,
  101695,
  101567.2,
  101581.5,
  101588.9,
  101701.3,
  101365.4,
  101482.9,
  101392.5,
  101241.8,
  100971,
  100957.2,
  100817.2,
  100865.1,
  100851.9,
  101118.3,
  101389.9,
  101572.1,
  101644.6,
  101627.4,
  101594.8,
  101690.5,
  101457.7,
  101280.5,
  101364.3,
  101475.8,
  101271.9,
  101008.1,
  100980.8,
  101012.9,
  100722.1,
  100548.8,
  100849.9,
  100705,
  100437,
  100736.3,
  101043.8,
  101435.1,
  101526.7,
  101634.4,
  101766.4,
  101926.8,
  101887.4,
  101897.4,
  101948.1,
  101883.7,
  101705.4,
  101624.5,
  101682,
  101795.8,
  101704.3,
  101591.9,
  101686.2,
  101820.6,
  101540,
  101347,
  101290.4,
  101307.5,
  101243.6,
  101648.3,
  101876.6,
  102126.3,
  102210.9,
  102226.1,
  102185.5,
  102279.9,
  102213.6,
  102081.3,
  102094.9,
  102297.5,
  102089.4,
  101951.6,
  101932.4,
  102041.8,
  101798.9,
  101633.2,
  101661.3,
  101766.2,
  101474.5,
  101355.8,
  101590.7,
  101715.2,
  101483.4,
  101424.6,
  101418.9,
  101537.9,
  101179.5,
  100850.1,
  100586,
  100628.7,
  100508.2,
  100632.2,
  100905.9,
  101246.3,
  101510.9,
  101743.3,
  101939.4,
  102211.4,
  102271.4,
  102245.1,
  102273.3,
  102351.3,
  102018.9,
  101764,
  101649.6,
  101598.2,
  101132,
  100911.5,
  100950.7,
  101008.7,
  100772.3,
  100622.6,
  100682.6,
  100873.5,
  100697.9,
  100616,
  100607.6,
  100849.5,
  100599.9,
  100522.4,
  100684.7,
  101094.9,
  101193.2,
  101243.9,
  101303.8,
  101413.4,
  101326.9,
  101199.9,
  100973.1,
  100839.2,
  100369.4,
  100316.6,
  100598,
  101143.7,
  101430.4,
  101665.9,
  101862.6,
  101963.3,
  101842.2,
  101727,
  101836.7,
  101909.9,
  101668.8,
  101522.4,
  101589.5,
  101601.3,
  101170.9,
  101062.4,
  101186.7,
  101220.5,
  101028.2,
  100652.7,
  100664.5,
  100912.6,
  101108.6,
  101317.5,
  101467.5,
  101733.2,
  101772.3,
  101478,
  101494.7,
  101598.7,
  101284.8,
  101084.7,
  101216.2,
  101462.1,
  101479.2,
  101395.7,
  101245.7,
  101162.3,
  100658.2,
  100427.4,
  100494.6,
  100574.2,
  100538.7,
  100675.8,
  100792.6,
  100882.5,
  100914.2,
  100843.5,
  100816.2,
  100883,
  100417.9,
  100674.1,
  100582.6,
  100797,
  100703.8,
  100792.1,
  100881.8,
  101122.2,
  101216.4,
  101436.7,
  101459,
  101755,
  101680.2,
  101734.7,
  101850.1,
  102000.4,
  101710.2,
  101572.9,
  101618.6,
  101630.9,
  101301.2,
  101079.4,
  101130.2,
  101171.1,
  100838.2,
  100737.1,
  100826.1,
  100936.1,
  100704.1,
  100765.8,
  100893.4,
  101028.5,
  100760.1,
  100829.8,
  101011.2,
  101186.1,
  100921.4,
  100821,
  100846.4,
  100904.3,
  100665.6,
  100553,
  100611.2,
  100776,
  100579.8,
  100529.2,
  100644.6,
  100874.4,
  100780.1,
  100830.3,
  100962.7,
  101023.3,
  100658.8,
  100747.3,
  100802.1,
  101051.4,
  101308.6,
  101362.5,
  101252.1,
  100971.3,
  100468.2,
  100035.4,
  99941.38,
  100354.5,
  100684.5,
  101267.8,
  101611.5,
  101970.4,
  102089,
  102086.9,
  102007.1,
  102093.3,
  101796.8,
  101505.6,
  101327.3,
  101252.6,
  100868.3,
  100726.9,
  100633.4,
  100761.9,
  100587.5,
  100756.9,
  100938.9,
  101224.7,
  101225.3,
  101196.2,
  101056.1,
  101108.6,
  100792.6,
  100569.5,
  100668,
  100847,
  100990.1,
  101124.7,
  101398,
  101691.3,
  101588.7,
  101562.8,
  101445.2,
  101377.9,
  101090.3,
  100911.3,
  100822.8,
  100867.6,
  100531,
  100539.5,
  100448.3,
  100687,
  100524.7,
  100511.9,
  100536,
  100946.2,
  100809,
  101097.8,
  100982.8,
  101238.3,
  101222.2,
  101398.1,
  101435.4,
  101654.6,
  101578.5,
  101584.1,
  101652.5,
  101730.1,
  101595,
  101404.7,
  101465.4,
  101523.9,
  101403.1,
  101357.9,
  101428,
  101613.1,
  101472.2,
  101394.9,
  101366.1,
  101520.8,
  101304.1,
  101217.8,
  101190.4,
  101277.3,
  101180.1,
  101091.3,
  101095.7,
  101216.9,
  101174.4,
  101233.4,
  101220.1,
  101270.7,
  100987.5,
  100821.1,
  100774.9,
  100918,
  100989.8,
  101134.1,
  101229.9,
  101644.9,
  101834.9,
  101985.9,
  102025.4,
  102181.3,
  102000.2,
  101797.2,
  101704.6,
  101733.8,
  101418.3,
  101219.4,
  101164.8,
  101094.4,
  100637.5,
  100540,
  100444.4,
  100247.9,
  99708.23,
  99539.55,
  99365.99,
  99928.23,
  100179.8,
  100590.5,
  100905.9,
  101148.5,
  101240.2,
  101333,
  101398,
  101537.9,
  101329.1,
  101200.4,
  101327.9,
  101646.1,
  101396.2,
  101264.6,
  101285.7,
  101504.5,
  101401.9,
  101394.2,
  101455.1,
  101502.8,
  101300.3,
  101132,
  101090.9,
  101099.9,
  100676.5,
  100584.8,
  100719.2,
  100877.1,
  101010.5,
  101096.9,
  101044.8,
  101037,
  101081.3,
  101347.9,
  101524.5,
  101857,
  102036.3,
  102157.9,
  102342.6,
  102479.8,
  102456.4,
  102461,
  102414.6,
  102431.7,
  102243.8,
  101976.5,
  101781.4,
  101844.3,
  101526.1,
  101260,
  101311,
  101339,
  101039.3,
  100935.7,
  101029.8,
  101067.9,
  100732.1,
  100709.9,
  100741.9,
  100724.6,
  100252.3,
  100306.9,
  100640.2,
  100962.7,
  100167,
  100887.9,
  100877.8,
  101319.8,
  101403.6,
  101544.7,
  101541.2,
  101607.2,
  101295.3,
  101175.2,
  100681.3,
  100640.1,
  100671,
  101066.7,
  101185.6,
  101374.6,
  101201.9,
  101179.3,
  101169.7,
  101276.6,
  101100,
  101144.4,
  101357.2,
  101691.7,
  101961.8,
  102214.1,
  102485.5,
  102751,
  102728.1,
  102609.7,
  102509.2,
  102558.5,
  102189.1,
  101854.8,
  101732.2,
  101608.6,
  101185.5,
  100978.8,
  100941.7,
  101498,
  101951.6,
  102294.2,
  102443.1,
  102629.3,
  102646,
  102490.8,
  102476.9,
  102541.9,
  102342.6,
  102201.8,
  102198.5,
  102298.6,
  102151,
  102147,
  102205.2,
  102372.9,
  102351.6,
  102345.8,
  102317.4,
  102366.9,
  102213.7,
  102113.5,
  102063.3,
  102029.1,
  101768.1,
  101615.1,
  101489.2,
  101596.7,
  101352.9,
  101446.3,
  101477.8,
  101579,
  101303,
  101225,
  101014.7,
  100666.1,
  100372.1,
  100123,
  99892.8,
  100108.6,
  100254.3,
  100559.8,
  100720,
  101010.9,
  101232.3,
  101549.8,
  101754.3,
  101944.6,
  101792.5,
  101700.7,
  101743.2,
  101927.1,
  101852.3,
  101994.8,
  102065.3,
  102178.5,
  102015,
  101882.1,
  101830,
  102047.2,
  101970.2,
  102055.5,
  102084.7,
  102346.1,
  102266.9,
  102216.1,
  102178.8,
  102315.7,
  102076.3,
  101920.6,
  101866.1,
  101926.4,
  101632.3,
  101465.3,
  101375.4,
  101464.4,
  101158.9,
  101068.4,
  100877.4,
  100856.9,
  100572.5,
  100619.2,
  100893,
  101054.8,
  101239,
  101594.3,
  101640.3,
  101837.4,
  101868.9,
  101878.4,
  101911.9,
  102014.6,
  101860.9,
  101818.4,
  101837.2,
  101991.1,
  101732.9,
  101706.2,
  101805.2,
  101867.6,
  101648.6,
  101743.1,
  101722.2,
  101691.9,
  101473.8,
  101310.1,
  101007.6,
  100775,
  100292.8,
  100491.1,
  100957,
  101251.6,
  101385.1,
  101390.2,
  101728.1,
  101852.7,
  101933.3,
  102144,
  102190.2,
  102245.5,
  101997.6,
  101734.9,
  101426.7,
  101364.3,
  100952.4,
  101126.5,
  101416.7,
  101731.6,
  101910.8,
  102189.3,
  102420.7,
  102511.1,
  102331.6,
  102148.8,
  101984.2,
  101942.5,
  101737.6,
  101570.8,
  101426.9,
  101484.7,
  101458.1,
  101724.3,
  101913,
  102126.9,
  102135.4,
  102166.9,
  102098.2,
  102044.8,
  101774.1,
  101560.6,
  101543.2,
  101561.8,
  101392.9,
  101375.1,
  101402.3,
  101427.1,
  101229.7,
  101208.1,
  101032.3,
  101006,
  101062.5,
  101137.8,
  100576.7,
  101159.4,
  101211,
  101412.1,
  101257.2,
  101580.2,
  101679.9,
  101848.4,
  102050.7,
  102107.7,
  102140.5,
  102070.5,
  101874.1,
  101778.8,
  101583.3,
  101556,
  101537.9,
  101601,
  101413,
  101421,
  101398.1,
  101394,
  101130.9,
  101211.5,
  101334.5,
  101453.3,
  101363.6,
  101363.9,
  101376.9,
  101622.6,
  101752.4,
  101878.8,
  101992.3,
  102128.1,
  102101.1,
  102064.4,
  101975.7,
  101919,
  101708.3,
  101658.7,
  101595.7,
  101496.4,
  101180.5,
  101118.6,
  100999.1,
  100718.9,
  100333.1,
  100536,
  100570.8,
  100667.9,
  100764,
  101320.6,
  101489.7,
  101657.8,
  101957.7,
  102452.9,
  102650.5,
  102785.2,
  102783.3,
  102766.4,
  102748.5,
  102775.8,
  102552.6,
  102565.4,
  102419.3,
  102277.4,
  101904.6,
  101869.9,
  101727.1,
  101729.6,
  101640.3,
  101693.7,
  101577.1,
  101412,
  100235,
  100296.6,
  100945.3,
  101379.2,
  101718.9,
  102204.9,
  102414,
  102594.5,
  102603.9,
  102375.4,
  102031.1,
  101674.3,
  101090.4,
  100920.2,
  101098.9,
  101692.8,
  102036,
  102248.9,
  102207.5,
  102133.9,
  101733.1,
  101566.7,
  101484,
  101494.6,
  101289.6,
  101346.8,
  101404.1,
  101551.7,
  101463.3,
  101502.7,
  101445.9,
  101553.1,
  101396.4,
  101452.3,
  101297.6,
  101178.4,
  100468.8,
  100637.2,
  100765.9,
  101083.7,
  101153.6,
  101349,
  101477.2,
  101812,
  102078.2,
  102308.5,
  102267.4,
  102145.2,
  101269.8,
  100599.5,
  100140.1,
  100844,
  101113.1,
  101521,
  101655.8,
  101773.1,
  101792.1,
  101863,
  101851.4,
  101992,
  102097.7,
  102415.1,
  102573.2,
  102684.8,
  102453.2,
  102493.2,
  102393.1,
  102409.9,
  102293.8,
  102305.9,
  102328.1,
  102508.7,
  102472.3,
  102422.4,
  102264.1,
  102196.3,
  101930.3,
  101790.2,
  101771.8,
  101817.7,
  101756.4,
  101942.7,
  102028.5,
  102120.2,
  102039.4,
  102157.9,
  101999.3,
  101971.2,
  101651.5,
  101562.1,
  101660.8,
  101677.6,
  101571.7,
  101607.8,
  101379.4,
  101183,
  100939.9,
  101348.5,
  101655.2,
  101945.4,
  102217.4,
  102621.8,
  102703.3,
  102813.8,
  102742.9,
  102755.7,
  102631.9,
  102534.9,
  102186.8,
  102168.6,
  102061.1,
  101974.4,
  101701.4,
  101674.5,
  101542.5,
  101688.9,
  101550.1,
  101901.1,
  102278.8,
  102409.4,
  102639.7,
  102564.7,
  102528.7,
  102411.1,
  102200.1,
  102098.8,
  101976.5,
  102107.3,
  101978.3,
  101979.3,
  101842.3,
  101810.9,
  101475.6,
  101449,
  101435.2,
  101449.8,
  101329,
  101477,
  101548.2,
  101545.3,
  101297,
  101300.6,
  101127.7,
  100898.8,
  100601.8,
  100400,
  100348,
  100693,
  100757,
  101006.4,
  101117.9,
  101205.4,
  101111.4,
  101245.6,
  101293.6,
  101535.1,
  101697.5,
  102057,
  102241.4,
  102297,
  102310.1,
  102419.5,
  102457.9,
  102424.3,
  102198.4,
  102321.7,
  102231.9,
  102210.6,
  102215.2,
  102429.6,
  102320.5,
  102304.1,
  102182.1,
  102037.8,
  101882.1,
  101790.5,
  101667.9,
  101717,
  101714.6,
  101811,
  101853.6,
  102023.8,
  101904,
  101910.3,
  101938.9,
  102261.2,
  102625.1,
  102815.8,
  102942.5,
  102893,
  102543.7,
  102249.1,
  101623.2,
  101327.2,
  100986.1,
  100805.2,
  100640.8,
  101125,
  101397.6,
  101524.9,
  101376.3,
  101330.5,
  101378.2,
  101520.7,
  101501.2,
  101678.5,
  101760.3,
  101950.4,
  102122.1,
  102451.6,
  102654,
  102800.1,
  102928.3,
  103070.7,
  103112.2,
  103148.1,
  103109.1,
  103073.1,
  102982,
  102886.7,
  102497.8,
  102292.9,
  102216,
  102201.8,
  102065.6,
  102239.8,
  102260.6,
  102346.2,
  102243.9,
  102193.8,
  102030.3,
  101955.3,
  101865.7,
  101783.8,
  101953.2,
  102129.1,
  102235.5,
  102453.3,
  102517.5,
  102563.7,
  102433.7,
  102372.4,
  102314.6,
  102386.9,
  102243.4,
  102174,
  101989.3,
  101866.4,
  101741.4,
  101760.8,
  101877.7,
  101847.1,
  101531.7,
  101535.9,
  101476.6,
  101522.9,
  101473.1,
  101453.1,
  101448.7,
  101467.3,
  101150.6,
  101162.4,
  101241.5,
  101463.7,
  101324,
  101408.3,
  101470.7,
  101680.6,
  101665.4,
  101709,
  101347.9,
  100850.7,
  100871.5,
  101193.6,
  101254.1,
  101617.7,
  101829.4,
  101996.5,
  101992,
  102077,
  101880.8,
  101990.1,
  101788.2,
  101589.8,
  101068.9,
  100975.3,
  101039,
  101163.2,
  101225,
  101636.9,
  101882.8,
  102149.2,
  102028.8,
  101774.1,
  101290,
  100983.1,
  100990.7,
  101587.3,
  102067.8,
  102385.3,
  102423.9,
  102498.5,
  102222,
  102031.8,
  101527.1,
  101444,
  101636.1,
  101922,
  102046.5,
  102220.1,
  102209.9,
  102266.1,
  102057.1,
  101731.7,
  101418.5,
  100954.4,
  100511,
  100456.9,
  100517.9,
  100960.9,
  101184.9,
  101501.5,
  101641.7,
  101931.4,
  102178.4,
  102482.3,
  102646.2,
  102801.9,
  102577,
  102190.8,
  101827,
  101734,
  101499.5,
  101760.7,
  101917.6,
  102322.3,
  102667.4,
  103056.4,
  103087,
  103299.6,
  103138,
  102989.4,
  102746.2,
  102674,
  102329.3,
  102204.8,
  102069.1,
  102041.2,
  101816.9,
  101703,
  101455.1,
  101425.3,
  101260.5,
  101446.9,
  101723.6,
  102327.4,
  102668.8,
  102939.1,
  102990.9,
  103079.8,
  103125.2,
  103021,
  102858.3,
  102652.1,
  102302.4,
  102034.4,
  102034.1,
  102136.8,
  102168.9,
  102201,
  102079.8,
  102046.8,
  101809.6,
  101857.5,
  101939.4,
  102047.4,
  101877,
  101754,
  101426.9,
  101197.8,
  100603.9,
  100503.4,
  100952.5,
  101402,
  101620.5,
  101797.8,
  101946,
  102332.2,
  102630.4,
  103109.6,
  103337.6,
  103451,
  103500.1,
  103509.1,
  103321.6,
  103171.7,
  103060.7,
  103151.6,
  103053.4,
  103042.7,
  102811.9,
  102687.2,
  102551.6,
  102574.3,
  102367,
  102217.9,
  102057.9,
  101995.1,
  101816.8,
  102041,
  102138.6,
  102270.3,
  102155.9,
  102199.8,
  102282.5,
  102440.4,
  102394.8,
  102425.7,
  102406.2,
  102612.4,
  102644,
  102746.8,
  102728.2,
  102845,
  102619.2,
  102534.7,
  102470.1,
  102438,
  102091,
  102028.8,
  101995.2,
  102044,
  101816.4,
  101737.6,
  101641.7,
  101646.9,
  101437.1,
  101384.7,
  101299.4,
  101387.8,
  101173.1,
  101109.3,
  100963.8,
  100903.2,
  100870.8,
  101098.2,
  101292,
  101711.8,
  101859,
  102150.9,
  102227.5,
  102475.2,
  102473.3,
  102761.1,
  102889.5,
  103040.3,
  102944.1,
  102975.6,
  102905.2,
  102944.1,
  102761.6,
  102857.9,
  102651.6,
  102607.8,
  102202.6,
  102079.7,
  101712.8,
  101682.7,
  101399.4,
  101327.6,
  101118.3,
  100852.1,
  100401.6,
  100560.7,
  101152.5,
  101429,
  101662.1,
  101827.7,
  102006.9,
  102072,
  101907.3,
  101818.7,
  101845.3,
  101858.3,
  101446.5,
  101446.8,
  101303.8,
  101342.2,
  101273.5,
  101313.4,
  101356.8,
  101446.8,
  101395.9,
  101390,
  101502.3,
  101618.7,
  101501.4,
  101422.7,
  101517.9,
  101782,
  101976.1,
  102265.9,
  102353.9,
  102608.5,
  102617.7,
  102696.6,
  102761.2,
  102930.2,
  102734,
  102643.6,
  102514.6,
  102361.8,
  102088.2,
  101961.7,
  101851.3,
  101643.2,
  101244.1,
  101122.8,
  101288,
  101455.4,
  101466.2,
  101668.3,
  101499.2,
  101786.4,
  101679.3,
  101788.3,
  101894.2,
  102081.4,
  101948.5,
  101887.9,
  101686,
  101844.7,
  101709.3,
  101630.3,
  101494.7,
  101495.2,
  100969.8,
  100787.1,
  100862.4,
  101253.2,
  101437.8,
  101802.4,
  101987.4,
  102330.5,
  102295.4,
  102343,
  102194.6,
  102244.4,
  101715.1,
  101443.2,
  101015.8,
  100890.2,
  100567.8,
  100975.6,
  101120.2,
  101205.2,
  101142.7,
  101082.2,
  100835.9,
  100794.2,
  100905.1,
  101042.1,
  101043.4,
  101186.7,
  101017.5,
  101025.4,
  101073.4,
  101397.1,
  101321.6,
  101579.5,
  101823,
  101958,
  101907.6,
  101862.9,
  101909.2,
  102078.9,
  101906.4,
  101951.9,
  102028.3,
  101999.9,
  101974.2,
  101955.7,
  102082.5,
  102155.1,
  102063,
  102111.2,
  102040.2,
  102204,
  102027.8,
  101894.7,
  101836.6,
  101883.1,
  101541.8,
  101439.7,
  101388.5,
  101155.8,
  100756.7,
  100623.4,
  100886,
  101299,
  101441.8,
  101551.9,
  101876,
  102213.1,
  102028,
  102059.7,
  102001.4,
  102152.7,
  101939.7,
  101910,
  101952.7,
  102005.2,
  101716.1,
  101660.8,
  101596.8,
  101418,
  101184.7,
  101363.3,
  101518.6,
  101234.8,
  101583.6,
  101309,
  101337,
  101221,
  100719.8,
  100465.4,
  100398.4,
  100977.2,
  101231,
  101565.9,
  101750.9,
  102076.6,
  102251.3,
  102341.5,
  102383.1,
  102379.9,
  102106.3,
  101909.6,
  101758.8,
  101727.1,
  101484.2,
  101280.4,
  101362.2,
  101148.8,
  100770.9,
  100384.8,
  100410.7,
  100453.9,
  100542.3,
  100700.1,
  100995.1,
  101268.5,
  101362.8,
  101501.9,
  101671.4,
  101721.5,
  101599.1,
  101518.5,
  101582.7,
  101634.2,
  101533.3,
  101495.1,
  101404.8,
  101412.2,
  101059.6,
  101013.7,
  100833.7,
  100810.2,
  100444.9,
  100188.9,
  99732.97,
  99971.02,
  100058.6,
  100142,
  100323.3,
  100462.1,
  100175.8,
  100192.9,
  100385.6,
  100504.7,
  100661.7,
  100918.4,
  101371.5,
  101708.2,
  101888.3,
  102060.5,
  102233.3,
  102314.5,
  102114.3,
  101980.4,
  101904.5,
  102037,
  101940.9,
  102117.6,
  102209.8,
  102439.2,
  102568.9,
  102563.7,
  102566.5,
  102671,
  102486.8,
  102306.8,
  102254.8,
  102191.4,
  101979,
  101808.2,
  101699.6,
  101790.8,
  101465.3,
  101419.9,
  101320.4,
  101419,
  101169.2,
  101057.9,
  101060.6,
  101006.6,
  100414,
  100480,
  100799.7,
  101218.6,
  100874.3,
  101364.3,
  101480.6,
  101278.1,
  101833.6,
  101641.1,
  101473.5,
  101724,
  101612,
  101571.1,
  101576.8,
  101673.9,
  101390.3,
  101190.2,
  101002.1,
  100793.9,
  100330.5,
  100208.7,
  100126.3,
  100259.3,
  100104,
  100325.6,
  100783.6,
  101353.7,
  101398.1,
  101536.8,
  101849.1,
  102051.5,
  102022.8,
  102074.3,
  102187.3,
  102290,
  102144.1,
  102014.7,
  101955.5,
  102050.2,
  101640.6,
  101432.3,
  101488.6,
  101650.6,
  101546.3,
  101475.3,
  101587.9,
  101608.3,
  101371,
  101387.7,
  101331.9,
  101267.7,
  101024.8,
  101037.6,
  101011.1,
  101102.2,
  100995.1,
  101032.3,
  101135.4,
  101323.2,
  101259.4,
  101201.4,
  101154.5,
  101147.1,
  100966.3,
  100671,
  100585.5,
  100421.9,
  99478.73,
  99242.36,
  99753.55,
  100158.5,
  100250.9,
  100580.4,
  100859.2,
  101072.9,
  100982.1,
  101061.3,
  101280.5,
  101499.9,
  101590.7,
  101787.7,
  101941.9,
  102112.9,
  101926,
  101887.2,
  101913.6,
  102071.2,
  101887,
  101881.2,
  101879.8,
  102022.2,
  101850.3,
  101756.4,
  101798.9,
  101755.7,
  101560.2,
  101451.4,
  101380.5,
  101331.5,
  101080.5,
  100986.6,
  100883.9,
  100939.1,
  100700.8,
  100676,
  100718.6,
  100861.4,
  100677.1,
  100661.2,
  100298,
  100293.5,
  100419.6,
  100520.3,
  100661.1,
  100681.4,
  100527.9,
  100491,
  100773.1,
  101001.1,
  101403.8,
  101770.9,
  101996.8,
  102205,
  102117.7,
  102047,
  101965,
  101821.1,
  101338.2,
  101062.8,
  100879,
  100612,
  100602.6,
  100778.9,
  100912,
  101001.1,
  100878.8,
  100763.3,
  100681.8,
  100836.3,
  100958.8,
  101160.3,
  101310.2,
  101439.3,
  101381.8,
  101304.8,
  101364.2,
  101280.8,
  100992.2,
  100929.6,
  101108.1,
  101413.2,
  101496.8,
  101598.4,
  101758.7,
  101922.6,
  101727.3,
  101622.2,
  101567.9,
  101543,
  101270.2,
  101158.7,
  101194.1,
  101359,
  101221.8,
  101266.1,
  101230,
  101180.9,
  100763.7,
  100593.4,
  100392.1,
  100390.1,
  99873.24,
  99843.04,
  100291.7,
  100725.6,
  100666.3,
  100726.4,
  100790.3,
  100696.9,
  100429.5,
  100192 ;

 time = 0.25, 0.5, 0.75, 1, 1.25, 1.5, 1.75, 2, 2.25, 2.5, 2.75, 3, 3.25, 
    3.5, 3.75, 4, 4.25, 4.5, 4.75, 5, 5.25, 5.5, 5.75, 6, 6.25, 6.5, 6.75, 7, 
    7.25, 7.5, 7.75, 8, 8.25, 8.5, 8.75, 9, 9.25, 9.5, 9.75, 10, 10.25, 10.5, 
    10.75, 11, 11.25, 11.5, 11.75, 12, 12.25, 12.5, 12.75, 13, 13.25, 13.5, 
    13.75, 14, 14.25, 14.5, 14.75, 15, 15.25, 15.5, 15.75, 16, 16.25, 16.5, 
    16.75, 17, 17.25, 17.5, 17.75, 18, 18.25, 18.5, 18.75, 19, 19.25, 19.5, 
    19.75, 20, 20.25, 20.5, 20.75, 21, 21.25, 21.5, 21.75, 22, 22.25, 22.5, 
    22.75, 23, 23.25, 23.5, 23.75, 24, 24.25, 24.5, 24.75, 25, 25.25, 25.5, 
    25.75, 26, 26.25, 26.5, 26.75, 27, 27.25, 27.5, 27.75, 28, 28.25, 28.5, 
    28.75, 29, 29.25, 29.5, 29.75, 30, 30.25, 30.5, 30.75, 31, 31.25, 31.5, 
    31.75, 32, 32.25, 32.5, 32.75, 33, 33.25, 33.5, 33.75, 34, 34.25, 34.5, 
    34.75, 35, 35.25, 35.5, 35.75, 36, 36.25, 36.5, 36.75, 37, 37.25, 37.5, 
    37.75, 38, 38.25, 38.5, 38.75, 39, 39.25, 39.5, 39.75, 40, 40.25, 40.5, 
    40.75, 41, 41.25, 41.5, 41.75, 42, 42.25, 42.5, 42.75, 43, 43.25, 43.5, 
    43.75, 44, 44.25, 44.5, 44.75, 45, 45.25, 45.5, 45.75, 46, 46.25, 46.5, 
    46.75, 47, 47.25, 47.5, 47.75, 48, 48.25, 48.5, 48.75, 49, 49.25, 49.5, 
    49.75, 50, 50.25, 50.5, 50.75, 51, 51.25, 51.5, 51.75, 52, 52.25, 52.5, 
    52.75, 53, 53.25, 53.5, 53.75, 54, 54.25, 54.5, 54.75, 55, 55.25, 55.5, 
    55.75, 56, 56.25, 56.5, 56.75, 57, 57.25, 57.5, 57.75, 58, 58.25, 58.5, 
    58.75, 59, 59.25, 59.5, 59.75, 60, 60.25, 60.5, 60.75, 61, 61.25, 61.5, 
    61.75, 62, 62.25, 62.5, 62.75, 63, 63.25, 63.5, 63.75, 64, 64.25, 64.5, 
    64.75, 65, 65.25, 65.5, 65.75, 66, 66.25, 66.5, 66.75, 67, 67.25, 67.5, 
    67.75, 68, 68.25, 68.5, 68.75, 69, 69.25, 69.5, 69.75, 70, 70.25, 70.5, 
    70.75, 71, 71.25, 71.5, 71.75, 72, 72.25, 72.5, 72.75, 73, 73.25, 73.5, 
    73.75, 74, 74.25, 74.5, 74.75, 75, 75.25, 75.5, 75.75, 76, 76.25, 76.5, 
    76.75, 77, 77.25, 77.5, 77.75, 78, 78.25, 78.5, 78.75, 79, 79.25, 79.5, 
    79.75, 80, 80.25, 80.5, 80.75, 81, 81.25, 81.5, 81.75, 82, 82.25, 82.5, 
    82.75, 83, 83.25, 83.5, 83.75, 84, 84.25, 84.5, 84.75, 85, 85.25, 85.5, 
    85.75, 86, 86.25, 86.5, 86.75, 87, 87.25, 87.5, 87.75, 88, 88.25, 88.5, 
    88.75, 89, 89.25, 89.5, 89.75, 90, 90.25, 90.5, 90.75, 91, 91.25, 91.5, 
    91.75, 92, 92.25, 92.5, 92.75, 93, 93.25, 93.5, 93.75, 94, 94.25, 94.5, 
    94.75, 95, 95.25, 95.5, 95.75, 96, 96.25, 96.5, 96.75, 97, 97.25, 97.5, 
    97.75, 98, 98.25, 98.5, 98.75, 99, 99.25, 99.5, 99.75, 100, 100.25, 
    100.5, 100.75, 101, 101.25, 101.5, 101.75, 102, 102.25, 102.5, 102.75, 
    103, 103.25, 103.5, 103.75, 104, 104.25, 104.5, 104.75, 105, 105.25, 
    105.5, 105.75, 106, 106.25, 106.5, 106.75, 107, 107.25, 107.5, 107.75, 
    108, 108.25, 108.5, 108.75, 109, 109.25, 109.5, 109.75, 110, 110.25, 
    110.5, 110.75, 111, 111.25, 111.5, 111.75, 112, 112.25, 112.5, 112.75, 
    113, 113.25, 113.5, 113.75, 114, 114.25, 114.5, 114.75, 115, 115.25, 
    115.5, 115.75, 116, 116.25, 116.5, 116.75, 117, 117.25, 117.5, 117.75, 
    118, 118.25, 118.5, 118.75, 119, 119.25, 119.5, 119.75, 120, 120.25, 
    120.5, 120.75, 121, 121.25, 121.5, 121.75, 122, 122.25, 122.5, 122.75, 
    123, 123.25, 123.5, 123.75, 124, 124.25, 124.5, 124.75, 125, 125.25, 
    125.5, 125.75, 126, 126.25, 126.5, 126.75, 127, 127.25, 127.5, 127.75, 
    128, 128.25, 128.5, 128.75, 129, 129.25, 129.5, 129.75, 130, 130.25, 
    130.5, 130.75, 131, 131.25, 131.5, 131.75, 132, 132.25, 132.5, 132.75, 
    133, 133.25, 133.5, 133.75, 134, 134.25, 134.5, 134.75, 135, 135.25, 
    135.5, 135.75, 136, 136.25, 136.5, 136.75, 137, 137.25, 137.5, 137.75, 
    138, 138.25, 138.5, 138.75, 139, 139.25, 139.5, 139.75, 140, 140.25, 
    140.5, 140.75, 141, 141.25, 141.5, 141.75, 142, 142.25, 142.5, 142.75, 
    143, 143.25, 143.5, 143.75, 144, 144.25, 144.5, 144.75, 145, 145.25, 
    145.5, 145.75, 146, 146.25, 146.5, 146.75, 147, 147.25, 147.5, 147.75, 
    148, 148.25, 148.5, 148.75, 149, 149.25, 149.5, 149.75, 150, 150.25, 
    150.5, 150.75, 151, 151.25, 151.5, 151.75, 152, 152.25, 152.5, 152.75, 
    153, 153.25, 153.5, 153.75, 154, 154.25, 154.5, 154.75, 155, 155.25, 
    155.5, 155.75, 156, 156.25, 156.5, 156.75, 157, 157.25, 157.5, 157.75, 
    158, 158.25, 158.5, 158.75, 159, 159.25, 159.5, 159.75, 160, 160.25, 
    160.5, 160.75, 161, 161.25, 161.5, 161.75, 162, 162.25, 162.5, 162.75, 
    163, 163.25, 163.5, 163.75, 164, 164.25, 164.5, 164.75, 165, 165.25, 
    165.5, 165.75, 166, 166.25, 166.5, 166.75, 167, 167.25, 167.5, 167.75, 
    168, 168.25, 168.5, 168.75, 169, 169.25, 169.5, 169.75, 170, 170.25, 
    170.5, 170.75, 171, 171.25, 171.5, 171.75, 172, 172.25, 172.5, 172.75, 
    173, 173.25, 173.5, 173.75, 174, 174.25, 174.5, 174.75, 175, 175.25, 
    175.5, 175.75, 176, 176.25, 176.5, 176.75, 177, 177.25, 177.5, 177.75, 
    178, 178.25, 178.5, 178.75, 179, 179.25, 179.5, 179.75, 180, 180.25, 
    180.5, 180.75, 181, 181.25, 181.5, 181.75, 182, 182.25, 182.5, 182.75, 
    183, 183.25, 183.5, 183.75, 184, 184.25, 184.5, 184.75, 185, 185.25, 
    185.5, 185.75, 186, 186.25, 186.5, 186.75, 187, 187.25, 187.5, 187.75, 
    188, 188.25, 188.5, 188.75, 189, 189.25, 189.5, 189.75, 190, 190.25, 
    190.5, 190.75, 191, 191.25, 191.5, 191.75, 192, 192.25, 192.5, 192.75, 
    193, 193.25, 193.5, 193.75, 194, 194.25, 194.5, 194.75, 195, 195.25, 
    195.5, 195.75, 196, 196.25, 196.5, 196.75, 197, 197.25, 197.5, 197.75, 
    198, 198.25, 198.5, 198.75, 199, 199.25, 199.5, 199.75, 200, 200.25, 
    200.5, 200.75, 201, 201.25, 201.5, 201.75, 202, 202.25, 202.5, 202.75, 
    203, 203.25, 203.5, 203.75, 204, 204.25, 204.5, 204.75, 205, 205.25, 
    205.5, 205.75, 206, 206.25, 206.5, 206.75, 207, 207.25, 207.5, 207.75, 
    208, 208.25, 208.5, 208.75, 209, 209.25, 209.5, 209.75, 210, 210.25, 
    210.5, 210.75, 211, 211.25, 211.5, 211.75, 212, 212.25, 212.5, 212.75, 
    213, 213.25, 213.5, 213.75, 214, 214.25, 214.5, 214.75, 215, 215.25, 
    215.5, 215.75, 216, 216.25, 216.5, 216.75, 217, 217.25, 217.5, 217.75, 
    218, 218.25, 218.5, 218.75, 219, 219.25, 219.5, 219.75, 220, 220.25, 
    220.5, 220.75, 221, 221.25, 221.5, 221.75, 222, 222.25, 222.5, 222.75, 
    223, 223.25, 223.5, 223.75, 224, 224.25, 224.5, 224.75, 225, 225.25, 
    225.5, 225.75, 226, 226.25, 226.5, 226.75, 227, 227.25, 227.5, 227.75, 
    228, 228.25, 228.5, 228.75, 229, 229.25, 229.5, 229.75, 230, 230.25, 
    230.5, 230.75, 231, 231.25, 231.5, 231.75, 232, 232.25, 232.5, 232.75, 
    233, 233.25, 233.5, 233.75, 234, 234.25, 234.5, 234.75, 235, 235.25, 
    235.5, 235.75, 236, 236.25, 236.5, 236.75, 237, 237.25, 237.5, 237.75, 
    238, 238.25, 238.5, 238.75, 239, 239.25, 239.5, 239.75, 240, 240.25, 
    240.5, 240.75, 241, 241.25, 241.5, 241.75, 242, 242.25, 242.5, 242.75, 
    243, 243.25, 243.5, 243.75, 244, 244.25, 244.5, 244.75, 245, 245.25, 
    245.5, 245.75, 246, 246.25, 246.5, 246.75, 247, 247.25, 247.5, 247.75, 
    248, 248.25, 248.5, 248.75, 249, 249.25, 249.5, 249.75, 250, 250.25, 
    250.5, 250.75, 251, 251.25, 251.5, 251.75, 252, 252.25, 252.5, 252.75, 
    253, 253.25, 253.5, 253.75, 254, 254.25, 254.5, 254.75, 255, 255.25, 
    255.5, 255.75, 256, 256.25, 256.5, 256.75, 257, 257.25, 257.5, 257.75, 
    258, 258.25, 258.5, 258.75, 259, 259.25, 259.5, 259.75, 260, 260.25, 
    260.5, 260.75, 261, 261.25, 261.5, 261.75, 262, 262.25, 262.5, 262.75, 
    263, 263.25, 263.5, 263.75, 264, 264.25, 264.5, 264.75, 265, 265.25, 
    265.5, 265.75, 266, 266.25, 266.5, 266.75, 267, 267.25, 267.5, 267.75, 
    268, 268.25, 268.5, 268.75, 269, 269.25, 269.5, 269.75, 270, 270.25, 
    270.5, 270.75, 271, 271.25, 271.5, 271.75, 272, 272.25, 272.5, 272.75, 
    273, 273.25, 273.5, 273.75, 274, 274.25, 274.5, 274.75, 275, 275.25, 
    275.5, 275.75, 276, 276.25, 276.5, 276.75, 277, 277.25, 277.5, 277.75, 
    278, 278.25, 278.5, 278.75, 279, 279.25, 279.5, 279.75, 280, 280.25, 
    280.5, 280.75, 281, 281.25, 281.5, 281.75, 282, 282.25, 282.5, 282.75, 
    283, 283.25, 283.5, 283.75, 284, 284.25, 284.5, 284.75, 285, 285.25, 
    285.5, 285.75, 286, 286.25, 286.5, 286.75, 287, 287.25, 287.5, 287.75, 
    288, 288.25, 288.5, 288.75, 289, 289.25, 289.5, 289.75, 290, 290.25, 
    290.5, 290.75, 291, 291.25, 291.5, 291.75, 292, 292.25, 292.5, 292.75, 
    293, 293.25, 293.5, 293.75, 294, 294.25, 294.5, 294.75, 295, 295.25, 
    295.5, 295.75, 296, 296.25, 296.5, 296.75, 297, 297.25, 297.5, 297.75, 
    298, 298.25, 298.5, 298.75, 299, 299.25, 299.5, 299.75, 300, 300.25, 
    300.5, 300.75, 301, 301.25, 301.5, 301.75, 302, 302.25, 302.5, 302.75, 
    303, 303.25, 303.5, 303.75, 304, 304.25, 304.5, 304.75, 305, 305.25, 
    305.5, 305.75, 306, 306.25, 306.5, 306.75, 307, 307.25, 307.5, 307.75, 
    308, 308.25, 308.5, 308.75, 309, 309.25, 309.5, 309.75, 310, 310.25, 
    310.5, 310.75, 311, 311.25, 311.5, 311.75, 312, 312.25, 312.5, 312.75, 
    313, 313.25, 313.5, 313.75, 314, 314.25, 314.5, 314.75, 315, 315.25, 
    315.5, 315.75, 316, 316.25, 316.5, 316.75, 317, 317.25, 317.5, 317.75, 
    318, 318.25, 318.5, 318.75, 319, 319.25, 319.5, 319.75, 320, 320.25, 
    320.5, 320.75, 321, 321.25, 321.5, 321.75, 322, 322.25, 322.5, 322.75, 
    323, 323.25, 323.5, 323.75, 324, 324.25, 324.5, 324.75, 325, 325.25, 
    325.5, 325.75, 326, 326.25, 326.5, 326.75, 327, 327.25, 327.5, 327.75, 
    328, 328.25, 328.5, 328.75, 329, 329.25, 329.5, 329.75, 330, 330.25, 
    330.5, 330.75, 331, 331.25, 331.5, 331.75, 332, 332.25, 332.5, 332.75, 
    333, 333.25, 333.5, 333.75, 334, 334.25, 334.5, 334.75, 335, 335.25, 
    335.5, 335.75, 336, 336.25, 336.5, 336.75, 337, 337.25, 337.5, 337.75, 
    338, 338.25, 338.5, 338.75, 339, 339.25, 339.5, 339.75, 340, 340.25, 
    340.5, 340.75, 341, 341.25, 341.5, 341.75, 342, 342.25, 342.5, 342.75, 
    343, 343.25, 343.5, 343.75, 344, 344.25, 344.5, 344.75, 345, 345.25, 
    345.5, 345.75, 346, 346.25, 346.5, 346.75, 347, 347.25, 347.5, 347.75, 
    348, 348.25, 348.5, 348.75, 349, 349.25, 349.5, 349.75, 350, 350.25, 
    350.5, 350.75, 351, 351.25, 351.5, 351.75, 352, 352.25, 352.5, 352.75, 
    353, 353.25, 353.5, 353.75, 354, 354.25, 354.5, 354.75, 355, 355.25, 
    355.5, 355.75, 356, 356.25, 356.5, 356.75, 357, 357.25, 357.5, 357.75, 
    358, 358.25, 358.5, 358.75, 359, 359.25, 359.5, 359.75, 360, 360.25, 
    360.5, 360.75, 361, 361.25, 361.5, 361.75, 362, 362.25, 362.5, 362.75, 
    363, 363.25, 363.5, 363.75, 364, 364.25, 364.5, 364.75, 365, 365.25, 
    365.5, 365.75, 366, 366.25, 366.5, 366.75, 367, 367.25, 367.5, 367.75, 
    368, 368.25, 368.5, 368.75, 369, 369.25, 369.5, 369.75, 370, 370.25, 
    370.5, 370.75, 371, 371.25, 371.5, 371.75, 372, 372.25, 372.5, 372.75, 
    373, 373.25, 373.5, 373.75, 374, 374.25, 374.5, 374.75, 375, 375.25, 
    375.5, 375.75, 376, 376.25, 376.5, 376.75, 377, 377.25, 377.5, 377.75, 
    378, 378.25, 378.5, 378.75, 379, 379.25, 379.5, 379.75, 380, 380.25, 
    380.5, 380.75, 381, 381.25, 381.5, 381.75, 382, 382.25, 382.5, 382.75, 
    383, 383.25, 383.5, 383.75, 384, 384.25, 384.5, 384.75, 385, 385.25, 
    385.5, 385.75, 386, 386.25, 386.5, 386.75, 387, 387.25, 387.5, 387.75, 
    388, 388.25, 388.5, 388.75, 389, 389.25, 389.5, 389.75, 390, 390.25, 
    390.5, 390.75, 391, 391.25, 391.5, 391.75, 392, 392.25, 392.5, 392.75, 
    393, 393.25, 393.5, 393.75, 394, 394.25, 394.5, 394.75, 395, 395.25, 
    395.5, 395.75, 396, 396.25, 396.5, 396.75, 397, 397.25, 397.5, 397.75, 
    398, 398.25, 398.5, 398.75, 399, 399.25, 399.5, 399.75, 400, 400.25, 
    400.5, 400.75, 401, 401.25, 401.5, 401.75, 402, 402.25, 402.5, 402.75, 
    403, 403.25, 403.5, 403.75, 404, 404.25, 404.5, 404.75, 405, 405.25, 
    405.5, 405.75, 406, 406.25, 406.5, 406.75, 407, 407.25, 407.5, 407.75, 
    408, 408.25, 408.5, 408.75, 409, 409.25, 409.5, 409.75, 410, 410.25, 
    410.5, 410.75, 411, 411.25, 411.5, 411.75, 412, 412.25, 412.5, 412.75, 
    413, 413.25, 413.5, 413.75, 414, 414.25, 414.5, 414.75, 415, 415.25, 
    415.5, 415.75, 416, 416.25, 416.5, 416.75, 417, 417.25, 417.5, 417.75, 
    418, 418.25, 418.5, 418.75, 419, 419.25, 419.5, 419.75, 420, 420.25, 
    420.5, 420.75, 421, 421.25, 421.5, 421.75, 422, 422.25, 422.5, 422.75, 
    423, 423.25, 423.5, 423.75, 424, 424.25, 424.5, 424.75, 425, 425.25, 
    425.5, 425.75, 426, 426.25, 426.5, 426.75, 427, 427.25, 427.5, 427.75, 
    428, 428.25, 428.5, 428.75, 429, 429.25, 429.5, 429.75, 430, 430.25, 
    430.5, 430.75, 431, 431.25, 431.5, 431.75, 432, 432.25, 432.5, 432.75, 
    433, 433.25, 433.5, 433.75, 434, 434.25, 434.5, 434.75, 435, 435.25, 
    435.5, 435.75, 436, 436.25, 436.5, 436.75, 437, 437.25, 437.5, 437.75, 
    438, 438.25, 438.5, 438.75, 439, 439.25, 439.5, 439.75, 440, 440.25, 
    440.5, 440.75, 441, 441.25, 441.5, 441.75, 442, 442.25, 442.5, 442.75, 
    443, 443.25, 443.5, 443.75, 444, 444.25, 444.5, 444.75, 445, 445.25, 
    445.5, 445.75, 446, 446.25, 446.5, 446.75, 447, 447.25, 447.5, 447.75, 
    448, 448.25, 448.5, 448.75, 449, 449.25, 449.5, 449.75, 450, 450.25, 
    450.5, 450.75, 451, 451.25, 451.5, 451.75, 452, 452.25, 452.5, 452.75, 
    453, 453.25, 453.5, 453.75, 454, 454.25, 454.5, 454.75, 455, 455.25, 
    455.5, 455.75, 456, 456.25, 456.5, 456.75, 457, 457.25, 457.5, 457.75, 
    458, 458.25, 458.5, 458.75, 459, 459.25, 459.5, 459.75, 460, 460.25, 
    460.5, 460.75, 461, 461.25, 461.5, 461.75, 462, 462.25, 462.5, 462.75, 
    463, 463.25, 463.5, 463.75, 464, 464.25, 464.5, 464.75, 465, 465.25, 
    465.5, 465.75, 466, 466.25, 466.5, 466.75, 467, 467.25, 467.5, 467.75, 
    468, 468.25, 468.5, 468.75, 469, 469.25, 469.5, 469.75, 470, 470.25, 
    470.5, 470.75, 471, 471.25, 471.5, 471.75, 472, 472.25, 472.5, 472.75, 
    473, 473.25, 473.5, 473.75, 474, 474.25, 474.5, 474.75, 475, 475.25, 
    475.5, 475.75, 476, 476.25, 476.5, 476.75, 477, 477.25, 477.5, 477.75, 
    478, 478.25, 478.5, 478.75, 479, 479.25, 479.5, 479.75, 480, 480.25, 
    480.5, 480.75, 481, 481.25, 481.5, 481.75, 482, 482.25, 482.5, 482.75, 
    483, 483.25, 483.5, 483.75, 484, 484.25, 484.5, 484.75, 485, 485.25, 
    485.5, 485.75, 486, 486.25, 486.5, 486.75, 487, 487.25, 487.5, 487.75, 
    488, 488.25, 488.5, 488.75, 489, 489.25, 489.5, 489.75, 490, 490.25, 
    490.5, 490.75, 491, 491.25, 491.5, 491.75, 492, 492.25, 492.5, 492.75, 
    493, 493.25, 493.5, 493.75, 494, 494.25, 494.5, 494.75, 495, 495.25, 
    495.5, 495.75, 496, 496.25, 496.5, 496.75, 497, 497.25, 497.5, 497.75, 
    498, 498.25, 498.5, 498.75, 499, 499.25, 499.5, 499.75, 500, 500.25, 
    500.5, 500.75, 501, 501.25, 501.5, 501.75, 502, 502.25, 502.5, 502.75, 
    503, 503.25, 503.5, 503.75, 504, 504.25, 504.5, 504.75, 505, 505.25, 
    505.5, 505.75, 506, 506.25, 506.5, 506.75, 507, 507.25, 507.5, 507.75, 
    508, 508.25, 508.5, 508.75, 509, 509.25, 509.5, 509.75, 510, 510.25, 
    510.5, 510.75, 511, 511.25, 511.5, 511.75, 512, 512.25, 512.5, 512.75, 
    513, 513.25, 513.5, 513.75, 514, 514.25, 514.5, 514.75, 515, 515.25, 
    515.5, 515.75, 516, 516.25, 516.5, 516.75, 517, 517.25, 517.5, 517.75, 
    518, 518.25, 518.5, 518.75, 519, 519.25, 519.5, 519.75, 520, 520.25, 
    520.5, 520.75, 521, 521.25, 521.5, 521.75, 522, 522.25, 522.5, 522.75, 
    523, 523.25, 523.5, 523.75, 524, 524.25, 524.5, 524.75, 525, 525.25, 
    525.5, 525.75, 526, 526.25, 526.5, 526.75, 527, 527.25, 527.5, 527.75, 
    528, 528.25, 528.5, 528.75, 529, 529.25, 529.5, 529.75, 530, 530.25, 
    530.5, 530.75, 531, 531.25, 531.5, 531.75, 532, 532.25, 532.5, 532.75, 
    533, 533.25, 533.5, 533.75, 534, 534.25, 534.5, 534.75, 535, 535.25, 
    535.5, 535.75, 536, 536.25, 536.5, 536.75, 537, 537.25, 537.5, 537.75, 
    538, 538.25, 538.5, 538.75, 539, 539.25, 539.5, 539.75, 540, 540.25, 
    540.5, 540.75, 541, 541.25, 541.5, 541.75, 542, 542.25, 542.5, 542.75, 
    543, 543.25, 543.5, 543.75, 544, 544.25, 544.5, 544.75, 545, 545.25, 
    545.5, 545.75, 546, 546.25, 546.5, 546.75, 547, 547.25, 547.5, 547.75, 
    548, 548.25, 548.5, 548.75, 549, 549.25, 549.5, 549.75, 550, 550.25, 
    550.5, 550.75, 551, 551.25, 551.5, 551.75, 552, 552.25, 552.5, 552.75, 
    553, 553.25, 553.5, 553.75, 554, 554.25, 554.5, 554.75, 555, 555.25, 
    555.5, 555.75, 556, 556.25, 556.5, 556.75, 557, 557.25, 557.5, 557.75, 
    558, 558.25, 558.5, 558.75, 559, 559.25, 559.5, 559.75, 560, 560.25, 
    560.5, 560.75, 561, 561.25, 561.5, 561.75, 562, 562.25, 562.5, 562.75, 
    563, 563.25, 563.5, 563.75, 564, 564.25, 564.5, 564.75, 565, 565.25, 
    565.5, 565.75, 566, 566.25, 566.5, 566.75, 567, 567.25, 567.5, 567.75, 
    568, 568.25, 568.5, 568.75, 569, 569.25, 569.5, 569.75, 570, 570.25, 
    570.5, 570.75, 571, 571.25, 571.5, 571.75, 572, 572.25, 572.5, 572.75, 
    573, 573.25, 573.5, 573.75, 574, 574.25, 574.5, 574.75, 575, 575.25, 
    575.5, 575.75, 576, 576.25, 576.5, 576.75, 577, 577.25, 577.5, 577.75, 
    578, 578.25, 578.5, 578.75, 579, 579.25, 579.5, 579.75, 580, 580.25, 
    580.5, 580.75, 581, 581.25, 581.5, 581.75, 582, 582.25, 582.5, 582.75, 
    583, 583.25, 583.5, 583.75, 584, 584.25, 584.5, 584.75, 585, 585.25, 
    585.5, 585.75, 586, 586.25, 586.5, 586.75, 587, 587.25, 587.5, 587.75, 
    588, 588.25, 588.5, 588.75, 589, 589.25, 589.5, 589.75, 590, 590.25, 
    590.5, 590.75, 591, 591.25, 591.5, 591.75, 592, 592.25, 592.5, 592.75, 
    593, 593.25, 593.5, 593.75, 594, 594.25, 594.5, 594.75, 595, 595.25, 
    595.5, 595.75, 596, 596.25, 596.5, 596.75, 597, 597.25, 597.5, 597.75, 
    598, 598.25, 598.5, 598.75, 599, 599.25, 599.5, 599.75, 600, 600.25, 
    600.5, 600.75, 601, 601.25, 601.5, 601.75, 602, 602.25, 602.5, 602.75, 
    603, 603.25, 603.5, 603.75, 604, 604.25, 604.5, 604.75, 605, 605.25, 
    605.5, 605.75, 606, 606.25, 606.5, 606.75, 607, 607.25, 607.5, 607.75, 
    608, 608.25, 608.5, 608.75, 609, 609.25, 609.5, 609.75, 610, 610.25, 
    610.5, 610.75, 611, 611.25, 611.5, 611.75, 612, 612.25, 612.5, 612.75, 
    613, 613.25, 613.5, 613.75, 614, 614.25, 614.5, 614.75, 615, 615.25, 
    615.5, 615.75, 616, 616.25, 616.5, 616.75, 617, 617.25, 617.5, 617.75, 
    618, 618.25, 618.5, 618.75, 619, 619.25, 619.5, 619.75, 620, 620.25, 
    620.5, 620.75, 621, 621.25, 621.5, 621.75, 622, 622.25, 622.5, 622.75, 
    623, 623.25, 623.5, 623.75, 624, 624.25, 624.5, 624.75, 625, 625.25, 
    625.5, 625.75, 626, 626.25, 626.5, 626.75, 627, 627.25, 627.5, 627.75, 
    628, 628.25, 628.5, 628.75, 629, 629.25, 629.5, 629.75, 630, 630.25, 
    630.5, 630.75, 631, 631.25, 631.5, 631.75, 632, 632.25, 632.5, 632.75, 
    633, 633.25, 633.5, 633.75, 634, 634.25, 634.5, 634.75, 635, 635.25, 
    635.5, 635.75, 636, 636.25, 636.5, 636.75, 637, 637.25, 637.5, 637.75, 
    638, 638.25, 638.5, 638.75, 639, 639.25, 639.5, 639.75, 640, 640.25, 
    640.5, 640.75, 641, 641.25, 641.5, 641.75, 642, 642.25, 642.5, 642.75, 
    643, 643.25, 643.5, 643.75, 644, 644.25, 644.5, 644.75, 645, 645.25, 
    645.5, 645.75, 646, 646.25, 646.5, 646.75, 647, 647.25, 647.5, 647.75, 
    648, 648.25, 648.5, 648.75, 649, 649.25, 649.5, 649.75, 650, 650.25, 
    650.5, 650.75, 651, 651.25, 651.5, 651.75, 652, 652.25, 652.5, 652.75, 
    653, 653.25, 653.5, 653.75, 654, 654.25, 654.5, 654.75, 655, 655.25, 
    655.5, 655.75, 656, 656.25, 656.5, 656.75, 657, 657.25, 657.5, 657.75, 
    658, 658.25, 658.5, 658.75, 659, 659.25, 659.5, 659.75, 660, 660.25, 
    660.5, 660.75, 661, 661.25, 661.5, 661.75, 662, 662.25, 662.5, 662.75, 
    663, 663.25, 663.5, 663.75, 664, 664.25, 664.5, 664.75, 665, 665.25, 
    665.5, 665.75, 666, 666.25, 666.5, 666.75, 667, 667.25, 667.5, 667.75, 
    668, 668.25, 668.5, 668.75, 669, 669.25, 669.5, 669.75, 670, 670.25, 
    670.5, 670.75, 671, 671.25, 671.5, 671.75, 672, 672.25, 672.5, 672.75, 
    673, 673.25, 673.5, 673.75, 674, 674.25, 674.5, 674.75, 675, 675.25, 
    675.5, 675.75, 676, 676.25, 676.5, 676.75, 677, 677.25, 677.5, 677.75, 
    678, 678.25, 678.5, 678.75, 679, 679.25, 679.5, 679.75, 680, 680.25, 
    680.5, 680.75, 681, 681.25, 681.5, 681.75, 682, 682.25, 682.5, 682.75, 
    683, 683.25, 683.5, 683.75, 684, 684.25, 684.5, 684.75, 685, 685.25, 
    685.5, 685.75, 686, 686.25, 686.5, 686.75, 687, 687.25, 687.5, 687.75, 
    688, 688.25, 688.5, 688.75, 689, 689.25, 689.5, 689.75, 690, 690.25, 
    690.5, 690.75, 691, 691.25, 691.5, 691.75, 692, 692.25, 692.5, 692.75, 
    693, 693.25, 693.5, 693.75, 694, 694.25, 694.5, 694.75, 695, 695.25, 
    695.5, 695.75, 696, 696.25, 696.5, 696.75, 697, 697.25, 697.5, 697.75, 
    698, 698.25, 698.5, 698.75, 699, 699.25, 699.5, 699.75, 700, 700.25, 
    700.5, 700.75, 701, 701.25, 701.5, 701.75, 702, 702.25, 702.5, 702.75, 
    703, 703.25, 703.5, 703.75, 704, 704.25, 704.5, 704.75, 705, 705.25, 
    705.5, 705.75, 706, 706.25, 706.5, 706.75, 707, 707.25, 707.5, 707.75, 
    708, 708.25, 708.5, 708.75, 709, 709.25, 709.5, 709.75, 710, 710.25, 
    710.5, 710.75, 711, 711.25, 711.5, 711.75, 712, 712.25, 712.5, 712.75, 
    713, 713.25, 713.5, 713.75, 714, 714.25, 714.5, 714.75, 715, 715.25, 
    715.5, 715.75, 716, 716.25, 716.5, 716.75, 717, 717.25, 717.5, 717.75, 
    718, 718.25, 718.5, 718.75, 719, 719.25, 719.5, 719.75, 720, 720.25, 
    720.5, 720.75, 721, 721.25, 721.5, 721.75, 722, 722.25, 722.5, 722.75, 
    723, 723.25, 723.5, 723.75, 724, 724.25, 724.5, 724.75, 725, 725.25, 
    725.5, 725.75, 726, 726.25, 726.5, 726.75, 727, 727.25, 727.5, 727.75, 
    728, 728.25, 728.5, 728.75, 729, 729.25, 729.5, 729.75, 730, 730.25, 
    730.5, 730.75, 731, 731.25, 731.5, 731.75, 732, 732.25, 732.5, 732.75, 
    733, 733.25, 733.5, 733.75, 734, 734.25, 734.5, 734.75, 735, 735.25, 
    735.5, 735.75, 736, 736.25, 736.5, 736.75, 737, 737.25, 737.5, 737.75, 
    738, 738.25, 738.5, 738.75, 739, 739.25, 739.5, 739.75, 740, 740.25, 
    740.5, 740.75, 741, 741.25, 741.5, 741.75, 742, 742.25, 742.5, 742.75, 
    743, 743.25, 743.5, 743.75, 744, 744.25, 744.5, 744.75, 745, 745.25, 
    745.5, 745.75, 746, 746.25, 746.5, 746.75, 747, 747.25, 747.5, 747.75, 
    748, 748.25, 748.5, 748.75, 749, 749.25, 749.5, 749.75, 750, 750.25, 
    750.5, 750.75, 751, 751.25, 751.5, 751.75, 752, 752.25, 752.5, 752.75, 
    753, 753.25, 753.5, 753.75, 754, 754.25, 754.5, 754.75, 755, 755.25, 
    755.5, 755.75, 756, 756.25, 756.5, 756.75, 757, 757.25, 757.5, 757.75, 
    758, 758.25, 758.5, 758.75, 759, 759.25, 759.5, 759.75, 760, 760.25, 
    760.5, 760.75, 761, 761.25, 761.5, 761.75, 762, 762.25, 762.5, 762.75, 
    763, 763.25, 763.5, 763.75, 764, 764.25, 764.5, 764.75, 765, 765.25, 
    765.5, 765.75, 766, 766.25, 766.5, 766.75, 767, 767.25, 767.5, 767.75, 
    768, 768.25, 768.5, 768.75, 769, 769.25, 769.5, 769.75, 770, 770.25, 
    770.5, 770.75, 771, 771.25, 771.5, 771.75, 772, 772.25, 772.5, 772.75, 
    773, 773.25, 773.5, 773.75, 774, 774.25, 774.5, 774.75, 775, 775.25, 
    775.5, 775.75, 776, 776.25, 776.5, 776.75, 777, 777.25, 777.5, 777.75, 
    778, 778.25, 778.5, 778.75, 779, 779.25, 779.5, 779.75, 780, 780.25, 
    780.5, 780.75, 781, 781.25, 781.5, 781.75, 782, 782.25, 782.5, 782.75, 
    783, 783.25, 783.5, 783.75, 784, 784.25, 784.5, 784.75, 785, 785.25, 
    785.5, 785.75, 786, 786.25, 786.5, 786.75, 787, 787.25, 787.5, 787.75, 
    788, 788.25, 788.5, 788.75, 789, 789.25, 789.5, 789.75, 790, 790.25, 
    790.5, 790.75, 791, 791.25, 791.5, 791.75, 792, 792.25, 792.5, 792.75, 
    793, 793.25, 793.5, 793.75, 794, 794.25, 794.5, 794.75, 795, 795.25, 
    795.5, 795.75, 796, 796.25, 796.5, 796.75, 797, 797.25, 797.5, 797.75, 
    798, 798.25, 798.5, 798.75, 799, 799.25, 799.5, 799.75, 800, 800.25, 
    800.5, 800.75, 801, 801.25, 801.5, 801.75, 802, 802.25, 802.5, 802.75, 
    803, 803.25, 803.5, 803.75, 804, 804.25, 804.5, 804.75, 805, 805.25, 
    805.5, 805.75, 806, 806.25, 806.5, 806.75, 807, 807.25, 807.5, 807.75, 
    808, 808.25, 808.5, 808.75, 809, 809.25, 809.5, 809.75, 810, 810.25, 
    810.5, 810.75, 811, 811.25, 811.5, 811.75, 812, 812.25, 812.5, 812.75, 
    813, 813.25, 813.5, 813.75, 814, 814.25, 814.5, 814.75, 815, 815.25, 
    815.5, 815.75, 816, 816.25, 816.5, 816.75, 817, 817.25, 817.5, 817.75, 
    818, 818.25, 818.5, 818.75, 819, 819.25, 819.5, 819.75, 820, 820.25, 
    820.5, 820.75, 821, 821.25, 821.5, 821.75, 822, 822.25, 822.5, 822.75, 
    823, 823.25, 823.5, 823.75, 824, 824.25, 824.5, 824.75, 825, 825.25, 
    825.5, 825.75, 826, 826.25, 826.5, 826.75, 827, 827.25, 827.5, 827.75, 
    828, 828.25, 828.5, 828.75, 829, 829.25, 829.5, 829.75, 830, 830.25, 
    830.5, 830.75, 831, 831.25, 831.5, 831.75, 832, 832.25, 832.5, 832.75, 
    833, 833.25, 833.5, 833.75, 834, 834.25, 834.5, 834.75, 835, 835.25, 
    835.5, 835.75, 836, 836.25, 836.5, 836.75, 837, 837.25, 837.5, 837.75, 
    838, 838.25, 838.5, 838.75, 839, 839.25, 839.5, 839.75, 840, 840.25, 
    840.5, 840.75, 841, 841.25, 841.5, 841.75, 842, 842.25, 842.5, 842.75, 
    843, 843.25, 843.5, 843.75, 844, 844.25, 844.5, 844.75, 845, 845.25, 
    845.5, 845.75, 846, 846.25, 846.5, 846.75, 847, 847.25, 847.5, 847.75, 
    848, 848.25, 848.5, 848.75, 849, 849.25, 849.5, 849.75, 850, 850.25, 
    850.5, 850.75, 851, 851.25, 851.5, 851.75, 852, 852.25, 852.5, 852.75, 
    853, 853.25, 853.5, 853.75, 854, 854.25, 854.5, 854.75, 855, 855.25, 
    855.5, 855.75, 856, 856.25, 856.5, 856.75, 857, 857.25, 857.5, 857.75, 
    858, 858.25, 858.5, 858.75, 859, 859.25, 859.5, 859.75, 860, 860.25, 
    860.5, 860.75, 861, 861.25, 861.5, 861.75, 862, 862.25, 862.5, 862.75, 
    863, 863.25, 863.5, 863.75, 864, 864.25, 864.5, 864.75, 865, 865.25, 
    865.5, 865.75, 866, 866.25, 866.5, 866.75, 867, 867.25, 867.5, 867.75, 
    868, 868.25, 868.5, 868.75, 869, 869.25, 869.5, 869.75, 870, 870.25, 
    870.5, 870.75, 871, 871.25, 871.5, 871.75, 872, 872.25, 872.5, 872.75, 
    873, 873.25, 873.5, 873.75, 874, 874.25, 874.5, 874.75, 875, 875.25, 
    875.5, 875.75, 876, 876.25, 876.5, 876.75, 877, 877.25, 877.5, 877.75, 
    878, 878.25, 878.5, 878.75, 879, 879.25, 879.5, 879.75, 880, 880.25, 
    880.5, 880.75, 881, 881.25, 881.5, 881.75, 882, 882.25, 882.5, 882.75, 
    883, 883.25, 883.5, 883.75, 884, 884.25, 884.5, 884.75, 885, 885.25, 
    885.5, 885.75, 886, 886.25, 886.5, 886.75, 887, 887.25, 887.5, 887.75, 
    888, 888.25, 888.5, 888.75, 889, 889.25, 889.5, 889.75, 890, 890.25, 
    890.5, 890.75, 891, 891.25, 891.5, 891.75, 892, 892.25, 892.5, 892.75, 
    893, 893.25, 893.5, 893.75, 894, 894.25, 894.5, 894.75, 895, 895.25, 
    895.5, 895.75, 896, 896.25, 896.5, 896.75, 897, 897.25, 897.5, 897.75, 
    898, 898.25, 898.5, 898.75, 899, 899.25, 899.5, 899.75, 900, 900.25, 
    900.5, 900.75, 901, 901.25, 901.5, 901.75, 902, 902.25, 902.5, 902.75, 
    903, 903.25, 903.5, 903.75, 904, 904.25, 904.5, 904.75, 905, 905.25, 
    905.5, 905.75, 906, 906.25, 906.5, 906.75, 907, 907.25, 907.5, 907.75, 
    908, 908.25, 908.5, 908.75, 909, 909.25, 909.5, 909.75, 910, 910.25, 
    910.5, 910.75, 911, 911.25, 911.5, 911.75, 912, 912.25, 912.5, 912.75, 
    913, 913.25, 913.5, 913.75, 914, 914.25, 914.5, 914.75, 915, 915.25, 
    915.5, 915.75, 916, 916.25, 916.5, 916.75, 917, 917.25, 917.5, 917.75, 
    918, 918.25, 918.5, 918.75, 919, 919.25, 919.5, 919.75, 920, 920.25, 
    920.5, 920.75, 921, 921.25, 921.5, 921.75, 922, 922.25, 922.5, 922.75, 
    923, 923.25, 923.5, 923.75, 924, 924.25, 924.5, 924.75, 925, 925.25, 
    925.5, 925.75, 926, 926.25, 926.5, 926.75, 927, 927.25, 927.5, 927.75, 
    928, 928.25, 928.5, 928.75, 929, 929.25, 929.5, 929.75, 930, 930.25, 
    930.5, 930.75, 931, 931.25, 931.5, 931.75, 932, 932.25, 932.5, 932.75, 
    933, 933.25, 933.5, 933.75, 934, 934.25, 934.5, 934.75, 935, 935.25, 
    935.5, 935.75, 936, 936.25, 936.5, 936.75, 937, 937.25, 937.5, 937.75, 
    938, 938.25, 938.5, 938.75, 939, 939.25, 939.5, 939.75, 940, 940.25, 
    940.5, 940.75, 941, 941.25, 941.5, 941.75, 942, 942.25, 942.5, 942.75, 
    943, 943.25, 943.5, 943.75, 944, 944.25, 944.5, 944.75, 945, 945.25, 
    945.5, 945.75, 946, 946.25, 946.5, 946.75, 947, 947.25, 947.5, 947.75, 
    948, 948.25, 948.5, 948.75, 949, 949.25, 949.5, 949.75, 950, 950.25, 
    950.5, 950.75, 951, 951.25, 951.5, 951.75, 952, 952.25, 952.5, 952.75, 
    953, 953.25, 953.5, 953.75, 954, 954.25, 954.5, 954.75, 955, 955.25, 
    955.5, 955.75, 956, 956.25, 956.5, 956.75, 957, 957.25, 957.5, 957.75, 
    958, 958.25, 958.5, 958.75, 959, 959.25, 959.5, 959.75, 960, 960.25, 
    960.5, 960.75, 961, 961.25, 961.5, 961.75, 962, 962.25, 962.5, 962.75, 
    963, 963.25, 963.5, 963.75, 964, 964.25, 964.5, 964.75, 965, 965.25, 
    965.5, 965.75, 966, 966.25, 966.5, 966.75, 967, 967.25, 967.5, 967.75, 
    968, 968.25, 968.5, 968.75, 969, 969.25, 969.5, 969.75, 970, 970.25, 
    970.5, 970.75, 971, 971.25, 971.5, 971.75, 972, 972.25, 972.5, 972.75, 
    973, 973.25, 973.5, 973.75, 974, 974.25, 974.5, 974.75, 975, 975.25, 
    975.5, 975.75, 976, 976.25, 976.5, 976.75, 977, 977.25, 977.5, 977.75, 
    978, 978.25, 978.5, 978.75, 979, 979.25, 979.5, 979.75, 980, 980.25, 
    980.5, 980.75, 981, 981.25, 981.5, 981.75, 982, 982.25, 982.5, 982.75, 
    983, 983.25, 983.5, 983.75, 984, 984.25, 984.5, 984.75, 985, 985.25, 
    985.5, 985.75, 986, 986.25, 986.5, 986.75, 987, 987.25, 987.5, 987.75, 
    988, 988.25, 988.5, 988.75, 989, 989.25, 989.5, 989.75, 990, 990.25, 
    990.5, 990.75, 991, 991.25, 991.5, 991.75, 992, 992.25, 992.5, 992.75, 
    993, 993.25, 993.5, 993.75, 994, 994.25, 994.5, 994.75, 995, 995.25, 
    995.5, 995.75, 996, 996.25, 996.5, 996.75, 997, 997.25, 997.5, 997.75, 
    998, 998.25, 998.5, 998.75, 999, 999.25, 999.5, 999.75, 1000, 1000.25, 
    1000.5, 1000.75, 1001, 1001.25, 1001.5, 1001.75, 1002, 1002.25, 1002.5, 
    1002.75, 1003, 1003.25, 1003.5, 1003.75, 1004, 1004.25, 1004.5, 1004.75, 
    1005, 1005.25, 1005.5, 1005.75, 1006, 1006.25, 1006.5, 1006.75, 1007, 
    1007.25, 1007.5, 1007.75, 1008, 1008.25, 1008.5, 1008.75, 1009, 1009.25, 
    1009.5, 1009.75, 1010, 1010.25, 1010.5, 1010.75, 1011, 1011.25, 1011.5, 
    1011.75, 1012, 1012.25, 1012.5, 1012.75, 1013, 1013.25, 1013.5, 1013.75, 
    1014, 1014.25, 1014.5, 1014.75, 1015, 1015.25, 1015.5, 1015.75, 1016, 
    1016.25, 1016.5, 1016.75, 1017, 1017.25, 1017.5, 1017.75, 1018, 1018.25, 
    1018.5, 1018.75, 1019, 1019.25, 1019.5, 1019.75, 1020, 1020.25, 1020.5, 
    1020.75, 1021, 1021.25, 1021.5, 1021.75, 1022, 1022.25, 1022.5, 1022.75, 
    1023, 1023.25, 1023.5, 1023.75, 1024, 1024.25, 1024.5, 1024.75, 1025, 
    1025.25, 1025.5, 1025.75, 1026, 1026.25, 1026.5, 1026.75, 1027, 1027.25, 
    1027.5, 1027.75, 1028, 1028.25, 1028.5, 1028.75, 1029, 1029.25, 1029.5, 
    1029.75, 1030, 1030.25, 1030.5, 1030.75, 1031, 1031.25, 1031.5, 1031.75, 
    1032, 1032.25, 1032.5, 1032.75, 1033, 1033.25, 1033.5, 1033.75, 1034, 
    1034.25, 1034.5, 1034.75, 1035, 1035.25, 1035.5, 1035.75, 1036, 1036.25, 
    1036.5, 1036.75, 1037, 1037.25, 1037.5, 1037.75, 1038, 1038.25, 1038.5, 
    1038.75, 1039, 1039.25, 1039.5, 1039.75, 1040, 1040.25, 1040.5, 1040.75, 
    1041, 1041.25, 1041.5, 1041.75, 1042, 1042.25, 1042.5, 1042.75, 1043, 
    1043.25, 1043.5, 1043.75, 1044, 1044.25, 1044.5, 1044.75, 1045, 1045.25, 
    1045.5, 1045.75, 1046, 1046.25, 1046.5, 1046.75, 1047, 1047.25, 1047.5, 
    1047.75, 1048, 1048.25, 1048.5, 1048.75, 1049, 1049.25, 1049.5, 1049.75, 
    1050, 1050.25, 1050.5, 1050.75, 1051, 1051.25, 1051.5, 1051.75, 1052, 
    1052.25, 1052.5, 1052.75, 1053, 1053.25, 1053.5, 1053.75, 1054, 1054.25, 
    1054.5, 1054.75, 1055, 1055.25, 1055.5, 1055.75, 1056, 1056.25, 1056.5, 
    1056.75, 1057, 1057.25, 1057.5, 1057.75, 1058, 1058.25, 1058.5, 1058.75, 
    1059, 1059.25, 1059.5, 1059.75, 1060, 1060.25, 1060.5, 1060.75, 1061, 
    1061.25, 1061.5, 1061.75, 1062, 1062.25, 1062.5, 1062.75, 1063, 1063.25, 
    1063.5, 1063.75, 1064, 1064.25, 1064.5, 1064.75, 1065, 1065.25, 1065.5, 
    1065.75, 1066, 1066.25, 1066.5, 1066.75, 1067, 1067.25, 1067.5, 1067.75, 
    1068, 1068.25, 1068.5, 1068.75, 1069, 1069.25, 1069.5, 1069.75, 1070, 
    1070.25, 1070.5, 1070.75, 1071, 1071.25, 1071.5, 1071.75, 1072, 1072.25, 
    1072.5, 1072.75, 1073, 1073.25, 1073.5, 1073.75, 1074, 1074.25, 1074.5, 
    1074.75, 1075, 1075.25, 1075.5, 1075.75, 1076, 1076.25, 1076.5, 1076.75, 
    1077, 1077.25, 1077.5, 1077.75, 1078, 1078.25, 1078.5, 1078.75, 1079, 
    1079.25, 1079.5, 1079.75, 1080, 1080.25, 1080.5, 1080.75, 1081, 1081.25, 
    1081.5, 1081.75, 1082, 1082.25, 1082.5, 1082.75, 1083, 1083.25, 1083.5, 
    1083.75, 1084, 1084.25, 1084.5, 1084.75, 1085, 1085.25, 1085.5, 1085.75, 
    1086, 1086.25, 1086.5, 1086.75, 1087, 1087.25, 1087.5, 1087.75, 1088, 
    1088.25, 1088.5, 1088.75, 1089, 1089.25, 1089.5, 1089.75, 1090, 1090.25, 
    1090.5, 1090.75, 1091, 1091.25, 1091.5, 1091.75, 1092, 1092.25, 1092.5, 
    1092.75, 1093, 1093.25, 1093.5, 1093.75, 1094, 1094.25, 1094.5, 1094.75, 
    1095, 1095.25, 1095.5, 1095.75, 1096, 1096.25, 1096.5, 1096.75, 1097, 
    1097.25, 1097.5, 1097.75, 1098, 1098.25, 1098.5, 1098.75, 1099, 1099.25, 
    1099.5, 1099.75, 1100, 1100.25, 1100.5, 1100.75, 1101, 1101.25, 1101.5, 
    1101.75, 1102, 1102.25, 1102.5, 1102.75, 1103, 1103.25, 1103.5, 1103.75, 
    1104, 1104.25, 1104.5, 1104.75, 1105, 1105.25, 1105.5, 1105.75, 1106, 
    1106.25, 1106.5, 1106.75, 1107, 1107.25, 1107.5, 1107.75, 1108, 1108.25, 
    1108.5, 1108.75, 1109, 1109.25, 1109.5, 1109.75, 1110, 1110.25, 1110.5, 
    1110.75, 1111, 1111.25, 1111.5, 1111.75, 1112, 1112.25, 1112.5, 1112.75, 
    1113, 1113.25, 1113.5, 1113.75, 1114, 1114.25, 1114.5, 1114.75, 1115, 
    1115.25, 1115.5, 1115.75, 1116, 1116.25, 1116.5, 1116.75, 1117, 1117.25, 
    1117.5, 1117.75, 1118, 1118.25, 1118.5, 1118.75, 1119, 1119.25, 1119.5, 
    1119.75, 1120, 1120.25, 1120.5, 1120.75, 1121, 1121.25, 1121.5, 1121.75, 
    1122, 1122.25, 1122.5, 1122.75, 1123, 1123.25, 1123.5, 1123.75, 1124, 
    1124.25, 1124.5, 1124.75, 1125, 1125.25, 1125.5, 1125.75, 1126, 1126.25, 
    1126.5, 1126.75, 1127, 1127.25, 1127.5, 1127.75, 1128, 1128.25, 1128.5, 
    1128.75, 1129, 1129.25, 1129.5, 1129.75, 1130, 1130.25, 1130.5, 1130.75, 
    1131, 1131.25, 1131.5, 1131.75, 1132, 1132.25, 1132.5, 1132.75, 1133, 
    1133.25, 1133.5, 1133.75, 1134, 1134.25, 1134.5, 1134.75, 1135, 1135.25, 
    1135.5, 1135.75, 1136, 1136.25, 1136.5, 1136.75, 1137, 1137.25, 1137.5, 
    1137.75, 1138, 1138.25, 1138.5, 1138.75, 1139, 1139.25, 1139.5, 1139.75, 
    1140, 1140.25, 1140.5, 1140.75, 1141, 1141.25, 1141.5, 1141.75, 1142, 
    1142.25, 1142.5, 1142.75, 1143, 1143.25, 1143.5, 1143.75, 1144, 1144.25, 
    1144.5, 1144.75, 1145, 1145.25, 1145.5, 1145.75, 1146, 1146.25, 1146.5, 
    1146.75, 1147, 1147.25, 1147.5, 1147.75, 1148, 1148.25, 1148.5, 1148.75, 
    1149, 1149.25, 1149.5, 1149.75, 1150, 1150.25, 1150.5, 1150.75, 1151, 
    1151.25, 1151.5, 1151.75, 1152, 1152.25, 1152.5, 1152.75, 1153, 1153.25, 
    1153.5, 1153.75, 1154, 1154.25, 1154.5, 1154.75, 1155, 1155.25, 1155.5, 
    1155.75, 1156, 1156.25, 1156.5, 1156.75, 1157, 1157.25, 1157.5, 1157.75, 
    1158, 1158.25, 1158.5, 1158.75, 1159, 1159.25, 1159.5, 1159.75, 1160, 
    1160.25, 1160.5, 1160.75, 1161, 1161.25, 1161.5, 1161.75, 1162, 1162.25, 
    1162.5, 1162.75, 1163, 1163.25, 1163.5, 1163.75, 1164, 1164.25, 1164.5, 
    1164.75, 1165, 1165.25, 1165.5, 1165.75, 1166, 1166.25, 1166.5, 1166.75, 
    1167, 1167.25, 1167.5, 1167.75, 1168, 1168.25, 1168.5, 1168.75, 1169, 
    1169.25, 1169.5, 1169.75, 1170, 1170.25, 1170.5, 1170.75, 1171, 1171.25, 
    1171.5, 1171.75, 1172, 1172.25, 1172.5, 1172.75, 1173, 1173.25, 1173.5, 
    1173.75, 1174, 1174.25, 1174.5, 1174.75, 1175, 1175.25, 1175.5, 1175.75, 
    1176, 1176.25, 1176.5, 1176.75, 1177, 1177.25, 1177.5, 1177.75, 1178, 
    1178.25, 1178.5, 1178.75, 1179, 1179.25, 1179.5, 1179.75, 1180, 1180.25, 
    1180.5, 1180.75, 1181, 1181.25, 1181.5, 1181.75, 1182, 1182.25, 1182.5, 
    1182.75, 1183, 1183.25, 1183.5, 1183.75, 1184, 1184.25, 1184.5, 1184.75, 
    1185, 1185.25, 1185.5, 1185.75, 1186, 1186.25, 1186.5, 1186.75, 1187, 
    1187.25, 1187.5, 1187.75, 1188, 1188.25, 1188.5, 1188.75, 1189, 1189.25, 
    1189.5, 1189.75, 1190, 1190.25, 1190.5, 1190.75, 1191, 1191.25, 1191.5, 
    1191.75, 1192, 1192.25, 1192.5, 1192.75, 1193, 1193.25, 1193.5, 1193.75, 
    1194, 1194.25, 1194.5, 1194.75, 1195, 1195.25, 1195.5, 1195.75, 1196, 
    1196.25, 1196.5, 1196.75, 1197, 1197.25, 1197.5, 1197.75, 1198, 1198.25, 
    1198.5, 1198.75, 1199, 1199.25, 1199.5, 1199.75, 1200, 1200.25, 1200.5, 
    1200.75, 1201, 1201.25, 1201.5, 1201.75, 1202, 1202.25, 1202.5, 1202.75, 
    1203, 1203.25, 1203.5, 1203.75, 1204, 1204.25, 1204.5, 1204.75, 1205, 
    1205.25, 1205.5, 1205.75, 1206, 1206.25, 1206.5, 1206.75, 1207, 1207.25, 
    1207.5, 1207.75, 1208, 1208.25, 1208.5, 1208.75, 1209, 1209.25, 1209.5, 
    1209.75, 1210, 1210.25, 1210.5, 1210.75, 1211, 1211.25, 1211.5, 1211.75, 
    1212, 1212.25, 1212.5, 1212.75, 1213, 1213.25, 1213.5, 1213.75, 1214, 
    1214.25, 1214.5, 1214.75, 1215, 1215.25, 1215.5, 1215.75, 1216, 1216.25, 
    1216.5, 1216.75, 1217, 1217.25, 1217.5, 1217.75, 1218, 1218.25, 1218.5, 
    1218.75, 1219, 1219.25, 1219.5, 1219.75, 1220, 1220.25, 1220.5, 1220.75, 
    1221, 1221.25, 1221.5, 1221.75, 1222, 1222.25, 1222.5, 1222.75, 1223, 
    1223.25, 1223.5, 1223.75, 1224, 1224.25, 1224.5, 1224.75, 1225, 1225.25, 
    1225.5, 1225.75, 1226, 1226.25, 1226.5, 1226.75, 1227, 1227.25, 1227.5, 
    1227.75, 1228, 1228.25, 1228.5, 1228.75, 1229, 1229.25, 1229.5, 1229.75, 
    1230, 1230.25, 1230.5, 1230.75, 1231, 1231.25, 1231.5, 1231.75, 1232, 
    1232.25, 1232.5, 1232.75, 1233, 1233.25, 1233.5, 1233.75, 1234, 1234.25, 
    1234.5, 1234.75, 1235, 1235.25, 1235.5, 1235.75, 1236, 1236.25, 1236.5, 
    1236.75, 1237, 1237.25, 1237.5, 1237.75, 1238, 1238.25, 1238.5, 1238.75, 
    1239, 1239.25, 1239.5, 1239.75, 1240, 1240.25, 1240.5, 1240.75, 1241, 
    1241.25, 1241.5, 1241.75, 1242, 1242.25, 1242.5, 1242.75, 1243, 1243.25, 
    1243.5, 1243.75, 1244, 1244.25, 1244.5, 1244.75, 1245, 1245.25, 1245.5, 
    1245.75, 1246, 1246.25, 1246.5, 1246.75, 1247, 1247.25, 1247.5, 1247.75, 
    1248, 1248.25, 1248.5, 1248.75, 1249, 1249.25, 1249.5, 1249.75, 1250, 
    1250.25, 1250.5, 1250.75, 1251, 1251.25, 1251.5, 1251.75, 1252, 1252.25, 
    1252.5, 1252.75, 1253, 1253.25, 1253.5, 1253.75, 1254, 1254.25, 1254.5, 
    1254.75, 1255, 1255.25, 1255.5, 1255.75, 1256, 1256.25, 1256.5, 1256.75, 
    1257, 1257.25, 1257.5, 1257.75, 1258, 1258.25, 1258.5, 1258.75, 1259, 
    1259.25, 1259.5, 1259.75, 1260, 1260.25, 1260.5, 1260.75, 1261, 1261.25, 
    1261.5, 1261.75, 1262, 1262.25, 1262.5, 1262.75, 1263, 1263.25, 1263.5, 
    1263.75, 1264, 1264.25, 1264.5, 1264.75, 1265, 1265.25, 1265.5, 1265.75, 
    1266, 1266.25, 1266.5, 1266.75, 1267, 1267.25, 1267.5, 1267.75, 1268, 
    1268.25, 1268.5, 1268.75, 1269, 1269.25, 1269.5, 1269.75, 1270, 1270.25, 
    1270.5, 1270.75, 1271, 1271.25, 1271.5, 1271.75, 1272, 1272.25, 1272.5, 
    1272.75, 1273, 1273.25, 1273.5, 1273.75, 1274, 1274.25, 1274.5, 1274.75, 
    1275, 1275.25, 1275.5, 1275.75, 1276, 1276.25, 1276.5, 1276.75, 1277, 
    1277.25, 1277.5, 1277.75, 1278, 1278.25, 1278.5, 1278.75, 1279, 1279.25, 
    1279.5, 1279.75, 1280, 1280.25, 1280.5, 1280.75, 1281, 1281.25, 1281.5, 
    1281.75, 1282, 1282.25, 1282.5, 1282.75, 1283, 1283.25, 1283.5, 1283.75, 
    1284, 1284.25, 1284.5, 1284.75, 1285, 1285.25, 1285.5, 1285.75, 1286, 
    1286.25, 1286.5, 1286.75, 1287, 1287.25, 1287.5, 1287.75, 1288, 1288.25, 
    1288.5, 1288.75, 1289, 1289.25, 1289.5, 1289.75, 1290, 1290.25, 1290.5, 
    1290.75, 1291, 1291.25, 1291.5, 1291.75, 1292, 1292.25, 1292.5, 1292.75, 
    1293, 1293.25, 1293.5, 1293.75, 1294, 1294.25, 1294.5, 1294.75, 1295, 
    1295.25, 1295.5, 1295.75, 1296, 1296.25, 1296.5, 1296.75, 1297, 1297.25, 
    1297.5, 1297.75, 1298, 1298.25, 1298.5, 1298.75, 1299, 1299.25, 1299.5, 
    1299.75, 1300, 1300.25, 1300.5, 1300.75, 1301, 1301.25, 1301.5, 1301.75, 
    1302, 1302.25, 1302.5, 1302.75, 1303, 1303.25, 1303.5, 1303.75, 1304, 
    1304.25, 1304.5, 1304.75, 1305, 1305.25, 1305.5, 1305.75, 1306, 1306.25, 
    1306.5, 1306.75, 1307, 1307.25, 1307.5, 1307.75, 1308, 1308.25, 1308.5, 
    1308.75, 1309, 1309.25, 1309.5, 1309.75, 1310, 1310.25, 1310.5, 1310.75, 
    1311, 1311.25, 1311.5, 1311.75, 1312, 1312.25, 1312.5, 1312.75, 1313, 
    1313.25, 1313.5, 1313.75, 1314, 1314.25, 1314.5, 1314.75, 1315, 1315.25, 
    1315.5, 1315.75, 1316, 1316.25, 1316.5, 1316.75, 1317, 1317.25, 1317.5, 
    1317.75, 1318, 1318.25, 1318.5, 1318.75, 1319, 1319.25, 1319.5, 1319.75, 
    1320, 1320.25, 1320.5, 1320.75, 1321, 1321.25, 1321.5, 1321.75, 1322, 
    1322.25, 1322.5, 1322.75, 1323, 1323.25, 1323.5, 1323.75, 1324, 1324.25, 
    1324.5, 1324.75, 1325, 1325.25, 1325.5, 1325.75, 1326, 1326.25, 1326.5, 
    1326.75, 1327, 1327.25, 1327.5, 1327.75, 1328, 1328.25, 1328.5, 1328.75, 
    1329, 1329.25, 1329.5, 1329.75, 1330, 1330.25, 1330.5, 1330.75, 1331, 
    1331.25, 1331.5, 1331.75, 1332, 1332.25, 1332.5, 1332.75, 1333, 1333.25, 
    1333.5, 1333.75, 1334, 1334.25, 1334.5, 1334.75, 1335, 1335.25, 1335.5, 
    1335.75, 1336, 1336.25, 1336.5, 1336.75, 1337, 1337.25, 1337.5, 1337.75, 
    1338, 1338.25, 1338.5, 1338.75, 1339, 1339.25, 1339.5, 1339.75, 1340, 
    1340.25, 1340.5, 1340.75, 1341, 1341.25, 1341.5, 1341.75, 1342, 1342.25, 
    1342.5, 1342.75, 1343, 1343.25, 1343.5, 1343.75, 1344, 1344.25, 1344.5, 
    1344.75, 1345, 1345.25, 1345.5, 1345.75, 1346, 1346.25, 1346.5, 1346.75, 
    1347, 1347.25, 1347.5, 1347.75, 1348, 1348.25, 1348.5, 1348.75, 1349, 
    1349.25, 1349.5, 1349.75, 1350, 1350.25, 1350.5, 1350.75, 1351, 1351.25, 
    1351.5, 1351.75, 1352, 1352.25, 1352.5, 1352.75, 1353, 1353.25, 1353.5, 
    1353.75, 1354, 1354.25, 1354.5, 1354.75, 1355, 1355.25, 1355.5, 1355.75, 
    1356, 1356.25, 1356.5, 1356.75, 1357, 1357.25, 1357.5, 1357.75, 1358, 
    1358.25, 1358.5, 1358.75, 1359, 1359.25, 1359.5, 1359.75, 1360, 1360.25, 
    1360.5, 1360.75, 1361, 1361.25, 1361.5, 1361.75, 1362, 1362.25, 1362.5, 
    1362.75, 1363, 1363.25, 1363.5, 1363.75, 1364, 1364.25, 1364.5, 1364.75, 
    1365, 1365.25, 1365.5, 1365.75, 1366, 1366.25, 1366.5, 1366.75, 1367, 
    1367.25, 1367.5, 1367.75, 1368, 1368.25, 1368.5, 1368.75, 1369, 1369.25, 
    1369.5, 1369.75, 1370, 1370.25, 1370.5, 1370.75, 1371, 1371.25, 1371.5, 
    1371.75, 1372, 1372.25, 1372.5, 1372.75, 1373, 1373.25, 1373.5, 1373.75, 
    1374, 1374.25, 1374.5, 1374.75, 1375, 1375.25, 1375.5, 1375.75, 1376, 
    1376.25, 1376.5, 1376.75, 1377, 1377.25, 1377.5, 1377.75, 1378, 1378.25, 
    1378.5, 1378.75, 1379, 1379.25, 1379.5, 1379.75, 1380, 1380.25, 1380.5, 
    1380.75, 1381, 1381.25, 1381.5, 1381.75, 1382, 1382.25, 1382.5, 1382.75, 
    1383, 1383.25, 1383.5, 1383.75, 1384, 1384.25, 1384.5, 1384.75, 1385, 
    1385.25, 1385.5, 1385.75, 1386, 1386.25, 1386.5, 1386.75, 1387, 1387.25, 
    1387.5, 1387.75, 1388, 1388.25, 1388.5, 1388.75, 1389, 1389.25, 1389.5, 
    1389.75, 1390, 1390.25, 1390.5, 1390.75, 1391, 1391.25, 1391.5, 1391.75, 
    1392, 1392.25, 1392.5, 1392.75, 1393, 1393.25, 1393.5, 1393.75, 1394, 
    1394.25, 1394.5, 1394.75, 1395, 1395.25, 1395.5, 1395.75, 1396, 1396.25, 
    1396.5, 1396.75, 1397, 1397.25, 1397.5, 1397.75, 1398, 1398.25, 1398.5, 
    1398.75, 1399, 1399.25, 1399.5, 1399.75, 1400, 1400.25, 1400.5, 1400.75, 
    1401, 1401.25, 1401.5, 1401.75, 1402, 1402.25, 1402.5, 1402.75, 1403, 
    1403.25, 1403.5, 1403.75, 1404, 1404.25, 1404.5, 1404.75, 1405, 1405.25, 
    1405.5, 1405.75, 1406, 1406.25, 1406.5, 1406.75, 1407, 1407.25, 1407.5, 
    1407.75, 1408, 1408.25, 1408.5, 1408.75, 1409, 1409.25, 1409.5, 1409.75, 
    1410, 1410.25, 1410.5, 1410.75, 1411, 1411.25, 1411.5, 1411.75, 1412, 
    1412.25, 1412.5, 1412.75, 1413, 1413.25, 1413.5, 1413.75, 1414, 1414.25, 
    1414.5, 1414.75, 1415, 1415.25, 1415.5, 1415.75, 1416, 1416.25, 1416.5, 
    1416.75, 1417, 1417.25, 1417.5, 1417.75, 1418, 1418.25, 1418.5, 1418.75, 
    1419, 1419.25, 1419.5, 1419.75, 1420, 1420.25, 1420.5, 1420.75, 1421, 
    1421.25, 1421.5, 1421.75, 1422, 1422.25, 1422.5, 1422.75, 1423, 1423.25, 
    1423.5, 1423.75, 1424, 1424.25, 1424.5, 1424.75, 1425, 1425.25, 1425.5, 
    1425.75, 1426, 1426.25, 1426.5, 1426.75, 1427, 1427.25, 1427.5, 1427.75, 
    1428, 1428.25, 1428.5, 1428.75, 1429, 1429.25, 1429.5, 1429.75, 1430, 
    1430.25, 1430.5, 1430.75, 1431, 1431.25, 1431.5, 1431.75, 1432, 1432.25, 
    1432.5, 1432.75, 1433, 1433.25, 1433.5, 1433.75, 1434, 1434.25, 1434.5, 
    1434.75, 1435, 1435.25, 1435.5, 1435.75, 1436, 1436.25, 1436.5, 1436.75, 
    1437, 1437.25, 1437.5, 1437.75, 1438, 1438.25, 1438.5, 1438.75, 1439, 
    1439.25, 1439.5, 1439.75, 1440, 1440.25, 1440.5, 1440.75, 1441, 1441.25, 
    1441.5, 1441.75, 1442, 1442.25, 1442.5, 1442.75, 1443, 1443.25, 1443.5, 
    1443.75, 1444, 1444.25, 1444.5, 1444.75, 1445, 1445.25, 1445.5, 1445.75, 
    1446, 1446.25, 1446.5, 1446.75, 1447, 1447.25, 1447.5, 1447.75, 1448, 
    1448.25, 1448.5, 1448.75, 1449, 1449.25, 1449.5, 1449.75, 1450, 1450.25, 
    1450.5, 1450.75, 1451, 1451.25, 1451.5, 1451.75, 1452, 1452.25, 1452.5, 
    1452.75, 1453, 1453.25, 1453.5, 1453.75, 1454, 1454.25, 1454.5, 1454.75, 
    1455, 1455.25, 1455.5, 1455.75, 1456, 1456.25, 1456.5, 1456.75, 1457, 
    1457.25, 1457.5, 1457.75, 1458, 1458.25, 1458.5, 1458.75, 1459, 1459.25, 
    1459.5, 1459.75, 1460, 1460.25, 1460.5, 1460.75, 1461, 1461.25, 1461.5, 
    1461.75, 1462, 1462.25, 1462.5, 1462.75, 1463, 1463.25, 1463.5, 1463.75, 
    1464, 1464.25, 1464.5, 1464.75, 1465, 1465.25, 1465.5, 1465.75, 1466, 
    1466.25, 1466.5, 1466.75, 1467, 1467.25, 1467.5, 1467.75, 1468, 1468.25, 
    1468.5, 1468.75, 1469, 1469.25, 1469.5, 1469.75, 1470, 1470.25, 1470.5, 
    1470.75, 1471, 1471.25, 1471.5, 1471.75, 1472, 1472.25, 1472.5, 1472.75, 
    1473, 1473.25, 1473.5, 1473.75, 1474, 1474.25, 1474.5, 1474.75, 1475, 
    1475.25, 1475.5, 1475.75, 1476, 1476.25, 1476.5, 1476.75, 1477, 1477.25, 
    1477.5, 1477.75, 1478, 1478.25, 1478.5, 1478.75, 1479, 1479.25, 1479.5, 
    1479.75, 1480, 1480.25, 1480.5, 1480.75, 1481, 1481.25, 1481.5, 1481.75, 
    1482, 1482.25, 1482.5, 1482.75, 1483, 1483.25, 1483.5, 1483.75, 1484, 
    1484.25, 1484.5, 1484.75, 1485, 1485.25, 1485.5, 1485.75, 1486, 1486.25, 
    1486.5, 1486.75, 1487, 1487.25, 1487.5, 1487.75, 1488, 1488.25, 1488.5, 
    1488.75, 1489, 1489.25, 1489.5, 1489.75, 1490, 1490.25, 1490.5, 1490.75, 
    1491, 1491.25, 1491.5, 1491.75, 1492, 1492.25, 1492.5, 1492.75, 1493, 
    1493.25, 1493.5, 1493.75, 1494, 1494.25, 1494.5, 1494.75, 1495, 1495.25, 
    1495.5, 1495.75, 1496, 1496.25, 1496.5, 1496.75, 1497, 1497.25, 1497.5, 
    1497.75, 1498, 1498.25, 1498.5, 1498.75, 1499, 1499.25, 1499.5, 1499.75, 
    1500, 1500.25, 1500.5, 1500.75, 1501, 1501.25, 1501.5, 1501.75, 1502, 
    1502.25, 1502.5, 1502.75, 1503, 1503.25, 1503.5, 1503.75, 1504, 1504.25, 
    1504.5, 1504.75, 1505, 1505.25, 1505.5, 1505.75, 1506, 1506.25, 1506.5, 
    1506.75, 1507, 1507.25, 1507.5, 1507.75, 1508, 1508.25, 1508.5, 1508.75, 
    1509, 1509.25, 1509.5, 1509.75, 1510, 1510.25, 1510.5, 1510.75, 1511, 
    1511.25, 1511.5, 1511.75, 1512, 1512.25, 1512.5, 1512.75, 1513, 1513.25, 
    1513.5, 1513.75, 1514, 1514.25, 1514.5, 1514.75, 1515, 1515.25, 1515.5, 
    1515.75, 1516, 1516.25, 1516.5, 1516.75, 1517, 1517.25, 1517.5, 1517.75, 
    1518, 1518.25, 1518.5, 1518.75, 1519, 1519.25, 1519.5, 1519.75, 1520, 
    1520.25, 1520.5, 1520.75, 1521, 1521.25, 1521.5, 1521.75, 1522, 1522.25, 
    1522.5, 1522.75, 1523, 1523.25, 1523.5, 1523.75, 1524, 1524.25, 1524.5, 
    1524.75, 1525, 1525.25, 1525.5, 1525.75, 1526, 1526.25, 1526.5, 1526.75, 
    1527, 1527.25, 1527.5, 1527.75, 1528, 1528.25, 1528.5, 1528.75, 1529, 
    1529.25, 1529.5, 1529.75, 1530, 1530.25, 1530.5, 1530.75, 1531, 1531.25, 
    1531.5, 1531.75, 1532, 1532.25, 1532.5, 1532.75, 1533, 1533.25, 1533.5, 
    1533.75, 1534, 1534.25, 1534.5, 1534.75, 1535, 1535.25, 1535.5, 1535.75, 
    1536, 1536.25, 1536.5, 1536.75, 1537, 1537.25, 1537.5, 1537.75, 1538, 
    1538.25, 1538.5, 1538.75, 1539, 1539.25, 1539.5, 1539.75, 1540, 1540.25, 
    1540.5, 1540.75, 1541, 1541.25, 1541.5, 1541.75, 1542, 1542.25, 1542.5, 
    1542.75, 1543, 1543.25, 1543.5, 1543.75, 1544, 1544.25, 1544.5, 1544.75, 
    1545, 1545.25, 1545.5, 1545.75, 1546, 1546.25, 1546.5, 1546.75, 1547, 
    1547.25, 1547.5, 1547.75, 1548, 1548.25, 1548.5, 1548.75, 1549, 1549.25, 
    1549.5, 1549.75, 1550, 1550.25, 1550.5, 1550.75, 1551, 1551.25, 1551.5, 
    1551.75, 1552, 1552.25, 1552.5, 1552.75, 1553, 1553.25, 1553.5, 1553.75, 
    1554, 1554.25, 1554.5, 1554.75, 1555, 1555.25, 1555.5, 1555.75, 1556, 
    1556.25, 1556.5, 1556.75, 1557, 1557.25, 1557.5, 1557.75, 1558, 1558.25, 
    1558.5, 1558.75, 1559, 1559.25, 1559.5, 1559.75, 1560, 1560.25, 1560.5, 
    1560.75, 1561, 1561.25, 1561.5, 1561.75, 1562, 1562.25, 1562.5, 1562.75, 
    1563, 1563.25, 1563.5, 1563.75, 1564, 1564.25, 1564.5, 1564.75, 1565, 
    1565.25, 1565.5, 1565.75, 1566, 1566.25, 1566.5, 1566.75, 1567, 1567.25, 
    1567.5, 1567.75, 1568, 1568.25, 1568.5, 1568.75, 1569, 1569.25, 1569.5, 
    1569.75, 1570, 1570.25, 1570.5, 1570.75, 1571, 1571.25, 1571.5, 1571.75, 
    1572, 1572.25, 1572.5, 1572.75, 1573, 1573.25, 1573.5, 1573.75, 1574, 
    1574.25, 1574.5, 1574.75, 1575, 1575.25, 1575.5, 1575.75, 1576, 1576.25, 
    1576.5, 1576.75, 1577, 1577.25, 1577.5, 1577.75, 1578, 1578.25, 1578.5, 
    1578.75, 1579, 1579.25, 1579.5, 1579.75, 1580, 1580.25, 1580.5, 1580.75, 
    1581, 1581.25, 1581.5, 1581.75, 1582, 1582.25, 1582.5, 1582.75, 1583, 
    1583.25, 1583.5, 1583.75, 1584, 1584.25, 1584.5, 1584.75, 1585, 1585.25, 
    1585.5, 1585.75, 1586, 1586.25, 1586.5, 1586.75, 1587, 1587.25, 1587.5, 
    1587.75, 1588, 1588.25, 1588.5, 1588.75, 1589, 1589.25, 1589.5, 1589.75, 
    1590, 1590.25, 1590.5, 1590.75, 1591, 1591.25, 1591.5, 1591.75, 1592, 
    1592.25, 1592.5, 1592.75, 1593, 1593.25, 1593.5, 1593.75, 1594, 1594.25, 
    1594.5, 1594.75, 1595, 1595.25, 1595.5, 1595.75, 1596, 1596.25, 1596.5, 
    1596.75, 1597, 1597.25, 1597.5, 1597.75, 1598, 1598.25, 1598.5, 1598.75, 
    1599, 1599.25, 1599.5, 1599.75, 1600, 1600.25, 1600.5, 1600.75, 1601, 
    1601.25, 1601.5, 1601.75, 1602, 1602.25, 1602.5, 1602.75, 1603, 1603.25, 
    1603.5, 1603.75, 1604, 1604.25, 1604.5, 1604.75, 1605, 1605.25, 1605.5, 
    1605.75, 1606, 1606.25, 1606.5, 1606.75, 1607, 1607.25, 1607.5, 1607.75, 
    1608, 1608.25, 1608.5, 1608.75, 1609, 1609.25, 1609.5, 1609.75, 1610, 
    1610.25, 1610.5, 1610.75, 1611, 1611.25, 1611.5, 1611.75, 1612, 1612.25, 
    1612.5, 1612.75, 1613, 1613.25, 1613.5, 1613.75, 1614, 1614.25, 1614.5, 
    1614.75, 1615, 1615.25, 1615.5, 1615.75, 1616, 1616.25, 1616.5, 1616.75, 
    1617, 1617.25, 1617.5, 1617.75, 1618, 1618.25, 1618.5, 1618.75, 1619, 
    1619.25, 1619.5, 1619.75, 1620, 1620.25, 1620.5, 1620.75, 1621, 1621.25, 
    1621.5, 1621.75, 1622, 1622.25, 1622.5, 1622.75, 1623, 1623.25, 1623.5, 
    1623.75, 1624, 1624.25, 1624.5, 1624.75, 1625, 1625.25, 1625.5, 1625.75, 
    1626, 1626.25, 1626.5, 1626.75, 1627, 1627.25, 1627.5, 1627.75, 1628, 
    1628.25, 1628.5, 1628.75, 1629, 1629.25, 1629.5, 1629.75, 1630, 1630.25, 
    1630.5, 1630.75, 1631, 1631.25, 1631.5, 1631.75, 1632, 1632.25, 1632.5, 
    1632.75, 1633, 1633.25, 1633.5, 1633.75, 1634, 1634.25, 1634.5, 1634.75, 
    1635, 1635.25, 1635.5, 1635.75, 1636, 1636.25, 1636.5, 1636.75, 1637, 
    1637.25, 1637.5, 1637.75, 1638, 1638.25, 1638.5, 1638.75, 1639, 1639.25, 
    1639.5, 1639.75, 1640, 1640.25, 1640.5, 1640.75, 1641, 1641.25, 1641.5, 
    1641.75, 1642, 1642.25, 1642.5, 1642.75, 1643, 1643.25, 1643.5, 1643.75, 
    1644, 1644.25, 1644.5, 1644.75, 1645, 1645.25, 1645.5, 1645.75, 1646, 
    1646.25, 1646.5, 1646.75, 1647, 1647.25, 1647.5, 1647.75, 1648, 1648.25, 
    1648.5, 1648.75, 1649, 1649.25, 1649.5, 1649.75, 1650, 1650.25, 1650.5, 
    1650.75, 1651, 1651.25, 1651.5, 1651.75, 1652, 1652.25, 1652.5, 1652.75, 
    1653, 1653.25, 1653.5, 1653.75, 1654, 1654.25, 1654.5, 1654.75, 1655, 
    1655.25, 1655.5, 1655.75, 1656, 1656.25, 1656.5, 1656.75, 1657, 1657.25, 
    1657.5, 1657.75, 1658, 1658.25, 1658.5, 1658.75, 1659, 1659.25, 1659.5, 
    1659.75, 1660, 1660.25, 1660.5, 1660.75, 1661, 1661.25, 1661.5, 1661.75, 
    1662, 1662.25, 1662.5, 1662.75, 1663, 1663.25, 1663.5, 1663.75, 1664, 
    1664.25, 1664.5, 1664.75, 1665, 1665.25, 1665.5, 1665.75, 1666, 1666.25, 
    1666.5, 1666.75, 1667, 1667.25, 1667.5, 1667.75, 1668, 1668.25, 1668.5, 
    1668.75, 1669, 1669.25, 1669.5, 1669.75, 1670, 1670.25, 1670.5, 1670.75, 
    1671, 1671.25, 1671.5, 1671.75, 1672, 1672.25, 1672.5, 1672.75, 1673, 
    1673.25, 1673.5, 1673.75, 1674, 1674.25, 1674.5, 1674.75, 1675, 1675.25, 
    1675.5, 1675.75, 1676, 1676.25, 1676.5, 1676.75, 1677, 1677.25, 1677.5, 
    1677.75, 1678, 1678.25, 1678.5, 1678.75, 1679, 1679.25, 1679.5, 1679.75, 
    1680, 1680.25, 1680.5, 1680.75, 1681, 1681.25, 1681.5, 1681.75, 1682, 
    1682.25, 1682.5, 1682.75, 1683, 1683.25, 1683.5, 1683.75, 1684, 1684.25, 
    1684.5, 1684.75, 1685, 1685.25, 1685.5, 1685.75, 1686, 1686.25, 1686.5, 
    1686.75, 1687, 1687.25, 1687.5, 1687.75, 1688, 1688.25, 1688.5, 1688.75, 
    1689, 1689.25, 1689.5, 1689.75, 1690, 1690.25, 1690.5, 1690.75, 1691, 
    1691.25, 1691.5, 1691.75, 1692, 1692.25, 1692.5, 1692.75, 1693, 1693.25, 
    1693.5, 1693.75, 1694, 1694.25, 1694.5, 1694.75, 1695, 1695.25, 1695.5, 
    1695.75, 1696, 1696.25, 1696.5, 1696.75, 1697, 1697.25, 1697.5, 1697.75, 
    1698, 1698.25, 1698.5, 1698.75, 1699, 1699.25, 1699.5, 1699.75, 1700, 
    1700.25, 1700.5, 1700.75, 1701, 1701.25, 1701.5, 1701.75, 1702, 1702.25, 
    1702.5, 1702.75, 1703, 1703.25, 1703.5, 1703.75, 1704, 1704.25, 1704.5, 
    1704.75, 1705, 1705.25, 1705.5, 1705.75, 1706, 1706.25, 1706.5, 1706.75, 
    1707, 1707.25, 1707.5, 1707.75, 1708, 1708.25, 1708.5, 1708.75, 1709, 
    1709.25, 1709.5, 1709.75, 1710, 1710.25, 1710.5, 1710.75, 1711, 1711.25, 
    1711.5, 1711.75, 1712, 1712.25, 1712.5, 1712.75, 1713, 1713.25, 1713.5, 
    1713.75, 1714, 1714.25, 1714.5, 1714.75, 1715, 1715.25, 1715.5, 1715.75, 
    1716, 1716.25, 1716.5, 1716.75, 1717, 1717.25, 1717.5, 1717.75, 1718, 
    1718.25, 1718.5, 1718.75, 1719, 1719.25, 1719.5, 1719.75, 1720, 1720.25, 
    1720.5, 1720.75, 1721, 1721.25, 1721.5, 1721.75, 1722, 1722.25, 1722.5, 
    1722.75, 1723, 1723.25, 1723.5, 1723.75, 1724, 1724.25, 1724.5, 1724.75, 
    1725, 1725.25, 1725.5, 1725.75, 1726, 1726.25, 1726.5, 1726.75, 1727, 
    1727.25, 1727.5, 1727.75, 1728, 1728.25, 1728.5, 1728.75, 1729, 1729.25, 
    1729.5, 1729.75, 1730, 1730.25, 1730.5, 1730.75, 1731, 1731.25, 1731.5, 
    1731.75, 1732, 1732.25, 1732.5, 1732.75, 1733, 1733.25, 1733.5, 1733.75, 
    1734, 1734.25, 1734.5, 1734.75, 1735, 1735.25, 1735.5, 1735.75, 1736, 
    1736.25, 1736.5, 1736.75, 1737, 1737.25, 1737.5, 1737.75, 1738, 1738.25, 
    1738.5, 1738.75, 1739, 1739.25, 1739.5, 1739.75, 1740, 1740.25, 1740.5, 
    1740.75, 1741, 1741.25, 1741.5, 1741.75, 1742, 1742.25, 1742.5, 1742.75, 
    1743, 1743.25, 1743.5, 1743.75, 1744, 1744.25, 1744.5, 1744.75, 1745, 
    1745.25, 1745.5, 1745.75, 1746, 1746.25, 1746.5, 1746.75, 1747, 1747.25, 
    1747.5, 1747.75, 1748, 1748.25, 1748.5, 1748.75, 1749, 1749.25, 1749.5, 
    1749.75, 1750, 1750.25, 1750.5, 1750.75, 1751, 1751.25, 1751.5, 1751.75, 
    1752, 1752.25, 1752.5, 1752.75, 1753, 1753.25, 1753.5, 1753.75, 1754, 
    1754.25, 1754.5, 1754.75, 1755, 1755.25, 1755.5, 1755.75, 1756, 1756.25, 
    1756.5, 1756.75, 1757, 1757.25, 1757.5, 1757.75, 1758, 1758.25, 1758.5, 
    1758.75, 1759, 1759.25, 1759.5, 1759.75, 1760, 1760.25, 1760.5, 1760.75, 
    1761, 1761.25, 1761.5, 1761.75, 1762, 1762.25, 1762.5, 1762.75, 1763, 
    1763.25, 1763.5, 1763.75, 1764, 1764.25, 1764.5, 1764.75, 1765, 1765.25, 
    1765.5, 1765.75, 1766, 1766.25, 1766.5, 1766.75, 1767, 1767.25, 1767.5, 
    1767.75, 1768, 1768.25, 1768.5, 1768.75, 1769, 1769.25, 1769.5, 1769.75, 
    1770, 1770.25, 1770.5, 1770.75, 1771, 1771.25, 1771.5, 1771.75, 1772, 
    1772.25, 1772.5, 1772.75, 1773, 1773.25, 1773.5, 1773.75, 1774, 1774.25, 
    1774.5, 1774.75, 1775, 1775.25, 1775.5, 1775.75, 1776, 1776.25, 1776.5, 
    1776.75, 1777, 1777.25, 1777.5, 1777.75, 1778, 1778.25, 1778.5, 1778.75, 
    1779, 1779.25, 1779.5, 1779.75, 1780, 1780.25, 1780.5, 1780.75, 1781, 
    1781.25, 1781.5, 1781.75, 1782, 1782.25, 1782.5, 1782.75, 1783, 1783.25, 
    1783.5, 1783.75, 1784, 1784.25, 1784.5, 1784.75, 1785, 1785.25, 1785.5, 
    1785.75, 1786, 1786.25, 1786.5, 1786.75, 1787, 1787.25, 1787.5, 1787.75, 
    1788, 1788.25, 1788.5, 1788.75, 1789, 1789.25, 1789.5, 1789.75, 1790, 
    1790.25, 1790.5, 1790.75, 1791, 1791.25, 1791.5, 1791.75, 1792, 1792.25, 
    1792.5, 1792.75, 1793, 1793.25, 1793.5, 1793.75, 1794, 1794.25, 1794.5, 
    1794.75, 1795, 1795.25, 1795.5, 1795.75, 1796, 1796.25, 1796.5, 1796.75, 
    1797, 1797.25, 1797.5, 1797.75, 1798, 1798.25, 1798.5, 1798.75, 1799, 
    1799.25, 1799.5, 1799.75, 1800, 1800.25, 1800.5, 1800.75, 1801, 1801.25, 
    1801.5, 1801.75, 1802, 1802.25, 1802.5, 1802.75, 1803, 1803.25, 1803.5, 
    1803.75, 1804, 1804.25, 1804.5, 1804.75, 1805, 1805.25, 1805.5, 1805.75, 
    1806, 1806.25, 1806.5, 1806.75, 1807, 1807.25, 1807.5, 1807.75, 1808, 
    1808.25, 1808.5, 1808.75, 1809, 1809.25, 1809.5, 1809.75, 1810, 1810.25, 
    1810.5, 1810.75, 1811, 1811.25, 1811.5, 1811.75, 1812, 1812.25, 1812.5, 
    1812.75, 1813, 1813.25, 1813.5, 1813.75, 1814, 1814.25, 1814.5, 1814.75, 
    1815, 1815.25, 1815.5, 1815.75, 1816, 1816.25, 1816.5, 1816.75, 1817, 
    1817.25, 1817.5, 1817.75, 1818, 1818.25, 1818.5, 1818.75, 1819, 1819.25, 
    1819.5, 1819.75, 1820, 1820.25, 1820.5, 1820.75, 1821, 1821.25, 1821.5, 
    1821.75, 1822, 1822.25, 1822.5, 1822.75, 1823, 1823.25, 1823.5, 1823.75, 
    1824, 1824.25, 1824.5, 1824.75, 1825 ;
}
