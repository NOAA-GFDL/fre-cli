netcdf \20030101.grid_spec.tile2 {
dimensions:
	grid_x = 97 ;
	grid_y = 97 ;
	time = UNLIMITED ; // (1 currently)
	grid_xt = 96 ;
	grid_yt = 96 ;
	phalf = 50 ;
variables:
	double grid_x(grid_x) ;
		grid_x:units = "degrees_E" ;
		grid_x:long_name = "cell corner longitude" ;
		grid_x:axis = "X" ;
	double grid_y(grid_y) ;
		grid_y:units = "degrees_N" ;
		grid_y:long_name = "cell corner latitude" ;
		grid_y:axis = "Y" ;
	double time(time) ;
		time:units = "days since 1870-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "JULIAN" ;
		time:calendar = "julian" ;
	double grid_xt(grid_xt) ;
		grid_xt:units = "degrees_E" ;
		grid_xt:long_name = "T-cell longitude" ;
		grid_xt:axis = "X" ;
	double grid_yt(grid_yt) ;
		grid_yt:units = "degrees_N" ;
		grid_yt:long_name = "T-cell latitude" ;
		grid_yt:axis = "Y" ;
	double phalf(phalf) ;
		phalf:units = "mb" ;
		phalf:long_name = "ref half pressure level" ;
		phalf:axis = "Z" ;
		phalf:positive = "down" ;
	float grid_lon(grid_y, grid_x) ;
		grid_lon:_FillValue = 1.e+20f ;
		grid_lon:missing_value = 1.e+20f ;
		grid_lon:units = "degrees_E" ;
		grid_lon:long_name = "longitude" ;
		grid_lon:cell_methods = "time: point" ;
	float grid_lat(grid_y, grid_x) ;
		grid_lat:_FillValue = 1.e+20f ;
		grid_lat:missing_value = 1.e+20f ;
		grid_lat:units = "degrees_N" ;
		grid_lat:long_name = "latitude" ;
		grid_lat:cell_methods = "time: point" ;
	float grid_lont(grid_yt, grid_xt) ;
		grid_lont:_FillValue = 1.e+20f ;
		grid_lont:missing_value = 1.e+20f ;
		grid_lont:units = "degrees_E" ;
		grid_lont:long_name = "longitude" ;
		grid_lont:cell_methods = "time: point" ;
	float grid_latt(grid_yt, grid_xt) ;
		grid_latt:_FillValue = 1.e+20f ;
		grid_latt:missing_value = 1.e+20f ;
		grid_latt:units = "degrees_N" ;
		grid_latt:long_name = "latitude" ;
		grid_latt:cell_methods = "time: point" ;
	float area(grid_yt, grid_xt) ;
		area:_FillValue = 1.e+20f ;
		area:missing_value = 1.e+20f ;
		area:units = "m**2" ;
		area:long_name = "cell area" ;
		area:cell_methods = "time: point" ;
	float bk(phalf) ;
		bk:_FillValue = 1.e+20f ;
		bk:missing_value = 1.e+20f ;
		bk:long_name = "vertical coordinate sigma value" ;
		bk:cell_methods = "time: point" ;
	float pk(phalf) ;
		pk:_FillValue = 1.e+20f ;
		pk:missing_value = 1.e+20f ;
		pk:units = "pascal" ;
		pk:long_name = "pressure part of the hybrid coordinate" ;
		pk:cell_methods = "time: point" ;
	float sftlf(grid_yt, grid_xt) ;
		sftlf:_FillValue = 1.e+20f ;
		sftlf:missing_value = 1.e+20f ;
		sftlf:units = "1.0" ;
		sftlf:long_name = "Fraction of the Grid Cell Occupied by Land" ;
		sftlf:cell_methods = "time: point" ;
		sftlf:cell_measures = "area: area" ;
		sftlf:standard_name = "land_area_fraction" ;
		sftlf:interp_method = "conserve_order1" ;
	float orog(grid_yt, grid_xt) ;
		orog:_FillValue = 1.e+20f ;
		orog:missing_value = 1.e+20f ;
		orog:units = "m" ;
		orog:long_name = "Surface Altitude" ;
		orog:cell_methods = "time: point" ;
		orog:cell_measures = "area: area" ;
		orog:standard_name = "surface_altitude" ;
		orog:interp_method = "conserve_order1" ;
	float land_mask(grid_yt, grid_xt) ;
		land_mask:_FillValue = 1.e+20f ;
		land_mask:missing_value = 1.e+20f ;
		land_mask:valid_range = -0.01f, 1.01f ;
		land_mask:long_name = "fractional amount of land" ;
		land_mask:cell_methods = "time: point" ;
		land_mask:interp_method = "conserve_order1" ;
	float zsurf(grid_yt, grid_xt) ;
		zsurf:_FillValue = 1.e+20f ;
		zsurf:missing_value = 1.e+20f ;
		zsurf:units = "m" ;
		zsurf:long_name = "surface height" ;
		zsurf:cell_methods = "time: point" ;

// global attributes:
		:title = "ESM4_longamip_D1_am4p2_proto7b_whiteCapsAlbedo_salt_SIS2" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
data:

 grid_x = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 
    20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 
    38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 
    56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 73, 
    74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 
    92, 93, 94, 95, 96, 97 ;

 grid_y = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 
    20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 
    38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 
    56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 73, 
    74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 
    92, 93, 94, 95, 96, 97 ;

 time = 0 ;

 grid_xt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 
    20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 
    38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 
    56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 73, 
    74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 
    92, 93, 94, 95, 96 ;

 grid_yt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 
    20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 
    38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 
    56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 73, 
    74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 
    92, 93, 94, 95, 96 ;

 phalf = 0.01, 0.0269722, 0.0517136, 0.0889455, 0.142479, 0.2207157, 
    0.3361283, 0.5048096, 0.7479993, 1.0940055, 1.580046, 2.2544108, 
    3.178956, 4.431935, 6.1111558, 8.3374392, 11.2583405, 15.0520759, 
    19.9315829, 26.1486254, 33.997842, 43.820624, 56.0087014, 71.0073115, 
    89.3178242, 111.4997021, 138.1716841, 170.012093, 207.7581856, 
    252.2033875, 304.1464563, 363.9522552, 430.6429622, 501.015122, 
    570.6113482, 635.806353, 694.8286462, 747.1992533, 793.0044191, 
    832.5750255, 866.4443202, 895.1917865, 919.4060705, 939.6860264, 
    956.4664631, 970.1833931, 981.1347983, 989.68, 995.9, 1000 ;

 grid_lon =
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125,
  35, 35.78278, 36.57269, 37.36979, 38.17411, 38.98572, 39.80465, 40.63093, 
    41.46459, 42.30565, 43.15412, 44.01001, 44.87331, 45.744, 46.62207, 
    47.50749, 48.40021, 49.30018, 50.20734, 51.12163, 52.04295, 52.97122, 
    53.90633, 54.84815, 55.79657, 56.75144, 57.71262, 58.67992, 59.65319, 
    60.63222, 61.61683, 62.60678, 63.60188, 64.60188, 65.60651, 66.61555, 
    67.62873, 68.64574, 69.66634, 70.69019, 71.71702, 72.7465, 73.77832, 
    74.81216, 75.84769, 76.88457, 77.92248, 78.96107, 80, 81.03893, 82.07752, 
    83.11543, 84.15231, 85.18784, 86.22168, 87.2535, 88.28298, 89.30981, 
    90.33366, 91.35426, 92.37127, 93.38445, 94.39349, 95.39812, 96.39812, 
    97.39321, 98.38318, 99.36778, 100.3468, 101.3201, 102.2874, 103.2486, 
    104.2034, 105.1518, 106.0937, 107.0288, 107.957, 108.8784, 109.7927, 
    110.6998, 111.5998, 112.4925, 113.3779, 114.256, 115.1267, 115.99, 
    116.8459, 117.6944, 118.5354, 119.3691, 120.1954, 121.0143, 121.8259, 
    122.6302, 123.4273, 124.2172, 125 ;

 grid_lat =
  -35.26439, -35.62921, -35.98892, -36.34341, -36.69255, -37.03624, 
    -37.37434, -37.70675, -38.03334, -38.354, -38.66859, -38.977, -39.27911, 
    -39.57478, -39.8639, -40.14635, -40.42199, -40.69072, -40.9524, 
    -41.20691, -41.45414, -41.69396, -41.92625, -42.15091, -42.36781, 
    -42.57683, -42.77788, -42.97084, -43.1556, -43.33206, -43.50012, 
    -43.65969, -43.81068, -43.95298, -44.08652, -44.21122, -44.32701, 
    -44.4338, -44.53154, -44.62016, -44.6996, -44.76982, -44.83077, 
    -44.88241, -44.9247, -44.95763, -44.98116, -44.99529, -45, -44.99529, 
    -44.98116, -44.95763, -44.9247, -44.88241, -44.83077, -44.76982, 
    -44.6996, -44.62016, -44.53154, -44.4338, -44.32701, -44.21122, 
    -44.08652, -43.95298, -43.81068, -43.65969, -43.50012, -43.33206, 
    -43.1556, -42.97084, -42.77788, -42.57683, -42.36781, -42.15091, 
    -41.92625, -41.69396, -41.45414, -41.20691, -40.9524, -40.69072, 
    -40.42199, -40.14635, -39.8639, -39.57478, -39.27911, -38.977, -38.66859, 
    -38.354, -38.03334, -37.70675, -37.37434, -37.03624, -36.69255, 
    -36.34341, -35.98892, -35.62921, -35.26439,
  -34.52972, -34.89117, -35.24767, -35.59911, -35.94537, -36.28631, 
    -36.62183, -36.95179, -37.27608, -37.59457, -37.90713, -38.21363, 
    -38.51395, -38.80796, -39.09554, -39.37654, -39.65086, -39.91835, 
    -40.1789, -40.43238, -40.67865, -40.9176, -41.14911, -41.37305, -41.5893, 
    -41.79774, -41.99827, -42.19077, -42.37512, -42.55122, -42.71897, 
    -42.87827, -43.02901, -43.17111, -43.30448, -43.42903, -43.54469, 
    -43.65138, -43.74903, -43.83758, -43.91697, -43.98714, -44.04806, 
    -44.09967, -44.14195, -44.17486, -44.19839, -44.21251, -44.21722, 
    -44.21251, -44.19839, -44.17486, -44.14195, -44.09967, -44.04806, 
    -43.98714, -43.91697, -43.83758, -43.74903, -43.65138, -43.54469, 
    -43.42903, -43.30448, -43.17111, -43.02901, -42.87827, -42.71897, 
    -42.55122, -42.37512, -42.19077, -41.99827, -41.79774, -41.5893, 
    -41.37305, -41.14911, -40.9176, -40.67865, -40.43238, -40.1789, 
    -39.91835, -39.65086, -39.37654, -39.09554, -38.80796, -38.51395, 
    -38.21363, -37.90713, -37.59457, -37.27608, -36.95179, -36.62183, 
    -36.28631, -35.94537, -35.59911, -35.24767, -34.89117, -34.52972,
  -33.79504, -34.15289, -34.50594, -34.8541, -35.19722, -35.53519, -35.86789, 
    -36.19517, -36.51693, -36.83301, -37.14331, -37.44768, -37.746, 
    -38.03813, -38.32394, -38.6033, -38.87608, -39.14214, -39.40136, 
    -39.6536, -39.89874, -40.13664, -40.36718, -40.59023, -40.80568, 
    -41.01338, -41.21324, -41.40512, -41.58892, -41.76453, -41.93184, 
    -42.09073, -42.24112, -42.38291, -42.516, -42.64032, -42.75576, 
    -42.86227, -42.95976, -43.04817, -43.12745, -43.19752, -43.25835, 
    -43.3099, -43.35213, -43.385, -43.4085, -43.4226, -43.42731, -43.4226, 
    -43.4085, -43.385, -43.35213, -43.3099, -43.25835, -43.19752, -43.12745, 
    -43.04817, -42.95976, -42.86227, -42.75576, -42.64032, -42.516, 
    -42.38291, -42.24112, -42.09073, -41.93184, -41.76453, -41.58892, 
    -41.40512, -41.21324, -41.01338, -40.80568, -40.59023, -40.36718, 
    -40.13664, -39.89874, -39.6536, -39.40136, -39.14214, -38.87608, 
    -38.6033, -38.32394, -38.03813, -37.746, -37.44768, -37.14331, -36.83301, 
    -36.51693, -36.19517, -35.86789, -35.53519, -35.19722, -34.8541, 
    -34.50594, -34.15289, -33.79504,
  -33.06036, -33.41436, -33.76374, -34.10837, -34.44813, -34.78289, 
    -35.11252, -35.4369, -35.75588, -36.06934, -36.37715, -36.67916, 
    -36.97525, -37.26529, -37.54912, -37.82662, -38.09766, -38.36209, 
    -38.61978, -38.87059, -39.1144, -39.35107, -39.58046, -39.80246, 
    -40.01692, -40.22372, -40.42275, -40.61388, -40.79699, -40.97196, 
    -41.13869, -41.29707, -41.44698, -41.58834, -41.72106, -41.84503, 
    -41.96017, -42.06641, -42.16367, -42.25187, -42.33097, -42.40089, 
    -42.4616, -42.51304, -42.55518, -42.58799, -42.61144, -42.62552, 
    -42.63021, -42.62552, -42.61144, -42.58799, -42.55518, -42.51304, 
    -42.4616, -42.40089, -42.33097, -42.25187, -42.16367, -42.06641, 
    -41.96017, -41.84503, -41.72106, -41.58834, -41.44698, -41.29707, 
    -41.13869, -40.97196, -40.79699, -40.61388, -40.42275, -40.22372, 
    -40.01692, -39.80246, -39.58046, -39.35107, -39.1144, -38.87059, 
    -38.61978, -38.36209, -38.09766, -37.82662, -37.54912, -37.26529, 
    -36.97525, -36.67916, -36.37715, -36.06934, -35.75588, -35.4369, 
    -35.11252, -34.78289, -34.44813, -34.10837, -33.76374, -33.41436, 
    -33.06036,
  -32.32569, -32.67561, -33.02107, -33.36194, -33.6981, -34.02942, -34.35575, 
    -34.67698, -34.99296, -35.30357, -35.60866, -35.90809, -36.20173, 
    -36.48944, -36.77109, -37.04652, -37.3156, -37.57819, -37.83415, 
    -38.08334, -38.32563, -38.56088, -38.78895, -39.00971, -39.22302, 
    -39.42876, -39.6268, -39.81702, -39.99928, -40.17348, -40.3395, 
    -40.49723, -40.64656, -40.78738, -40.91961, -41.04314, -41.15789, 
    -41.26377, -41.36071, -41.44865, -41.5275, -41.59722, -41.65775, 
    -41.70904, -41.75106, -41.78378, -41.80717, -41.82121, -41.82589, 
    -41.82121, -41.80717, -41.78378, -41.75106, -41.70904, -41.65775, 
    -41.59722, -41.5275, -41.44865, -41.36071, -41.26377, -41.15789, 
    -41.04314, -40.91961, -40.78738, -40.64656, -40.49723, -40.3395, 
    -40.17348, -39.99928, -39.81702, -39.6268, -39.42876, -39.22302, 
    -39.00971, -38.78895, -38.56088, -38.32563, -38.08334, -37.83415, 
    -37.57819, -37.3156, -37.04652, -36.77109, -36.48944, -36.20173, 
    -35.90809, -35.60866, -35.30357, -34.99296, -34.67698, -34.35575, 
    -34.02942, -33.6981, -33.36194, -33.02107, -32.67561, -32.32569,
  -31.59101, -31.93662, -32.27793, -32.61481, -32.94714, -33.27477, 
    -33.59758, -33.91543, -34.22818, -34.5357, -34.83784, -35.13448, 
    -35.42545, -35.71062, -35.98985, -36.26299, -36.52991, -36.79046, 
    -37.04449, -37.29186, -37.53244, -37.76608, -37.99264, -38.21198, 
    -38.42397, -38.62848, -38.82537, -39.01452, -39.1958, -39.36908, 
    -39.53426, -39.69121, -39.83982, -39.97999, -40.11162, -40.23461, 
    -40.34887, -40.45432, -40.55087, -40.63845, -40.717, -40.78645, 
    -40.84675, -40.89785, -40.93972, -40.97232, -40.99562, -41.00961, 
    -41.01428, -41.00961, -40.99562, -40.97232, -40.93972, -40.89785, 
    -40.84675, -40.78645, -40.717, -40.63845, -40.55087, -40.45432, 
    -40.34887, -40.23461, -40.11162, -39.97999, -39.83982, -39.69121, 
    -39.53426, -39.36908, -39.1958, -39.01452, -38.82537, -38.62848, 
    -38.42397, -38.21198, -37.99264, -37.76608, -37.53244, -37.29186, 
    -37.04449, -36.79046, -36.52991, -36.26299, -35.98985, -35.71062, 
    -35.42545, -35.13448, -34.83784, -34.5357, -34.22818, -33.91543, 
    -33.59758, -33.27477, -32.94714, -32.61481, -32.27793, -31.93662, 
    -31.59101,
  -30.85634, -31.19741, -31.53433, -31.86699, -32.19525, -32.51897, 
    -32.83802, -33.15226, -33.46156, -33.76576, -34.06473, -34.35833, 
    -34.64641, -34.92882, -35.20542, -35.47607, -35.74061, -35.9989, 
    -36.2508, -36.49615, -36.73482, -36.96666, -37.19153, -37.40928, 
    -37.61977, -37.82288, -38.01846, -38.20639, -38.38652, -38.55875, 
    -38.72294, -38.87898, -39.02676, -39.16616, -39.29708, -39.41943, 
    -39.5331, -39.63801, -39.73409, -39.82125, -39.89942, -39.96855, 
    -40.02857, -40.07944, -40.12112, -40.15358, -40.17678, -40.1907, 
    -40.19535, -40.1907, -40.17678, -40.15358, -40.12112, -40.07944, 
    -40.02857, -39.96855, -39.89942, -39.82125, -39.73409, -39.63801, 
    -39.5331, -39.41943, -39.29708, -39.16616, -39.02676, -38.87898, 
    -38.72294, -38.55875, -38.38652, -38.20639, -38.01846, -37.82288, 
    -37.61977, -37.40928, -37.19153, -36.96666, -36.73482, -36.49615, 
    -36.2508, -35.9989, -35.74061, -35.47607, -35.20542, -34.92882, 
    -34.64641, -34.35833, -34.06473, -33.76576, -33.46156, -33.15226, 
    -32.83802, -32.51897, -32.19525, -31.86699, -31.53433, -31.19741, 
    -30.85634,
  -30.12167, -30.45796, -30.79028, -31.11849, -31.44245, -31.76203, -32.0771, 
    -32.3875, -32.6931, -32.99376, -33.28933, -33.57967, -33.86464, 
    -34.14407, -34.41782, -34.68575, -34.94771, -35.20354, -35.45309, 
    -35.69623, -35.9328, -36.16264, -36.38563, -36.6016, -36.81043, 
    -37.01196, -37.20607, -37.39261, -37.57145, -37.74247, -37.90554, 
    -38.06054, -38.20735, -38.34586, -38.47596, -38.59755, -38.71054, 
    -38.81484, -38.91036, -38.99702, -39.07475, -39.1435, -39.20319, 
    -39.25378, -39.29524, -39.32752, -39.3506, -39.36445, -39.36907, 
    -39.36445, -39.3506, -39.32752, -39.29524, -39.25378, -39.20319, 
    -39.1435, -39.07475, -38.99702, -38.91036, -38.81484, -38.71054, 
    -38.59755, -38.47596, -38.34586, -38.20735, -38.06054, -37.90554, 
    -37.74247, -37.57145, -37.39261, -37.20607, -37.01196, -36.81043, 
    -36.6016, -36.38563, -36.16264, -35.9328, -35.69623, -35.45309, 
    -35.20354, -34.94771, -34.68575, -34.41782, -34.14407, -33.86464, 
    -33.57967, -33.28933, -32.99376, -32.6931, -32.3875, -32.0771, -31.76203, 
    -31.44245, -31.11849, -30.79028, -30.45796, -30.12167,
  -29.38699, -29.7183, -30.04578, -30.36931, -30.68875, -31.00396, -31.31481, 
    -31.62114, -31.92283, -32.21972, -32.51167, -32.79853, -33.08015, 
    -33.35638, -33.62707, -33.89207, -34.15122, -34.40438, -34.6514, 
    -34.89211, -35.12637, -35.35404, -35.57495, -35.78897, -35.99594, 
    -36.19573, -36.38819, -36.57319, -36.75058, -36.92025, -37.08205, 
    -37.23587, -37.38158, -37.51908, -37.64825, -37.76899, -37.8812, 
    -37.98478, -38.07965, -38.16574, -38.24297, -38.31126, -38.37057, 
    -38.42085, -38.46204, -38.49412, -38.51705, -38.53082, -38.53541, 
    -38.53082, -38.51705, -38.49412, -38.46204, -38.42085, -38.37057, 
    -38.31126, -38.24297, -38.16574, -38.07965, -37.98478, -37.8812, 
    -37.76899, -37.64825, -37.51908, -37.38158, -37.23587, -37.08205, 
    -36.92025, -36.75058, -36.57319, -36.38819, -36.19573, -35.99594, 
    -35.78897, -35.57495, -35.35404, -35.12637, -34.89211, -34.6514, 
    -34.40438, -34.15122, -33.89207, -33.62707, -33.35638, -33.08015, 
    -32.79853, -32.51167, -32.21972, -31.92283, -31.62114, -31.31481, 
    -31.00396, -30.68875, -30.36931, -30.04578, -29.7183, -29.38699,
  -28.65232, -28.97841, -29.30084, -29.61947, -29.93416, -30.24478, 
    -30.55118, -30.85322, -31.15076, -31.44366, -31.73176, -32.01491, 
    -32.29297, -32.56578, -32.83318, -33.09504, -33.35118, -33.60146, 
    -33.84572, -34.08381, -34.31557, -34.54086, -34.75951, -34.97139, 
    -35.17633, -35.3742, -35.56485, -35.74813, -35.92393, -36.09208, 
    -36.25248, -36.40498, -36.54947, -36.68583, -36.81395, -36.93372, 
    -37.04504, -37.14782, -37.24197, -37.3274, -37.40405, -37.47184, 
    -37.53071, -37.58062, -37.62151, -37.65335, -37.67612, -37.68979, 
    -37.69435, -37.68979, -37.67612, -37.65335, -37.62151, -37.58062, 
    -37.53071, -37.47184, -37.40405, -37.3274, -37.24197, -37.14782, 
    -37.04504, -36.93372, -36.81395, -36.68583, -36.54947, -36.40498, 
    -36.25248, -36.09208, -35.92393, -35.74813, -35.56485, -35.3742, 
    -35.17633, -34.97139, -34.75951, -34.54086, -34.31557, -34.08381, 
    -33.84572, -33.60146, -33.35118, -33.09504, -32.83318, -32.56578, 
    -32.29297, -32.01491, -31.73176, -31.44366, -31.15076, -30.85322, 
    -30.55118, -30.24478, -29.93416, -29.61947, -29.30084, -28.97841, 
    -28.65232,
  -27.91764, -28.23831, -28.55546, -28.86897, -29.17869, -29.48449, 
    -29.78622, -30.08375, -30.37692, -30.6656, -30.94962, -31.22885, 
    -31.50312, -31.77229, -32.03619, -32.29469, -32.5476, -32.79479, 
    -33.03609, -33.27135, -33.50042, -33.72313, -33.93933, -34.14888, 
    -34.35161, -34.54738, -34.73605, -34.91746, -35.09149, -35.25799, 
    -35.41682, -35.56787, -35.71101, -35.8461, -35.97306, -36.09175, 
    -36.20208, -36.30396, -36.39729, -36.48199, -36.55799, -36.62521, 
    -36.68359, -36.73308, -36.77364, -36.80522, -36.8278, -36.84136, 
    -36.84588, -36.84136, -36.8278, -36.80522, -36.77364, -36.73308, 
    -36.68359, -36.62521, -36.55799, -36.48199, -36.39729, -36.30396, 
    -36.20208, -36.09175, -35.97306, -35.8461, -35.71101, -35.56787, 
    -35.41682, -35.25799, -35.09149, -34.91746, -34.73605, -34.54738, 
    -34.35161, -34.14888, -33.93933, -33.72313, -33.50042, -33.27135, 
    -33.03609, -32.79479, -32.5476, -32.29469, -32.03619, -31.77229, 
    -31.50312, -31.22885, -30.94962, -30.6656, -30.37692, -30.08375, 
    -29.78622, -29.48449, -29.17869, -28.86897, -28.55546, -28.23831, 
    -27.91764,
  -27.18297, -27.49799, -27.80966, -28.11782, -28.42235, -28.72311, 
    -29.01996, -29.31275, -29.60133, -29.88556, -30.16529, -30.44036, 
    -30.71063, -30.97594, -31.23613, -31.49104, -31.74052, -31.98441, 
    -32.22254, -32.45477, -32.68093, -32.90088, -33.11443, -33.32146, 
    -33.5218, -33.7153, -33.90181, -34.08119, -34.25329, -34.41798, 
    -34.57511, -34.72456, -34.8662, -34.99992, -35.12558, -35.24308, 
    -35.35233, -35.45321, -35.54563, -35.62952, -35.70479, -35.77137, 
    -35.8292, -35.87823, -35.91842, -35.94971, -35.97208, -35.98551, 
    -35.98999, -35.98551, -35.97208, -35.94971, -35.91842, -35.87823, 
    -35.8292, -35.77137, -35.70479, -35.62952, -35.54563, -35.45321, 
    -35.35233, -35.24308, -35.12558, -34.99992, -34.8662, -34.72456, 
    -34.57511, -34.41798, -34.25329, -34.08119, -33.90181, -33.7153, 
    -33.5218, -33.32146, -33.11443, -32.90088, -32.68093, -32.45477, 
    -32.22254, -31.98441, -31.74052, -31.49104, -31.23613, -30.97594, 
    -30.71063, -30.44036, -30.16529, -29.88556, -29.60133, -29.31275, 
    -29.01996, -28.72311, -28.42235, -28.11782, -27.80966, -27.49799, 
    -27.18297,
  -26.44829, -26.75747, -27.06343, -27.36604, -27.66517, -27.96067, 
    -28.25241, -28.54023, -28.82401, -29.10357, -29.37879, -29.64949, 
    -29.91554, -30.17676, -30.43301, -30.68413, -30.92996, -31.17034, 
    -31.4051, -31.63409, -31.85715, -32.07413, -32.28485, -32.48917, 
    -32.68693, -32.87798, -33.06216, -33.23934, -33.40936, -33.57207, 
    -33.72735, -33.87507, -34.01508, -34.14728, -34.27153, -34.38773, 
    -34.49578, -34.59556, -34.68699, -34.76999, -34.84446, -34.91034, 
    -34.96757, -35.01609, -35.05586, -35.08683, -35.10897, -35.12226, 
    -35.12669, -35.12226, -35.10897, -35.08683, -35.05586, -35.01609, 
    -34.96757, -34.91034, -34.84446, -34.76999, -34.68699, -34.59556, 
    -34.49578, -34.38773, -34.27153, -34.14728, -34.01508, -33.87507, 
    -33.72735, -33.57207, -33.40936, -33.23934, -33.06216, -32.87798, 
    -32.68693, -32.48917, -32.28485, -32.07413, -31.85715, -31.63409, 
    -31.4051, -31.17034, -30.92996, -30.68413, -30.43301, -30.17676, 
    -29.91554, -29.64949, -29.37879, -29.10357, -28.82401, -28.54023, 
    -28.25241, -27.96067, -27.66517, -27.36604, -27.06343, -26.75747, 
    -26.44829,
  -25.71362, -26.01674, -26.31679, -26.61363, -26.90714, -27.19717, 
    -27.48358, -27.76624, -28.04498, -28.31966, -28.59014, -28.85626, 
    -29.11786, -29.37479, -29.62689, -29.874, -30.11596, -30.35262, -30.5838, 
    -30.80936, -31.02912, -31.24292, -31.45062, -31.65205, -31.84704, 
    -32.03546, -32.21714, -32.39194, -32.55971, -32.7203, -32.87358, 
    -33.01942, -33.15767, -33.28822, -33.41094, -33.52573, -33.63246, 
    -33.73105, -33.8214, -33.90341, -33.97701, -34.04213, -34.0987, 
    -34.14666, -34.18597, -34.21658, -34.23848, -34.25162, -34.256, 
    -34.25162, -34.23848, -34.21658, -34.18597, -34.14666, -34.0987, 
    -34.04213, -33.97701, -33.90341, -33.8214, -33.73105, -33.63246, 
    -33.52573, -33.41094, -33.28822, -33.15767, -33.01942, -32.87358, 
    -32.7203, -32.55971, -32.39194, -32.21714, -32.03546, -31.84704, 
    -31.65205, -31.45062, -31.24292, -31.02912, -30.80936, -30.5838, 
    -30.35262, -30.11596, -29.874, -29.62689, -29.37479, -29.11786, 
    -28.85626, -28.59014, -28.31966, -28.04498, -27.76624, -27.48358, 
    -27.19717, -26.90714, -26.61363, -26.31679, -26.01674, -25.71362,
  -24.97894, -25.2758, -25.56974, -25.86061, -26.14829, -26.43264, -26.71351, 
    -26.99077, -27.26427, -27.53386, -27.79938, -28.0607, -28.31764, 
    -28.57006, -28.81779, -29.06068, -29.29857, -29.5313, -29.75869, 
    -29.9806, -30.19686, -30.4073, -30.61178, -30.81012, -31.00217, 
    -31.18778, -31.36679, -31.53904, -31.7044, -31.86271, -32.01384, 
    -32.15764, -32.29399, -32.42276, -32.54383, -32.65709, -32.76241, 
    -32.85971, -32.94887, -33.02983, -33.10248, -33.16676, -33.22261, 
    -33.26997, -33.30878, -33.33901, -33.36062, -33.3736, -33.37793, 
    -33.3736, -33.36062, -33.33901, -33.30878, -33.26997, -33.22261, 
    -33.16676, -33.10248, -33.02983, -32.94887, -32.85971, -32.76241, 
    -32.65709, -32.54383, -32.42276, -32.29399, -32.15764, -32.01384, 
    -31.86271, -31.7044, -31.53904, -31.36679, -31.18778, -31.00217, 
    -30.81012, -30.61178, -30.4073, -30.19686, -29.9806, -29.75869, -29.5313, 
    -29.29857, -29.06068, -28.81779, -28.57006, -28.31764, -28.0607, 
    -27.79938, -27.53386, -27.26427, -26.99077, -26.71351, -26.43264, 
    -26.14829, -25.86061, -25.56974, -25.2758, -24.97894,
  -24.24427, -24.53467, -24.82229, -25.10699, -25.38863, -25.66709, 
    -25.94222, -26.21387, -26.48191, -26.74619, -27.00655, -27.26284, 
    -27.51491, -27.76261, -28.00576, -28.24422, -28.47782, -28.70641, 
    -28.92981, -29.14787, -29.36043, -29.56732, -29.76838, -29.96344, 
    -30.15236, -30.33498, -30.51114, -30.68068, -30.84346, -30.99933, 
    -31.14815, -31.28979, -31.4241, -31.55096, -31.67025, -31.78186, 
    -31.88566, -31.98156, -32.06945, -32.14926, -32.22089, -32.28428, 
    -32.33934, -32.38604, -32.42432, -32.45413, -32.47544, -32.48825, 
    -32.49251, -32.48825, -32.47544, -32.45413, -32.42432, -32.38604, 
    -32.33934, -32.28428, -32.22089, -32.14926, -32.06945, -31.98156, 
    -31.88566, -31.78186, -31.67025, -31.55096, -31.4241, -31.28979, 
    -31.14815, -30.99933, -30.84346, -30.68068, -30.51114, -30.33498, 
    -30.15236, -29.96344, -29.76838, -29.56732, -29.36043, -29.14787, 
    -28.92981, -28.70641, -28.47782, -28.24422, -28.00576, -27.76261, 
    -27.51491, -27.26284, -27.00655, -26.74619, -26.48191, -26.21387, 
    -25.94222, -25.66709, -25.38863, -25.10699, -24.82229, -24.53467, 
    -24.24427,
  -23.50959, -23.79335, -24.07445, -24.35277, -24.62818, -24.90054, 
    -25.16972, -25.43556, -25.69794, -25.95669, -26.21167, -26.46273, 
    -26.70972, -26.95247, -27.19084, -27.42466, -27.65377, -27.87801, 
    -28.09721, -28.31122, -28.51988, -28.72301, -28.92046, -29.11207, 
    -29.29767, -29.47712, -29.65025, -29.8169, -29.97694, -30.13022, 
    -30.27658, -30.4159, -30.54803, -30.67286, -30.79025, -30.90008, 
    -31.00225, -31.09665, -31.18319, -31.26176, -31.33229, -31.39471, 
    -31.44894, -31.49493, -31.53263, -31.56199, -31.58298, -31.59559, 
    -31.59979, -31.59559, -31.58298, -31.56199, -31.53263, -31.49493, 
    -31.44894, -31.39471, -31.33229, -31.26176, -31.18319, -31.09665, 
    -31.00225, -30.90008, -30.79025, -30.67286, -30.54803, -30.4159, 
    -30.27658, -30.13022, -29.97694, -29.8169, -29.65025, -29.47712, 
    -29.29767, -29.11207, -28.92046, -28.72301, -28.51988, -28.31122, 
    -28.09721, -27.87801, -27.65377, -27.42466, -27.19084, -26.95247, 
    -26.70972, -26.46273, -26.21167, -25.95669, -25.69794, -25.43556, 
    -25.16972, -24.90054, -24.62818, -24.35277, -24.07445, -23.79335, 
    -23.50959,
  -22.77492, -23.05183, -23.32623, -23.59798, -23.86696, -24.13302, 
    -24.39604, -24.65587, -24.91236, -25.16539, -25.41478, -25.6604, 
    -25.9021, -26.13971, -26.37307, -26.60204, -26.82645, -27.04614, 
    -27.26094, -27.47071, -27.67526, -27.87444, -28.06809, -28.25605, 
    -28.43815, -28.61425, -28.78417, -28.94778, -29.10491, -29.25543, 
    -29.39919, -29.53604, -29.66586, -29.78851, -29.90387, -30.01182, 
    -30.11224, -30.20505, -30.29012, -30.36738, -30.43673, -30.49811, 
    -30.55145, -30.59668, -30.63375, -30.66263, -30.68328, -30.69568, 
    -30.69982, -30.69568, -30.68328, -30.66263, -30.63375, -30.59668, 
    -30.55145, -30.49811, -30.43673, -30.36738, -30.29012, -30.20505, 
    -30.11224, -30.01182, -29.90387, -29.78851, -29.66586, -29.53604, 
    -29.39919, -29.25543, -29.10491, -28.94778, -28.78417, -28.61425, 
    -28.43815, -28.25605, -28.06809, -27.87444, -27.67526, -27.47071, 
    -27.26094, -27.04614, -26.82645, -26.60204, -26.37307, -26.13971, 
    -25.9021, -25.6604, -25.41478, -25.16539, -24.91236, -24.65587, 
    -24.39604, -24.13302, -23.86696, -23.59798, -23.32623, -23.05183, 
    -22.77492,
  -22.04024, -22.31014, -22.57764, -22.84263, -23.10497, -23.36455, -23.6212, 
    -23.87482, -24.12524, -24.37232, -24.61593, -24.85591, -25.0921, 
    -25.32435, -25.55252, -25.77643, -25.99593, -26.21087, -26.42107, 
    -26.62638, -26.82663, -27.02167, -27.21133, -27.39545, -27.57387, 
    -27.74643, -27.91298, -28.07337, -28.22743, -28.37503, -28.51603, 
    -28.65027, -28.77763, -28.89797, -29.01118, -29.11712, -29.2157, 
    -29.3068, -29.39032, -29.46618, -29.53428, -29.59455, -29.64693, 
    -29.69135, -29.72776, -29.75613, -29.77641, -29.78859, -29.79265, 
    -29.78859, -29.77641, -29.75613, -29.72776, -29.69135, -29.64693, 
    -29.59455, -29.53428, -29.46618, -29.39032, -29.3068, -29.2157, 
    -29.11712, -29.01118, -28.89797, -28.77763, -28.65027, -28.51603, 
    -28.37503, -28.22743, -28.07337, -27.91298, -27.74643, -27.57387, 
    -27.39545, -27.21133, -27.02167, -26.82663, -26.62638, -26.42107, 
    -26.21087, -25.99593, -25.77643, -25.55252, -25.32435, -25.0921, 
    -24.85591, -24.61593, -24.37232, -24.12524, -23.87482, -23.6212, 
    -23.36455, -23.10497, -22.84263, -22.57764, -22.31014, -22.04024,
  -21.30557, -21.56826, -21.82868, -22.08672, -22.34225, -22.59513, 
    -22.84524, -23.09244, -23.33659, -23.57754, -23.81515, -24.04927, 
    -24.27976, -24.50646, -24.72922, -24.94787, -25.16227, -25.37224, 
    -25.57764, -25.77831, -25.97407, -26.16477, -26.35024, -26.53034, 
    -26.70489, -26.87375, -27.03675, -27.19374, -27.34457, -27.4891, 
    -27.62718, -27.75867, -27.88343, -28.00133, -28.11226, -28.21608, 
    -28.3127, -28.40199, -28.48387, -28.55823, -28.625, -28.6841, -28.73546, 
    -28.77902, -28.81473, -28.84255, -28.86244, -28.87439, -28.87837, 
    -28.87439, -28.86244, -28.84255, -28.81473, -28.77902, -28.73546, 
    -28.6841, -28.625, -28.55823, -28.48387, -28.40199, -28.3127, -28.21608, 
    -28.11226, -28.00133, -27.88343, -27.75867, -27.62718, -27.4891, 
    -27.34457, -27.19374, -27.03675, -26.87375, -26.70489, -26.53034, 
    -26.35024, -26.16477, -25.97407, -25.77831, -25.57764, -25.37224, 
    -25.16227, -24.94787, -24.72922, -24.50646, -24.27976, -24.04927, 
    -23.81515, -23.57754, -23.33659, -23.09244, -22.84524, -22.59513, 
    -22.34225, -22.08672, -21.82868, -21.56826, -21.30557,
  -20.57089, -20.8262, -21.07937, -21.33028, -21.5788, -21.82482, -22.06818, 
    -22.30877, -22.54645, -22.78106, -23.01249, -23.24056, -23.46515, 
    -23.68609, -23.90323, -24.11643, -24.32551, -24.53034, -24.73074, 
    -24.92656, -25.11763, -25.3038, -25.48491, -25.6608, -25.8313, -25.99627, 
    -26.15555, -26.30898, -26.45642, -26.59771, -26.73272, -26.86131, 
    -26.98333, -27.09867, -27.20719, -27.30877, -27.40331, -27.4907, 
    -27.57083, -27.64362, -27.70898, -27.76684, -27.81712, -27.85977, 
    -27.89473, -27.92197, -27.94145, -27.95315, -27.95705, -27.95315, 
    -27.94145, -27.92197, -27.89473, -27.85977, -27.81712, -27.76684, 
    -27.70898, -27.64362, -27.57083, -27.4907, -27.40331, -27.30877, 
    -27.20719, -27.09867, -26.98333, -26.86131, -26.73272, -26.59771, 
    -26.45642, -26.30898, -26.15555, -25.99627, -25.8313, -25.6608, 
    -25.48491, -25.3038, -25.11763, -24.92656, -24.73074, -24.53034, 
    -24.32551, -24.11643, -23.90323, -23.68609, -23.46515, -23.24056, 
    -23.01249, -22.78106, -22.54645, -22.30877, -22.06818, -21.82482, 
    -21.5788, -21.33028, -21.07937, -20.8262, -20.57089,
  -19.83622, -20.08398, -20.32972, -20.57332, -20.81466, -21.05361, 
    -21.29005, -21.52384, -21.75485, -21.98295, -22.20798, -22.42981, 
    -22.6483, -22.86328, -23.07462, -23.28216, -23.48574, -23.68522, 
    -23.88042, -24.0712, -24.2574, -24.43885, -24.6154, -24.7869, -24.95318, 
    -25.11408, -25.26947, -25.41917, -25.56305, -25.70096, -25.83275, 
    -25.95829, -26.07744, -26.19007, -26.29606, -26.39529, -26.48764, 
    -26.57302, -26.65132, -26.72244, -26.78632, -26.84286, -26.892, 
    -26.93369, -26.96786, -26.99449, -27.01353, -27.02497, -27.02878, 
    -27.02497, -27.01353, -26.99449, -26.96786, -26.93369, -26.892, 
    -26.84286, -26.78632, -26.72244, -26.65132, -26.57302, -26.48764, 
    -26.39529, -26.29606, -26.19007, -26.07744, -25.95829, -25.83275, 
    -25.70096, -25.56305, -25.41917, -25.26947, -25.11408, -24.95318, 
    -24.7869, -24.6154, -24.43885, -24.2574, -24.0712, -23.88042, -23.68522, 
    -23.48574, -23.28216, -23.07462, -22.86328, -22.6483, -22.42981, 
    -22.20798, -21.98295, -21.75485, -21.52384, -21.29005, -21.05361, 
    -20.81466, -20.57332, -20.32972, -20.08398, -19.83622,
  -19.10155, -19.34159, -19.57973, -19.81585, -20.04982, -20.28154, 
    -20.51087, -20.73768, -20.96184, -21.18322, -21.40168, -21.61708, 
    -21.82927, -22.03811, -22.24345, -22.44514, -22.64302, -22.83695, 
    -23.02677, -23.21232, -23.39345, -23.57, -23.74181, -23.90874, -24.07061, 
    -24.22728, -24.3786, -24.52441, -24.66457, -24.79893, -24.92736, 
    -25.0497, -25.16584, -25.27564, -25.37897, -25.47573, -25.56579, 
    -25.64905, -25.72542, -25.7948, -25.85711, -25.91227, -25.96022, 
    -26.00089, -26.03424, -26.06021, -26.0788, -26.08995, -26.09367, 
    -26.08995, -26.0788, -26.06021, -26.03424, -26.00089, -25.96022, 
    -25.91227, -25.85711, -25.7948, -25.72542, -25.64905, -25.56579, 
    -25.47573, -25.37897, -25.27564, -25.16584, -25.0497, -24.92736, 
    -24.79893, -24.66457, -24.52441, -24.3786, -24.22728, -24.07061, 
    -23.90874, -23.74181, -23.57, -23.39345, -23.21232, -23.02677, -22.83695, 
    -22.64302, -22.44514, -22.24345, -22.03811, -21.82927, -21.61708, 
    -21.40168, -21.18322, -20.96184, -20.73768, -20.51087, -20.28154, 
    -20.04982, -19.81585, -19.57973, -19.34159, -19.10155,
  -18.36687, -18.59904, -18.82941, -19.05788, -19.28433, -19.50863, 
    -19.73068, -19.95033, -20.16746, -20.38194, -20.59364, -20.80241, 
    -21.00812, -21.21062, -21.40977, -21.60542, -21.79742, -21.98561, 
    -22.16986, -22.35, -22.52588, -22.69734, -22.86423, -23.0264, -23.18369, 
    -23.33596, -23.48304, -23.6248, -23.76108, -23.89175, -24.01665, 
    -24.13567, -24.24865, -24.35549, -24.45604, -24.55021, -24.63787, 
    -24.71892, -24.79326, -24.86081, -24.92148, -24.97519, -25.02188, 
    -25.06149, -25.09396, -25.11926, -25.13736, -25.14822, -25.15185, 
    -25.14822, -25.13736, -25.11926, -25.09396, -25.06149, -25.02188, 
    -24.97519, -24.92148, -24.86081, -24.79326, -24.71892, -24.63787, 
    -24.55021, -24.45604, -24.35549, -24.24865, -24.13567, -24.01665, 
    -23.89175, -23.76108, -23.6248, -23.48304, -23.33596, -23.18369, 
    -23.0264, -22.86423, -22.69734, -22.52588, -22.35, -22.16986, -21.98561, 
    -21.79742, -21.60542, -21.40977, -21.21062, -21.00812, -20.80241, 
    -20.59364, -20.38194, -20.16746, -19.95033, -19.73068, -19.50863, 
    -19.28433, -19.05788, -18.82941, -18.59904, -18.36687,
  -17.63219, -17.85633, -18.07879, -18.29944, -18.51819, -18.73492, -18.9495, 
    -19.16182, -19.37174, -19.57915, -19.7839, -19.98587, -20.18491, 
    -20.38089, -20.57367, -20.76309, -20.94901, -21.13129, -21.30978, 
    -21.48432, -21.65476, -21.82095, -21.98275, -22.13999, -22.29253, 
    -22.44022, -22.5829, -22.72045, -22.85269, -22.97951, -23.10075, 
    -23.21629, -23.32599, -23.42973, -23.52739, -23.61885, -23.704, 
    -23.78273, -23.85496, -23.92059, -23.97954, -24.03174, -24.07711, 
    -24.1156, -24.14717, -24.17175, -24.18934, -24.19991, -24.20343, 
    -24.19991, -24.18934, -24.17175, -24.14717, -24.1156, -24.07711, 
    -24.03174, -23.97954, -23.92059, -23.85496, -23.78273, -23.704, 
    -23.61885, -23.52739, -23.42973, -23.32599, -23.21629, -23.10075, 
    -22.97951, -22.85269, -22.72045, -22.5829, -22.44022, -22.29253, 
    -22.13999, -21.98275, -21.82095, -21.65476, -21.48432, -21.30978, 
    -21.13129, -20.94901, -20.76309, -20.57367, -20.38089, -20.18491, 
    -19.98587, -19.7839, -19.57915, -19.37174, -19.16182, -18.9495, 
    -18.73492, -18.51819, -18.29944, -18.07879, -17.85633, -17.63219,
  -16.89752, -17.11348, -17.32786, -17.54054, -17.75143, -17.96042, 
    -18.16737, -18.37219, -18.57473, -18.77489, -18.97252, -19.16751, 
    -19.35971, -19.54898, -19.7352, -19.91821, -20.09789, -20.27407, 
    -20.44661, -20.61537, -20.7802, -20.94095, -21.09747, -21.24961, 
    -21.39723, -21.54018, -21.6783, -21.81147, -21.93953, -22.06234, 
    -22.17978, -22.2917, -22.39799, -22.49851, -22.59314, -22.68178, 
    -22.76431, -22.84064, -22.91066, -22.97429, -23.03145, -23.08206, 
    -23.12605, -23.16338, -23.19399, -23.21784, -23.2349, -23.24514, 
    -23.24856, -23.24514, -23.2349, -23.21784, -23.19399, -23.16338, 
    -23.12605, -23.08206, -23.03145, -22.97429, -22.91066, -22.84064, 
    -22.76431, -22.68178, -22.59314, -22.49851, -22.39799, -22.2917, 
    -22.17978, -22.06234, -21.93953, -21.81147, -21.6783, -21.54018, 
    -21.39723, -21.24961, -21.09747, -20.94095, -20.7802, -20.61537, 
    -20.44661, -20.27407, -20.09789, -19.91821, -19.7352, -19.54898, 
    -19.35971, -19.16751, -18.97252, -18.77489, -18.57473, -18.37219, 
    -18.16737, -17.96042, -17.75143, -17.54054, -17.32786, -17.11348, 
    -16.89752,
  -16.16285, -16.37048, -16.57663, -16.7812, -16.98408, -17.18516, -17.38433, 
    -17.58147, -17.77647, -17.96921, -18.15956, -18.34738, -18.53256, 
    -18.71496, -18.89445, -19.07088, -19.24412, -19.41402, -19.58045, 
    -19.74325, -19.9023, -20.05743, -20.20851, -20.35538, -20.49791, 
    -20.63595, -20.76936, -20.89799, -21.02171, -21.14038, -21.25386, 
    -21.36204, -21.46477, -21.56195, -21.65344, -21.73915, -21.81896, 
    -21.89278, -21.9605, -22.02205, -22.07734, -22.1263, -22.16886, 
    -22.20498, -22.23459, -22.25766, -22.27417, -22.28408, -22.28739, 
    -22.28408, -22.27417, -22.25766, -22.23459, -22.20498, -22.16886, 
    -22.1263, -22.07734, -22.02205, -21.9605, -21.89278, -21.81896, 
    -21.73915, -21.65344, -21.56195, -21.46477, -21.36204, -21.25386, 
    -21.14038, -21.02171, -20.89799, -20.76936, -20.63595, -20.49791, 
    -20.35538, -20.20851, -20.05743, -19.9023, -19.74325, -19.58045, 
    -19.41402, -19.24412, -19.07088, -18.89445, -18.71496, -18.53256, 
    -18.34738, -18.15956, -17.96921, -17.77647, -17.58147, -17.38433, 
    -17.18516, -16.98408, -16.7812, -16.57663, -16.37048, -16.16285,
  -15.42817, -15.62734, -15.82513, -16.02143, -16.21614, -16.40917, -16.6004, 
    -16.78971, -16.97701, -17.16216, -17.34505, -17.52556, -17.70355, 
    -17.8789, -18.05148, -18.22116, -18.38779, -18.55125, -18.71139, 
    -18.86807, -19.02115, -19.1705, -19.31597, -19.45741, -19.59469, 
    -19.72766, -19.85619, -19.98014, -20.09937, -20.21375, -20.32315, 
    -20.42744, -20.5265, -20.6202, -20.70844, -20.79111, -20.8681, -20.9393, 
    -21.00464, -21.06402, -21.11737, -21.16462, -21.20569, -21.24054, 
    -21.26912, -21.29139, -21.30732, -21.31689, -21.32008, -21.31689, 
    -21.30732, -21.29139, -21.26912, -21.24054, -21.20569, -21.16462, 
    -21.11737, -21.06402, -21.00464, -20.9393, -20.8681, -20.79111, 
    -20.70844, -20.6202, -20.5265, -20.42744, -20.32315, -20.21375, 
    -20.09937, -19.98014, -19.85619, -19.72766, -19.59469, -19.45741, 
    -19.31597, -19.1705, -19.02115, -18.86807, -18.71139, -18.55125, 
    -18.38779, -18.22116, -18.05148, -17.8789, -17.70355, -17.52556, 
    -17.34505, -17.16216, -16.97701, -16.78971, -16.6004, -16.40917, 
    -16.21614, -16.02143, -15.82513, -15.62734, -15.42817,
  -14.6935, -14.88407, -15.07335, -15.26124, -15.44765, -15.63248, -15.81561, 
    -15.99695, -16.17639, -16.3538, -16.52908, -16.7021, -16.87274, 
    -17.04088, -17.20639, -17.36914, -17.52901, -17.68585, -17.83953, 
    -17.98992, -18.13688, -18.28028, -18.41997, -18.55582, -18.68769, 
    -18.81544, -18.93895, -19.05806, -19.17266, -19.28261, -19.38778, 
    -19.48806, -19.58331, -19.67343, -19.7583, -19.83782, -19.91188, 
    -19.98038, -20.04325, -20.10039, -20.15172, -20.19719, -20.23672, 
    -20.27026, -20.29777, -20.3192, -20.33454, -20.34374, -20.34682, 
    -20.34374, -20.33454, -20.3192, -20.29777, -20.27026, -20.23672, 
    -20.19719, -20.15172, -20.10039, -20.04325, -19.98038, -19.91188, 
    -19.83782, -19.7583, -19.67343, -19.58331, -19.48806, -19.38778, 
    -19.28261, -19.17266, -19.05806, -18.93895, -18.81544, -18.68769, 
    -18.55582, -18.41997, -18.28028, -18.13688, -17.98992, -17.83953, 
    -17.68585, -17.52901, -17.36914, -17.20639, -17.04088, -16.87274, 
    -16.7021, -16.52908, -16.3538, -16.17639, -15.99695, -15.81561, 
    -15.63248, -15.44765, -15.26124, -15.07335, -14.88407, -14.6935,
  -13.95882, -14.14067, -14.32132, -14.50067, -14.67863, -14.85512, 
    -15.03002, -15.20323, -15.37465, -15.54417, -15.71168, -15.87706, 
    -16.0402, -16.20097, -16.35925, -16.51492, -16.66785, -16.81791, 
    -16.96498, -17.10892, -17.2496, -17.38689, -17.52065, -17.65075, 
    -17.77705, -17.89944, -18.01776, -18.1319, -18.24172, -18.34711, 
    -18.44792, -18.54405, -18.63538, -18.7218, -18.80319, -18.87945, 
    -18.95048, -19.0162, -19.0765, -19.13132, -19.18058, -19.2242, -19.26213, 
    -19.29432, -19.32071, -19.34128, -19.356, -19.36483, -19.36778, 
    -19.36483, -19.356, -19.34128, -19.32071, -19.29432, -19.26213, -19.2242, 
    -19.18058, -19.13132, -19.0765, -19.0162, -18.95048, -18.87945, 
    -18.80319, -18.7218, -18.63538, -18.54405, -18.44792, -18.34711, 
    -18.24172, -18.1319, -18.01776, -17.89944, -17.77705, -17.65075, 
    -17.52065, -17.38689, -17.2496, -17.10892, -16.96498, -16.81791, 
    -16.66785, -16.51492, -16.35925, -16.20097, -16.0402, -15.87706, 
    -15.71168, -15.54417, -15.37465, -15.20323, -15.03002, -14.85512, 
    -14.67863, -14.50067, -14.32132, -14.14067, -13.95882,
  -13.22415, -13.39715, -13.56903, -13.73972, -13.90911, -14.07711, 
    -14.24364, -14.40859, -14.57185, -14.73334, -14.89293, -15.05052, 
    -15.20599, -15.35924, -15.51014, -15.65857, -15.80442, -15.94755, 
    -16.08784, -16.22518, -16.35942, -16.49044, -16.61812, -16.74232, 
    -16.86292, -16.97978, -17.09279, -17.20181, -17.30672, -17.4074, 
    -17.50373, -17.5956, -17.68288, -17.76548, -17.84328, -17.91618, 
    -17.9841, -18.04693, -18.1046, -18.15702, -18.20412, -18.24584, 
    -18.28212, -18.31291, -18.33815, -18.35783, -18.3719, -18.38036, 
    -18.38318, -18.38036, -18.3719, -18.35783, -18.33815, -18.31291, 
    -18.28212, -18.24584, -18.20412, -18.15702, -18.1046, -18.04693, 
    -17.9841, -17.91618, -17.84328, -17.76548, -17.68288, -17.5956, 
    -17.50373, -17.4074, -17.30672, -17.20181, -17.09279, -16.97978, 
    -16.86292, -16.74232, -16.61812, -16.49044, -16.35942, -16.22518, 
    -16.08784, -15.94755, -15.80442, -15.65857, -15.51014, -15.35924, 
    -15.20599, -15.05052, -14.89293, -14.73334, -14.57185, -14.40859, 
    -14.24364, -14.07711, -13.90911, -13.73972, -13.56903, -13.39715, 
    -13.22415,
  -12.48947, -12.65351, -12.81652, -12.97841, -13.1391, -13.2985, -13.45652, 
    -13.61306, -13.76804, -13.92135, -14.07288, -14.22254, -14.37021, 
    -14.51579, -14.65916, -14.8002, -14.93881, -15.07486, -15.20823, 
    -15.33881, -15.46647, -15.59108, -15.71253, -15.83068, -15.94542, 
    -16.05663, -16.16418, -16.26795, -16.36782, -16.46367, -16.55539, 
    -16.64287, -16.72599, -16.80466, -16.87877, -16.94822, -17.01292, 
    -17.07278, -17.12773, -17.17768, -17.22256, -17.26232, -17.2969, 
    -17.32624, -17.3503, -17.36906, -17.38247, -17.39053, -17.39322, 
    -17.39053, -17.38247, -17.36906, -17.3503, -17.32624, -17.2969, 
    -17.26232, -17.22256, -17.17768, -17.12773, -17.07278, -17.01292, 
    -16.94822, -16.87877, -16.80466, -16.72599, -16.64287, -16.55539, 
    -16.46367, -16.36782, -16.26795, -16.16418, -16.05663, -15.94542, 
    -15.83068, -15.71253, -15.59108, -15.46647, -15.33881, -15.20823, 
    -15.07486, -14.93881, -14.8002, -14.65916, -14.51579, -14.37021, 
    -14.22254, -14.07288, -13.92135, -13.76804, -13.61306, -13.45652, 
    -13.2985, -13.1391, -12.97841, -12.81652, -12.65351, -12.48947,
  -11.7548, -11.90976, -12.06378, -12.21676, -12.36863, -12.5193, -12.66869, 
    -12.81671, -12.96326, -13.10826, -13.2516, -13.39319, -13.53292, 
    -13.67069, -13.80638, -13.9399, -14.07113, -14.19996, -14.32627, 
    -14.44994, -14.57087, -14.68893, -14.804, -14.91598, -15.02473, 
    -15.13014, -15.2321, -15.33048, -15.42518, -15.51608, -15.60307, 
    -15.68605, -15.7649, -15.83954, -15.90985, -15.97575, -16.03714, 
    -16.09396, -16.1461, -16.19351, -16.23612, -16.27386, -16.30668, 
    -16.33454, -16.35738, -16.37519, -16.38792, -16.39557, -16.39812, 
    -16.39557, -16.38792, -16.37519, -16.35738, -16.33454, -16.30668, 
    -16.27386, -16.23612, -16.19351, -16.1461, -16.09396, -16.03714, 
    -15.97575, -15.90985, -15.83954, -15.7649, -15.68605, -15.60307, 
    -15.51608, -15.42518, -15.33048, -15.2321, -15.13014, -15.02473, 
    -14.91598, -14.804, -14.68893, -14.57087, -14.44994, -14.32627, 
    -14.19996, -14.07113, -13.9399, -13.80638, -13.67069, -13.53292, 
    -13.39319, -13.2516, -13.10826, -12.96326, -12.81671, -12.66869, 
    -12.5193, -12.36863, -12.21676, -12.06378, -11.90976, -11.7548,
  -11.02012, -11.16591, -11.31083, -11.45479, -11.59772, -11.73955, 
    -11.88019, -12.01956, -12.15757, -12.29414, -12.42916, -12.56255, 
    -12.6942, -12.82403, -12.95192, -13.07777, -13.20149, -13.32295, 
    -13.44206, -13.5587, -13.67276, -13.78413, -13.8927, -13.99836, 
    -14.10098, -14.20047, -14.29671, -14.38959, -14.479, -14.56483, 
    -14.64697, -14.72534, -14.79981, -14.87031, -14.93673, -14.99899, 
    -15.05699, -15.11067, -15.15995, -15.20475, -15.24501, -15.28068, 
    -15.3117, -15.33803, -15.35962, -15.37645, -15.38849, -15.39572, 
    -15.39813, -15.39572, -15.38849, -15.37645, -15.35962, -15.33803, 
    -15.3117, -15.28068, -15.24501, -15.20475, -15.15995, -15.11067, 
    -15.05699, -14.99899, -14.93673, -14.87031, -14.79981, -14.72534, 
    -14.64697, -14.56483, -14.479, -14.38959, -14.29671, -14.20047, 
    -14.10098, -13.99836, -13.8927, -13.78413, -13.67276, -13.5587, 
    -13.44206, -13.32295, -13.20149, -13.07777, -12.95192, -12.82403, 
    -12.6942, -12.56255, -12.42916, -12.29414, -12.15757, -12.01956, 
    -11.88019, -11.73955, -11.59772, -11.45479, -11.31083, -11.16591, 
    -11.02012,
  -10.28545, -10.42197, -10.55768, -10.69252, -10.82641, -10.95929, 
    -11.09107, -11.22167, -11.35102, -11.47903, -11.60561, -11.73068, 
    -11.85414, -11.97589, -12.09585, -12.21391, -12.32998, -12.44396, 
    -12.55573, -12.66521, -12.77227, -12.87683, -12.97877, -13.07798, 
    -13.17436, -13.2678, -13.3582, -13.44545, -13.52945, -13.61009, 
    -13.68729, -13.76093, -13.83093, -13.89719, -13.95963, -14.01815, 
    -14.07269, -14.12316, -14.16949, -14.21162, -14.24948, -14.28303, 
    -14.3122, -14.33696, -14.35726, -14.37309, -14.38441, -14.39121, 
    -14.39348, -14.39121, -14.38441, -14.37309, -14.35726, -14.33696, 
    -14.3122, -14.28303, -14.24948, -14.21162, -14.16949, -14.12316, 
    -14.07269, -14.01815, -13.95963, -13.89719, -13.83093, -13.76093, 
    -13.68729, -13.61009, -13.52945, -13.44545, -13.3582, -13.2678, 
    -13.17436, -13.07798, -12.97877, -12.87683, -12.77227, -12.66521, 
    -12.55573, -12.44396, -12.32998, -12.21391, -12.09585, -11.97589, 
    -11.85414, -11.73068, -11.60561, -11.47903, -11.35102, -11.22167, 
    -11.09107, -10.95929, -10.82641, -10.69252, -10.55768, -10.42197, 
    -10.28545,
  -9.550773, -9.677926, -9.804344, -9.929964, -10.05472, -10.17854, 
    -10.30135, -10.42309, -10.54366, -10.66301, -10.78103, -10.89766, 
    -11.0128, -11.12637, -11.23828, -11.34843, -11.45673, -11.5631, 
    -11.66742, -11.7696, -11.86955, -11.96717, -12.06235, -12.155, -12.24501, 
    -12.33229, -12.41673, -12.49824, -12.57673, -12.65208, -12.72422, 
    -12.79304, -12.85847, -12.9204, -12.97877, -13.03348, -13.08447, 
    -13.13165, -13.17497, -13.21437, -13.24977, -13.28114, -13.30842, 
    -13.33158, -13.35057, -13.36537, -13.37596, -13.38232, -13.38444, 
    -13.38232, -13.37596, -13.36537, -13.35057, -13.33158, -13.30842, 
    -13.28114, -13.24977, -13.21437, -13.17497, -13.13165, -13.08447, 
    -13.03348, -12.97877, -12.9204, -12.85847, -12.79304, -12.72422, 
    -12.65208, -12.57673, -12.49824, -12.41673, -12.33229, -12.24501, 
    -12.155, -12.06235, -11.96717, -11.86955, -11.7696, -11.66742, -11.5631, 
    -11.45673, -11.34843, -11.23828, -11.12637, -11.0128, -10.89766, 
    -10.78103, -10.66301, -10.54366, -10.42309, -10.30135, -10.17854, 
    -10.05472, -9.929964, -9.804344, -9.677926, -9.550773,
  -8.816097, -8.933801, -9.050837, -9.167146, -9.282667, -9.397336, 
    -9.511086, -9.623848, -9.735553, -9.846126, -9.955491, -10.06357, 
    -10.17029, -10.27556, -10.3793, -10.48143, -10.58185, -10.68048, 
    -10.77724, -10.87202, -10.96474, -11.0553, -11.14361, -11.22959, 
    -11.31312, -11.39412, -11.47251, -11.54817, -11.62103, -11.691, 
    -11.75798, -11.82189, -11.88264, -11.94017, -11.99438, -12.0452, 
    -12.09256, -12.1364, -12.17664, -12.21324, -12.24614, -12.27528, 
    -12.30063, -12.32215, -12.3398, -12.35355, -12.36339, -12.3693, 
    -12.37127, -12.3693, -12.36339, -12.35355, -12.3398, -12.32215, 
    -12.30063, -12.27528, -12.24614, -12.21324, -12.17664, -12.1364, 
    -12.09256, -12.0452, -11.99438, -11.94017, -11.88264, -11.82189, 
    -11.75798, -11.691, -11.62103, -11.54817, -11.47251, -11.39412, 
    -11.31312, -11.22959, -11.14361, -11.0553, -10.96474, -10.87202, 
    -10.77724, -10.68048, -10.58185, -10.48143, -10.3793, -10.27556, 
    -10.17029, -10.06357, -9.955491, -9.846126, -9.735553, -9.623848, 
    -9.511086, -9.397336, -9.282667, -9.167146, -9.050837, -8.933801, 
    -8.816097,
  -8.081423, -8.189597, -8.297169, -8.404083, -8.510284, -8.615713, 
    -8.720308, -8.824006, -8.926742, -9.028447, -9.129053, -9.228487, 
    -9.326677, -9.423547, -9.519018, -9.613013, -9.705451, -9.79625, 
    -9.885328, -9.972599, -10.05798, -10.14138, -10.22272, -10.30191, 
    -10.37886, -10.45349, -10.52571, -10.59543, -10.66257, -10.72705, 
    -10.78878, -10.84769, -10.90369, -10.95672, -11.0067, -11.05355, 
    -11.09722, -11.13764, -11.17476, -11.2085, -11.23884, -11.26572, 
    -11.2891, -11.30894, -11.32522, -11.33791, -11.34698, -11.35243, 
    -11.35425, -11.35243, -11.34698, -11.33791, -11.32522, -11.30894, 
    -11.2891, -11.26572, -11.23884, -11.2085, -11.17476, -11.13764, 
    -11.09722, -11.05355, -11.0067, -10.95672, -10.90369, -10.84769, 
    -10.78878, -10.72705, -10.66257, -10.59543, -10.52571, -10.45349, 
    -10.37886, -10.30191, -10.22272, -10.14138, -10.05798, -9.972599, 
    -9.885328, -9.79625, -9.705451, -9.613013, -9.519018, -9.423547, 
    -9.326677, -9.228487, -9.129053, -9.028447, -8.926742, -8.824006, 
    -8.720308, -8.615713, -8.510284, -8.404083, -8.297169, -8.189597, 
    -8.081423,
  -7.346748, -7.445321, -7.543353, -7.640796, -7.737598, -7.833705, 
    -7.929061, -8.023608, -8.117288, -8.210036, -8.30179, -8.392486, 
    -8.482054, -8.570426, -8.657532, -8.743299, -8.827652, -8.910519, 
    -8.99182, -9.071482, -9.149424, -9.225567, -9.299832, -9.372141, 
    -9.442413, -9.510569, -9.576528, -9.640213, -9.701547, -9.760451, 
    -9.816853, -9.870676, -9.92185, -9.970306, -10.01598, -10.0588, 
    -10.09871, -10.13566, -10.16958, -10.20043, -10.22816, -10.25273, 
    -10.2741, -10.29224, -10.30712, -10.31872, -10.32702, -10.332, -10.33367, 
    -10.332, -10.32702, -10.31872, -10.30712, -10.29224, -10.2741, -10.25273, 
    -10.22816, -10.20043, -10.16958, -10.13566, -10.09871, -10.0588, 
    -10.01598, -9.970306, -9.92185, -9.870676, -9.816853, -9.760451, 
    -9.701547, -9.640213, -9.576528, -9.510569, -9.442413, -9.372141, 
    -9.299832, -9.225567, -9.149424, -9.071482, -8.99182, -8.910519, 
    -8.827652, -8.743299, -8.657532, -8.570426, -8.482054, -8.392486, 
    -8.30179, -8.210036, -8.117288, -8.023608, -7.929061, -7.833705, 
    -7.737598, -7.640796, -7.543353, -7.445321, -7.346748,
  -6.612073, -6.700978, -6.789403, -6.877304, -6.964634, -7.051345, 
    -7.137385, -7.222704, -7.307246, -7.390956, -7.473776, -7.555646, 
    -7.636507, -7.716295, -7.794946, -7.872395, -7.948575, -8.023417, 
    -8.096853, -8.168813, -8.239225, -8.308019, -8.375121, -8.44046, 
    -8.503963, -8.565559, -8.625175, -8.682739, -8.738181, -8.791431, 
    -8.842422, -8.891085, -8.937356, -8.981172, -9.02247, -9.061195, 
    -9.097291, -9.130703, -9.161384, -9.189286, -9.21437, -9.236594, 
    -9.255927, -9.272337, -9.285798, -9.29629, -9.303797, -9.308306, 
    -9.30981, -9.308306, -9.303797, -9.29629, -9.285798, -9.272337, 
    -9.255927, -9.236594, -9.21437, -9.189286, -9.161384, -9.130703, 
    -9.097291, -9.061195, -9.02247, -8.981172, -8.937356, -8.891085, 
    -8.842422, -8.791431, -8.738181, -8.682739, -8.625175, -8.565559, 
    -8.503963, -8.44046, -8.375121, -8.308019, -8.239225, -8.168813, 
    -8.096853, -8.023417, -7.948575, -7.872395, -7.794946, -7.716295, 
    -7.636507, -7.555646, -7.473776, -7.390956, -7.307246, -7.222704, 
    -7.137385, -7.051345, -6.964634, -6.877304, -6.789403, -6.700978, 
    -6.612073,
  -5.877398, -5.956575, -6.035332, -6.113627, -6.19142, -6.268667, -6.345323, 
    -6.421341, -6.496675, -6.571271, -6.645081, -6.718051, -6.790126, 
    -6.86125, -6.931367, -7.000417, -7.068341, -7.135077, -7.200565, 
    -7.26474, -7.327541, -7.388902, -7.448759, -7.507047, -7.563702, 
    -7.618658, -7.671851, -7.723217, -7.772693, -7.820215, -7.865723, 
    -7.909157, -7.950458, -7.989569, -8.026436, -8.061007, -8.09323, 
    -8.123061, -8.150454, -8.175366, -8.197762, -8.217607, -8.23487, 
    -8.249522, -8.261543, -8.270913, -8.277617, -8.281642, -8.282985, 
    -8.281642, -8.277617, -8.270913, -8.261543, -8.249522, -8.23487, 
    -8.217607, -8.197762, -8.175366, -8.150454, -8.123061, -8.09323, 
    -8.061007, -8.026436, -7.989569, -7.950458, -7.909157, -7.865723, 
    -7.820215, -7.772693, -7.723217, -7.671851, -7.618658, -7.563702, 
    -7.507047, -7.448759, -7.388902, -7.327541, -7.26474, -7.200565, 
    -7.135077, -7.068341, -7.000417, -6.931367, -6.86125, -6.790126, 
    -6.718051, -6.645081, -6.571271, -6.496675, -6.421341, -6.345323, 
    -6.268667, -6.19142, -6.113627, -6.035332, -5.956575, -5.877398,
  -5.142724, -5.21212, -5.281153, -5.349786, -5.417983, -5.485706, -5.552916, 
    -5.619571, -5.68563, -5.751048, -5.815781, -5.87978, -5.943, -6.00539, 
    -6.066901, -6.12748, -6.187074, -6.245632, -6.303097, -6.359414, 
    -6.414529, -6.468383, -6.520922, -6.572086, -6.621819, -6.670065, 
    -6.716765, -6.761864, -6.805305, -6.847034, -6.886996, -6.925138, 
    -6.96141, -6.995759, -7.02814, -7.058504, -7.086808, -7.113011, 
    -7.137073, -7.158958, -7.178632, -7.196066, -7.211231, -7.224104, 
    -7.234665, -7.242897, -7.248786, -7.252323, -7.253503, -7.252323, 
    -7.248786, -7.242897, -7.234665, -7.224104, -7.211231, -7.196066, 
    -7.178632, -7.158958, -7.137073, -7.113011, -7.086808, -7.058504, 
    -7.02814, -6.995759, -6.96141, -6.925138, -6.886996, -6.847034, 
    -6.805305, -6.761864, -6.716765, -6.670065, -6.621819, -6.572086, 
    -6.520922, -6.468383, -6.414529, -6.359414, -6.303097, -6.245632, 
    -6.187074, -6.12748, -6.066901, -6.00539, -5.943, -5.87978, -5.815781, 
    -5.751048, -5.68563, -5.619571, -5.552916, -5.485706, -5.417983, 
    -5.349786, -5.281153, -5.21212, -5.142724,
  -4.408049, -4.467618, -4.526879, -4.5858, -4.64435, -4.702497, -4.760206, 
    -4.817443, -4.874171, -4.930352, -4.985948, -5.040917, -5.095221, 
    -5.148814, -5.201655, -5.253699, -5.304901, -5.355214, -5.404592, 
    -5.452987, -5.50035, -5.546633, -5.591787, -5.635764, -5.678512, 
    -5.719984, -5.760129, -5.7989, -5.836247, -5.872125, -5.906484, 
    -5.939281, -5.970469, -6.000007, -6.027852, -6.053965, -6.078306, 
    -6.100842, -6.121536, -6.140359, -6.157281, -6.172276, -6.18532, 
    -6.196393, -6.205477, -6.212557, -6.217623, -6.220666, -6.221681, 
    -6.220666, -6.217623, -6.212557, -6.205477, -6.196393, -6.18532, 
    -6.172276, -6.157281, -6.140359, -6.121536, -6.100842, -6.078306, 
    -6.053965, -6.027852, -6.000007, -5.970469, -5.939281, -5.906484, 
    -5.872125, -5.836247, -5.7989, -5.760129, -5.719984, -5.678512, 
    -5.635764, -5.591787, -5.546633, -5.50035, -5.452987, -5.404592, 
    -5.355214, -5.304901, -5.253699, -5.201655, -5.148814, -5.095221, 
    -5.040917, -4.985948, -4.930352, -4.874171, -4.817443, -4.760206, 
    -4.702497, -4.64435, -4.5858, -4.526879, -4.467618, -4.408049,
  -3.673374, -3.723077, -3.772523, -3.82169, -3.870549, -3.919074, -3.967237, 
    -4.015007, -4.062356, -4.10925, -4.155657, -4.201545, -4.246879, 
    -4.291623, -4.335741, -4.379195, -4.421948, -4.463961, -4.505196, 
    -4.545611, -4.585167, -4.623823, -4.661538, -4.69827, -4.733978, 
    -4.768622, -4.802159, -4.834549, -4.865752, -4.895727, -4.924435, 
    -4.951838, -4.977899, -5.002581, -5.025849, -5.047671, -5.068013, 
    -5.086846, -5.104141, -5.119872, -5.134015, -5.146547, -5.15745, 
    -5.166705, -5.174297, -5.180215, -5.184449, -5.186993, -5.187841, 
    -5.186993, -5.184449, -5.180215, -5.174297, -5.166705, -5.15745, 
    -5.146547, -5.134015, -5.119872, -5.104141, -5.086846, -5.068013, 
    -5.047671, -5.025849, -5.002581, -4.977899, -4.951838, -4.924435, 
    -4.895727, -4.865752, -4.834549, -4.802159, -4.768622, -4.733978, 
    -4.69827, -4.661538, -4.623823, -4.585167, -4.545611, -4.505196, 
    -4.463961, -4.421948, -4.379195, -4.335741, -4.291623, -4.246879, 
    -4.201545, -4.155657, -4.10925, -4.062356, -4.015007, -3.967237, 
    -3.919074, -3.870549, -3.82169, -3.772523, -3.723077, -3.673374,
  -2.938699, -2.978501, -3.0181, -3.057476, -3.096608, -3.135473, -3.17405, 
    -3.212315, -3.250242, -3.287808, -3.324986, -3.361748, -3.398068, 
    -3.433917, -3.469266, -3.504085, -3.538343, -3.57201, -3.605054, 
    -3.637443, -3.669145, -3.700126, -3.730354, -3.759796, -3.788419, 
    -3.816189, -3.843073, -3.869038, -3.894052, -3.918083, -3.941099, 
    -3.963069, -3.983964, -4.003754, -4.022411, -4.039908, -4.05622, 
    -4.071321, -4.08519, -4.097805, -4.109146, -4.119196, -4.127939, 
    -4.135361, -4.14145, -4.146196, -4.149592, -4.151631, -4.152311, 
    -4.151631, -4.149592, -4.146196, -4.14145, -4.135361, -4.127939, 
    -4.119196, -4.109146, -4.097805, -4.08519, -4.071321, -4.05622, 
    -4.039908, -4.022411, -4.003754, -3.983964, -3.963069, -3.941099, 
    -3.918083, -3.894052, -3.869038, -3.843073, -3.816189, -3.788419, 
    -3.759796, -3.730354, -3.700126, -3.669145, -3.637443, -3.605054, 
    -3.57201, -3.538343, -3.504085, -3.469266, -3.433917, -3.398068, 
    -3.361748, -3.324986, -3.287808, -3.250242, -3.212315, -3.17405, 
    -3.135473, -3.096608, -3.057476, -3.0181, -2.978501, -2.938699,
  -2.204024, -2.233899, -2.263623, -2.29318, -2.322554, -2.35173, -2.38069, 
    -2.409416, -2.437891, -2.466094, -2.494007, -2.52161, -2.548881, 
    -2.575799, -2.602343, -2.628489, -2.654216, -2.679499, -2.704315, 
    -2.72864, -2.752449, -2.775718, -2.798423, -2.820537, -2.842036, 
    -2.862896, -2.883091, -2.902596, -2.921387, -2.93944, -2.956731, 
    -2.973237, -2.988935, -3.003803, -3.017821, -3.030967, -3.043222, 
    -3.054569, -3.06499, -3.074468, -3.08299, -3.090542, -3.097111, 
    -3.102689, -3.107264, -3.11083, -3.113382, -3.114914, -3.115426, 
    -3.114914, -3.113382, -3.11083, -3.107264, -3.102689, -3.097111, 
    -3.090542, -3.08299, -3.074468, -3.06499, -3.054569, -3.043222, 
    -3.030967, -3.017821, -3.003803, -2.988935, -2.973237, -2.956731, 
    -2.93944, -2.921387, -2.902596, -2.883091, -2.862896, -2.842036, 
    -2.820537, -2.798423, -2.775718, -2.752449, -2.72864, -2.704315, 
    -2.679499, -2.654216, -2.628489, -2.602343, -2.575799, -2.548881, 
    -2.52161, -2.494007, -2.466094, -2.437891, -2.409416, -2.38069, -2.35173, 
    -2.322554, -2.29318, -2.263623, -2.233899, -2.204024,
  -1.46935, -1.489277, -1.509105, -1.528821, -1.548416, -1.56788, -1.587199, 
    -1.606363, -1.62536, -1.644176, -1.662799, -1.681216, -1.699411, 
    -1.717372, -1.735083, -1.752529, -1.769696, -1.786567, -1.803126, 
    -1.819359, -1.835248, -1.850776, -1.865928, -1.880687, -1.895035, 
    -1.908957, -1.922435, -1.935454, -1.947996, -1.960045, -1.971586, 
    -1.982603, -1.993082, -2.003006, -2.012363, -2.021138, -2.029319, 
    -2.036894, -2.04385, -2.050177, -2.055866, -2.060907, -2.065293, 
    -2.069016, -2.07207, -2.074451, -2.076154, -2.077178, -2.077519, 
    -2.077178, -2.076154, -2.074451, -2.07207, -2.069016, -2.065293, 
    -2.060907, -2.055866, -2.050177, -2.04385, -2.036894, -2.029319, 
    -2.021138, -2.012363, -2.003006, -1.993082, -1.982603, -1.971586, 
    -1.960045, -1.947996, -1.935454, -1.922435, -1.908957, -1.895035, 
    -1.880687, -1.865928, -1.850776, -1.835248, -1.819359, -1.803126, 
    -1.786567, -1.769696, -1.752529, -1.735083, -1.717372, -1.699411, 
    -1.681216, -1.662799, -1.644176, -1.62536, -1.606363, -1.587199, 
    -1.56788, -1.548416, -1.528821, -1.509105, -1.489277, -1.46935,
  -0.7346748, -0.744642, -0.7545591, -0.7644209, -0.7742223, -0.7839577, 
    -0.7936214, -0.8032075, -0.8127099, -0.8221223, -0.8314381, -0.8406506, 
    -0.8497528, -0.8587376, -0.8675976, -0.8763254, -0.8849133, -0.8933536, 
    -0.9016382, -0.9097592, -0.9177083, -0.9254774, -0.9330581, -0.9404421, 
    -0.947621, -0.9545865, -0.9613302, -0.9678438, -0.9741191, -0.9801481, 
    -0.9859229, -0.9914355, -0.9966785, -1.001644, -1.006326, -1.010717, 
    -1.014811, -1.018601, -1.022082, -1.025248, -1.028095, -1.030618, 
    -1.032812, -1.034675, -1.036204, -1.037395, -1.038247, -1.038759, 
    -1.03893, -1.038759, -1.038247, -1.037395, -1.036204, -1.034675, 
    -1.032812, -1.030618, -1.028095, -1.025248, -1.022082, -1.018601, 
    -1.014811, -1.010717, -1.006326, -1.001644, -0.9966785, -0.9914355, 
    -0.9859229, -0.9801481, -0.9741191, -0.9678438, -0.9613302, -0.9545865, 
    -0.947621, -0.9404421, -0.9330581, -0.9254774, -0.9177083, -0.9097592, 
    -0.9016382, -0.8933536, -0.8849133, -0.8763254, -0.8675976, -0.8587376, 
    -0.8497528, -0.8406506, -0.8314381, -0.8221223, -0.8127099, -0.8032075, 
    -0.7936214, -0.7839577, -0.7742223, -0.7644209, -0.7545591, -0.744642, 
    -0.7346748,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.7346748, 0.744642, 0.7545591, 0.7644209, 0.7742223, 0.7839577, 0.7936214, 
    0.8032075, 0.8127099, 0.8221223, 0.8314381, 0.8406506, 0.8497528, 
    0.8587376, 0.8675976, 0.8763254, 0.8849133, 0.8933536, 0.9016382, 
    0.9097592, 0.9177083, 0.9254774, 0.9330581, 0.9404421, 0.947621, 
    0.9545865, 0.9613302, 0.9678438, 0.9741191, 0.9801481, 0.9859229, 
    0.9914355, 0.9966785, 1.001644, 1.006326, 1.010717, 1.014811, 1.018601, 
    1.022082, 1.025248, 1.028095, 1.030618, 1.032812, 1.034675, 1.036204, 
    1.037395, 1.038247, 1.038759, 1.03893, 1.038759, 1.038247, 1.037395, 
    1.036204, 1.034675, 1.032812, 1.030618, 1.028095, 1.025248, 1.022082, 
    1.018601, 1.014811, 1.010717, 1.006326, 1.001644, 0.9966785, 0.9914355, 
    0.9859229, 0.9801481, 0.9741191, 0.9678438, 0.9613302, 0.9545865, 
    0.947621, 0.9404421, 0.9330581, 0.9254774, 0.9177083, 0.9097592, 
    0.9016382, 0.8933536, 0.8849133, 0.8763254, 0.8675976, 0.8587376, 
    0.8497528, 0.8406506, 0.8314381, 0.8221223, 0.8127099, 0.8032075, 
    0.7936214, 0.7839577, 0.7742223, 0.7644209, 0.7545591, 0.744642, 0.7346748,
  1.46935, 1.489277, 1.509105, 1.528821, 1.548416, 1.56788, 1.587199, 
    1.606363, 1.62536, 1.644176, 1.662799, 1.681216, 1.699411, 1.717372, 
    1.735083, 1.752529, 1.769696, 1.786567, 1.803126, 1.819359, 1.835248, 
    1.850776, 1.865928, 1.880687, 1.895035, 1.908957, 1.922435, 1.935454, 
    1.947996, 1.960045, 1.971586, 1.982603, 1.993082, 2.003006, 2.012363, 
    2.021138, 2.029319, 2.036894, 2.04385, 2.050177, 2.055866, 2.060907, 
    2.065293, 2.069016, 2.07207, 2.074451, 2.076154, 2.077178, 2.077519, 
    2.077178, 2.076154, 2.074451, 2.07207, 2.069016, 2.065293, 2.060907, 
    2.055866, 2.050177, 2.04385, 2.036894, 2.029319, 2.021138, 2.012363, 
    2.003006, 1.993082, 1.982603, 1.971586, 1.960045, 1.947996, 1.935454, 
    1.922435, 1.908957, 1.895035, 1.880687, 1.865928, 1.850776, 1.835248, 
    1.819359, 1.803126, 1.786567, 1.769696, 1.752529, 1.735083, 1.717372, 
    1.699411, 1.681216, 1.662799, 1.644176, 1.62536, 1.606363, 1.587199, 
    1.56788, 1.548416, 1.528821, 1.509105, 1.489277, 1.46935,
  2.204024, 2.233899, 2.263623, 2.29318, 2.322554, 2.35173, 2.38069, 
    2.409416, 2.437891, 2.466094, 2.494007, 2.52161, 2.548881, 2.575799, 
    2.602343, 2.628489, 2.654216, 2.679499, 2.704315, 2.72864, 2.752449, 
    2.775718, 2.798423, 2.820537, 2.842036, 2.862896, 2.883091, 2.902596, 
    2.921387, 2.93944, 2.956731, 2.973237, 2.988935, 3.003803, 3.017821, 
    3.030967, 3.043222, 3.054569, 3.06499, 3.074468, 3.08299, 3.090542, 
    3.097111, 3.102689, 3.107264, 3.11083, 3.113382, 3.114914, 3.115426, 
    3.114914, 3.113382, 3.11083, 3.107264, 3.102689, 3.097111, 3.090542, 
    3.08299, 3.074468, 3.06499, 3.054569, 3.043222, 3.030967, 3.017821, 
    3.003803, 2.988935, 2.973237, 2.956731, 2.93944, 2.921387, 2.902596, 
    2.883091, 2.862896, 2.842036, 2.820537, 2.798423, 2.775718, 2.752449, 
    2.72864, 2.704315, 2.679499, 2.654216, 2.628489, 2.602343, 2.575799, 
    2.548881, 2.52161, 2.494007, 2.466094, 2.437891, 2.409416, 2.38069, 
    2.35173, 2.322554, 2.29318, 2.263623, 2.233899, 2.204024,
  2.938699, 2.978501, 3.0181, 3.057476, 3.096608, 3.135473, 3.17405, 
    3.212315, 3.250242, 3.287808, 3.324986, 3.361748, 3.398068, 3.433917, 
    3.469266, 3.504085, 3.538343, 3.57201, 3.605054, 3.637443, 3.669145, 
    3.700126, 3.730354, 3.759796, 3.788419, 3.816189, 3.843073, 3.869038, 
    3.894052, 3.918083, 3.941099, 3.963069, 3.983964, 4.003754, 4.022411, 
    4.039908, 4.05622, 4.071321, 4.08519, 4.097805, 4.109146, 4.119196, 
    4.127939, 4.135361, 4.14145, 4.146196, 4.149592, 4.151631, 4.152311, 
    4.151631, 4.149592, 4.146196, 4.14145, 4.135361, 4.127939, 4.119196, 
    4.109146, 4.097805, 4.08519, 4.071321, 4.05622, 4.039908, 4.022411, 
    4.003754, 3.983964, 3.963069, 3.941099, 3.918083, 3.894052, 3.869038, 
    3.843073, 3.816189, 3.788419, 3.759796, 3.730354, 3.700126, 3.669145, 
    3.637443, 3.605054, 3.57201, 3.538343, 3.504085, 3.469266, 3.433917, 
    3.398068, 3.361748, 3.324986, 3.287808, 3.250242, 3.212315, 3.17405, 
    3.135473, 3.096608, 3.057476, 3.0181, 2.978501, 2.938699,
  3.673374, 3.723077, 3.772523, 3.82169, 3.870549, 3.919074, 3.967237, 
    4.015007, 4.062356, 4.10925, 4.155657, 4.201545, 4.246879, 4.291623, 
    4.335741, 4.379195, 4.421948, 4.463961, 4.505196, 4.545611, 4.585167, 
    4.623823, 4.661538, 4.69827, 4.733978, 4.768622, 4.802159, 4.834549, 
    4.865752, 4.895727, 4.924435, 4.951838, 4.977899, 5.002581, 5.025849, 
    5.047671, 5.068013, 5.086846, 5.104141, 5.119872, 5.134015, 5.146547, 
    5.15745, 5.166705, 5.174297, 5.180215, 5.184449, 5.186993, 5.187841, 
    5.186993, 5.184449, 5.180215, 5.174297, 5.166705, 5.15745, 5.146547, 
    5.134015, 5.119872, 5.104141, 5.086846, 5.068013, 5.047671, 5.025849, 
    5.002581, 4.977899, 4.951838, 4.924435, 4.895727, 4.865752, 4.834549, 
    4.802159, 4.768622, 4.733978, 4.69827, 4.661538, 4.623823, 4.585167, 
    4.545611, 4.505196, 4.463961, 4.421948, 4.379195, 4.335741, 4.291623, 
    4.246879, 4.201545, 4.155657, 4.10925, 4.062356, 4.015007, 3.967237, 
    3.919074, 3.870549, 3.82169, 3.772523, 3.723077, 3.673374,
  4.408049, 4.467618, 4.526879, 4.5858, 4.64435, 4.702497, 4.760206, 
    4.817443, 4.874171, 4.930352, 4.985948, 5.040917, 5.095221, 5.148814, 
    5.201655, 5.253699, 5.304901, 5.355214, 5.404592, 5.452987, 5.50035, 
    5.546633, 5.591787, 5.635764, 5.678512, 5.719984, 5.760129, 5.7989, 
    5.836247, 5.872125, 5.906484, 5.939281, 5.970469, 6.000007, 6.027852, 
    6.053965, 6.078306, 6.100842, 6.121536, 6.140359, 6.157281, 6.172276, 
    6.18532, 6.196393, 6.205477, 6.212557, 6.217623, 6.220666, 6.221681, 
    6.220666, 6.217623, 6.212557, 6.205477, 6.196393, 6.18532, 6.172276, 
    6.157281, 6.140359, 6.121536, 6.100842, 6.078306, 6.053965, 6.027852, 
    6.000007, 5.970469, 5.939281, 5.906484, 5.872125, 5.836247, 5.7989, 
    5.760129, 5.719984, 5.678512, 5.635764, 5.591787, 5.546633, 5.50035, 
    5.452987, 5.404592, 5.355214, 5.304901, 5.253699, 5.201655, 5.148814, 
    5.095221, 5.040917, 4.985948, 4.930352, 4.874171, 4.817443, 4.760206, 
    4.702497, 4.64435, 4.5858, 4.526879, 4.467618, 4.408049,
  5.142724, 5.21212, 5.281153, 5.349786, 5.417983, 5.485706, 5.552916, 
    5.619571, 5.68563, 5.751048, 5.815781, 5.87978, 5.943, 6.00539, 6.066901, 
    6.12748, 6.187074, 6.245632, 6.303097, 6.359414, 6.414529, 6.468383, 
    6.520922, 6.572086, 6.621819, 6.670065, 6.716765, 6.761864, 6.805305, 
    6.847034, 6.886996, 6.925138, 6.96141, 6.995759, 7.02814, 7.058504, 
    7.086808, 7.113011, 7.137073, 7.158958, 7.178632, 7.196066, 7.211231, 
    7.224104, 7.234665, 7.242897, 7.248786, 7.252323, 7.253503, 7.252323, 
    7.248786, 7.242897, 7.234665, 7.224104, 7.211231, 7.196066, 7.178632, 
    7.158958, 7.137073, 7.113011, 7.086808, 7.058504, 7.02814, 6.995759, 
    6.96141, 6.925138, 6.886996, 6.847034, 6.805305, 6.761864, 6.716765, 
    6.670065, 6.621819, 6.572086, 6.520922, 6.468383, 6.414529, 6.359414, 
    6.303097, 6.245632, 6.187074, 6.12748, 6.066901, 6.00539, 5.943, 5.87978, 
    5.815781, 5.751048, 5.68563, 5.619571, 5.552916, 5.485706, 5.417983, 
    5.349786, 5.281153, 5.21212, 5.142724,
  5.877398, 5.956575, 6.035332, 6.113627, 6.19142, 6.268667, 6.345323, 
    6.421341, 6.496675, 6.571271, 6.645081, 6.718051, 6.790126, 6.86125, 
    6.931367, 7.000417, 7.068341, 7.135077, 7.200565, 7.26474, 7.327541, 
    7.388902, 7.448759, 7.507047, 7.563702, 7.618658, 7.671851, 7.723217, 
    7.772693, 7.820215, 7.865723, 7.909157, 7.950458, 7.989569, 8.026436, 
    8.061007, 8.09323, 8.123061, 8.150454, 8.175366, 8.197762, 8.217607, 
    8.23487, 8.249522, 8.261543, 8.270913, 8.277617, 8.281642, 8.282985, 
    8.281642, 8.277617, 8.270913, 8.261543, 8.249522, 8.23487, 8.217607, 
    8.197762, 8.175366, 8.150454, 8.123061, 8.09323, 8.061007, 8.026436, 
    7.989569, 7.950458, 7.909157, 7.865723, 7.820215, 7.772693, 7.723217, 
    7.671851, 7.618658, 7.563702, 7.507047, 7.448759, 7.388902, 7.327541, 
    7.26474, 7.200565, 7.135077, 7.068341, 7.000417, 6.931367, 6.86125, 
    6.790126, 6.718051, 6.645081, 6.571271, 6.496675, 6.421341, 6.345323, 
    6.268667, 6.19142, 6.113627, 6.035332, 5.956575, 5.877398,
  6.612073, 6.700978, 6.789403, 6.877304, 6.964634, 7.051345, 7.137385, 
    7.222704, 7.307246, 7.390956, 7.473776, 7.555646, 7.636507, 7.716295, 
    7.794946, 7.872395, 7.948575, 8.023417, 8.096853, 8.168813, 8.239225, 
    8.308019, 8.375121, 8.44046, 8.503963, 8.565559, 8.625175, 8.682739, 
    8.738181, 8.791431, 8.842422, 8.891085, 8.937356, 8.981172, 9.02247, 
    9.061195, 9.097291, 9.130703, 9.161384, 9.189286, 9.21437, 9.236594, 
    9.255927, 9.272337, 9.285798, 9.29629, 9.303797, 9.308306, 9.30981, 
    9.308306, 9.303797, 9.29629, 9.285798, 9.272337, 9.255927, 9.236594, 
    9.21437, 9.189286, 9.161384, 9.130703, 9.097291, 9.061195, 9.02247, 
    8.981172, 8.937356, 8.891085, 8.842422, 8.791431, 8.738181, 8.682739, 
    8.625175, 8.565559, 8.503963, 8.44046, 8.375121, 8.308019, 8.239225, 
    8.168813, 8.096853, 8.023417, 7.948575, 7.872395, 7.794946, 7.716295, 
    7.636507, 7.555646, 7.473776, 7.390956, 7.307246, 7.222704, 7.137385, 
    7.051345, 6.964634, 6.877304, 6.789403, 6.700978, 6.612073,
  7.346748, 7.445321, 7.543353, 7.640796, 7.737598, 7.833705, 7.929061, 
    8.023608, 8.117288, 8.210036, 8.30179, 8.392486, 8.482054, 8.570426, 
    8.657532, 8.743299, 8.827652, 8.910519, 8.99182, 9.071482, 9.149424, 
    9.225567, 9.299832, 9.372141, 9.442413, 9.510569, 9.576528, 9.640213, 
    9.701547, 9.760451, 9.816853, 9.870676, 9.92185, 9.970306, 10.01598, 
    10.0588, 10.09871, 10.13566, 10.16958, 10.20043, 10.22816, 10.25273, 
    10.2741, 10.29224, 10.30712, 10.31872, 10.32702, 10.332, 10.33367, 
    10.332, 10.32702, 10.31872, 10.30712, 10.29224, 10.2741, 10.25273, 
    10.22816, 10.20043, 10.16958, 10.13566, 10.09871, 10.0588, 10.01598, 
    9.970306, 9.92185, 9.870676, 9.816853, 9.760451, 9.701547, 9.640213, 
    9.576528, 9.510569, 9.442413, 9.372141, 9.299832, 9.225567, 9.149424, 
    9.071482, 8.99182, 8.910519, 8.827652, 8.743299, 8.657532, 8.570426, 
    8.482054, 8.392486, 8.30179, 8.210036, 8.117288, 8.023608, 7.929061, 
    7.833705, 7.737598, 7.640796, 7.543353, 7.445321, 7.346748,
  8.081423, 8.189597, 8.297169, 8.404083, 8.510284, 8.615713, 8.720308, 
    8.824006, 8.926742, 9.028447, 9.129053, 9.228487, 9.326677, 9.423547, 
    9.519018, 9.613013, 9.705451, 9.79625, 9.885328, 9.972599, 10.05798, 
    10.14138, 10.22272, 10.30191, 10.37886, 10.45349, 10.52571, 10.59543, 
    10.66257, 10.72705, 10.78878, 10.84769, 10.90369, 10.95672, 11.0067, 
    11.05355, 11.09722, 11.13764, 11.17476, 11.2085, 11.23884, 11.26572, 
    11.2891, 11.30894, 11.32522, 11.33791, 11.34698, 11.35243, 11.35425, 
    11.35243, 11.34698, 11.33791, 11.32522, 11.30894, 11.2891, 11.26572, 
    11.23884, 11.2085, 11.17476, 11.13764, 11.09722, 11.05355, 11.0067, 
    10.95672, 10.90369, 10.84769, 10.78878, 10.72705, 10.66257, 10.59543, 
    10.52571, 10.45349, 10.37886, 10.30191, 10.22272, 10.14138, 10.05798, 
    9.972599, 9.885328, 9.79625, 9.705451, 9.613013, 9.519018, 9.423547, 
    9.326677, 9.228487, 9.129053, 9.028447, 8.926742, 8.824006, 8.720308, 
    8.615713, 8.510284, 8.404083, 8.297169, 8.189597, 8.081423,
  8.816097, 8.933801, 9.050837, 9.167146, 9.282667, 9.397336, 9.511086, 
    9.623848, 9.735553, 9.846126, 9.955491, 10.06357, 10.17029, 10.27556, 
    10.3793, 10.48143, 10.58185, 10.68048, 10.77724, 10.87202, 10.96474, 
    11.0553, 11.14361, 11.22959, 11.31312, 11.39412, 11.47251, 11.54817, 
    11.62103, 11.691, 11.75798, 11.82189, 11.88264, 11.94017, 11.99438, 
    12.0452, 12.09256, 12.1364, 12.17664, 12.21324, 12.24614, 12.27528, 
    12.30063, 12.32215, 12.3398, 12.35355, 12.36339, 12.3693, 12.37127, 
    12.3693, 12.36339, 12.35355, 12.3398, 12.32215, 12.30063, 12.27528, 
    12.24614, 12.21324, 12.17664, 12.1364, 12.09256, 12.0452, 11.99438, 
    11.94017, 11.88264, 11.82189, 11.75798, 11.691, 11.62103, 11.54817, 
    11.47251, 11.39412, 11.31312, 11.22959, 11.14361, 11.0553, 10.96474, 
    10.87202, 10.77724, 10.68048, 10.58185, 10.48143, 10.3793, 10.27556, 
    10.17029, 10.06357, 9.955491, 9.846126, 9.735553, 9.623848, 9.511086, 
    9.397336, 9.282667, 9.167146, 9.050837, 8.933801, 8.816097,
  9.550773, 9.677926, 9.804344, 9.929964, 10.05472, 10.17854, 10.30135, 
    10.42309, 10.54366, 10.66301, 10.78103, 10.89766, 11.0128, 11.12637, 
    11.23828, 11.34843, 11.45673, 11.5631, 11.66742, 11.7696, 11.86955, 
    11.96717, 12.06235, 12.155, 12.24501, 12.33229, 12.41673, 12.49824, 
    12.57673, 12.65208, 12.72422, 12.79304, 12.85847, 12.9204, 12.97877, 
    13.03348, 13.08447, 13.13165, 13.17497, 13.21437, 13.24977, 13.28114, 
    13.30842, 13.33158, 13.35057, 13.36537, 13.37596, 13.38232, 13.38444, 
    13.38232, 13.37596, 13.36537, 13.35057, 13.33158, 13.30842, 13.28114, 
    13.24977, 13.21437, 13.17497, 13.13165, 13.08447, 13.03348, 12.97877, 
    12.9204, 12.85847, 12.79304, 12.72422, 12.65208, 12.57673, 12.49824, 
    12.41673, 12.33229, 12.24501, 12.155, 12.06235, 11.96717, 11.86955, 
    11.7696, 11.66742, 11.5631, 11.45673, 11.34843, 11.23828, 11.12637, 
    11.0128, 10.89766, 10.78103, 10.66301, 10.54366, 10.42309, 10.30135, 
    10.17854, 10.05472, 9.929964, 9.804344, 9.677926, 9.550773,
  10.28545, 10.42197, 10.55768, 10.69252, 10.82641, 10.95929, 11.09107, 
    11.22167, 11.35102, 11.47903, 11.60561, 11.73068, 11.85414, 11.97589, 
    12.09585, 12.21391, 12.32998, 12.44396, 12.55573, 12.66521, 12.77227, 
    12.87683, 12.97877, 13.07798, 13.17436, 13.2678, 13.3582, 13.44545, 
    13.52945, 13.61009, 13.68729, 13.76093, 13.83093, 13.89719, 13.95963, 
    14.01815, 14.07269, 14.12316, 14.16949, 14.21162, 14.24948, 14.28303, 
    14.3122, 14.33696, 14.35726, 14.37309, 14.38441, 14.39121, 14.39348, 
    14.39121, 14.38441, 14.37309, 14.35726, 14.33696, 14.3122, 14.28303, 
    14.24948, 14.21162, 14.16949, 14.12316, 14.07269, 14.01815, 13.95963, 
    13.89719, 13.83093, 13.76093, 13.68729, 13.61009, 13.52945, 13.44545, 
    13.3582, 13.2678, 13.17436, 13.07798, 12.97877, 12.87683, 12.77227, 
    12.66521, 12.55573, 12.44396, 12.32998, 12.21391, 12.09585, 11.97589, 
    11.85414, 11.73068, 11.60561, 11.47903, 11.35102, 11.22167, 11.09107, 
    10.95929, 10.82641, 10.69252, 10.55768, 10.42197, 10.28545,
  11.02012, 11.16591, 11.31083, 11.45479, 11.59772, 11.73955, 11.88019, 
    12.01956, 12.15757, 12.29414, 12.42916, 12.56255, 12.6942, 12.82403, 
    12.95192, 13.07777, 13.20149, 13.32295, 13.44206, 13.5587, 13.67276, 
    13.78413, 13.8927, 13.99836, 14.10098, 14.20047, 14.29671, 14.38959, 
    14.479, 14.56483, 14.64697, 14.72534, 14.79981, 14.87031, 14.93673, 
    14.99899, 15.05699, 15.11067, 15.15995, 15.20475, 15.24501, 15.28068, 
    15.3117, 15.33803, 15.35962, 15.37645, 15.38849, 15.39572, 15.39813, 
    15.39572, 15.38849, 15.37645, 15.35962, 15.33803, 15.3117, 15.28068, 
    15.24501, 15.20475, 15.15995, 15.11067, 15.05699, 14.99899, 14.93673, 
    14.87031, 14.79981, 14.72534, 14.64697, 14.56483, 14.479, 14.38959, 
    14.29671, 14.20047, 14.10098, 13.99836, 13.8927, 13.78413, 13.67276, 
    13.5587, 13.44206, 13.32295, 13.20149, 13.07777, 12.95192, 12.82403, 
    12.6942, 12.56255, 12.42916, 12.29414, 12.15757, 12.01956, 11.88019, 
    11.73955, 11.59772, 11.45479, 11.31083, 11.16591, 11.02012,
  11.7548, 11.90976, 12.06378, 12.21676, 12.36863, 12.5193, 12.66869, 
    12.81671, 12.96326, 13.10826, 13.2516, 13.39319, 13.53292, 13.67069, 
    13.80638, 13.9399, 14.07113, 14.19996, 14.32627, 14.44994, 14.57087, 
    14.68893, 14.804, 14.91598, 15.02473, 15.13014, 15.2321, 15.33048, 
    15.42518, 15.51608, 15.60307, 15.68605, 15.7649, 15.83954, 15.90985, 
    15.97575, 16.03714, 16.09396, 16.1461, 16.19351, 16.23612, 16.27386, 
    16.30668, 16.33454, 16.35738, 16.37519, 16.38792, 16.39557, 16.39812, 
    16.39557, 16.38792, 16.37519, 16.35738, 16.33454, 16.30668, 16.27386, 
    16.23612, 16.19351, 16.1461, 16.09396, 16.03714, 15.97575, 15.90985, 
    15.83954, 15.7649, 15.68605, 15.60307, 15.51608, 15.42518, 15.33048, 
    15.2321, 15.13014, 15.02473, 14.91598, 14.804, 14.68893, 14.57087, 
    14.44994, 14.32627, 14.19996, 14.07113, 13.9399, 13.80638, 13.67069, 
    13.53292, 13.39319, 13.2516, 13.10826, 12.96326, 12.81671, 12.66869, 
    12.5193, 12.36863, 12.21676, 12.06378, 11.90976, 11.7548,
  12.48947, 12.65351, 12.81652, 12.97841, 13.1391, 13.2985, 13.45652, 
    13.61306, 13.76804, 13.92135, 14.07288, 14.22254, 14.37021, 14.51579, 
    14.65916, 14.8002, 14.93881, 15.07486, 15.20823, 15.33881, 15.46647, 
    15.59108, 15.71253, 15.83068, 15.94542, 16.05663, 16.16418, 16.26795, 
    16.36782, 16.46367, 16.55539, 16.64287, 16.72599, 16.80466, 16.87877, 
    16.94822, 17.01292, 17.07278, 17.12773, 17.17768, 17.22256, 17.26232, 
    17.2969, 17.32624, 17.3503, 17.36906, 17.38247, 17.39053, 17.39322, 
    17.39053, 17.38247, 17.36906, 17.3503, 17.32624, 17.2969, 17.26232, 
    17.22256, 17.17768, 17.12773, 17.07278, 17.01292, 16.94822, 16.87877, 
    16.80466, 16.72599, 16.64287, 16.55539, 16.46367, 16.36782, 16.26795, 
    16.16418, 16.05663, 15.94542, 15.83068, 15.71253, 15.59108, 15.46647, 
    15.33881, 15.20823, 15.07486, 14.93881, 14.8002, 14.65916, 14.51579, 
    14.37021, 14.22254, 14.07288, 13.92135, 13.76804, 13.61306, 13.45652, 
    13.2985, 13.1391, 12.97841, 12.81652, 12.65351, 12.48947,
  13.22415, 13.39715, 13.56903, 13.73972, 13.90911, 14.07711, 14.24364, 
    14.40859, 14.57185, 14.73334, 14.89293, 15.05052, 15.20599, 15.35924, 
    15.51014, 15.65857, 15.80442, 15.94755, 16.08784, 16.22518, 16.35942, 
    16.49044, 16.61812, 16.74232, 16.86292, 16.97978, 17.09279, 17.20181, 
    17.30672, 17.4074, 17.50373, 17.5956, 17.68288, 17.76548, 17.84328, 
    17.91618, 17.9841, 18.04693, 18.1046, 18.15702, 18.20412, 18.24584, 
    18.28212, 18.31291, 18.33815, 18.35783, 18.3719, 18.38036, 18.38318, 
    18.38036, 18.3719, 18.35783, 18.33815, 18.31291, 18.28212, 18.24584, 
    18.20412, 18.15702, 18.1046, 18.04693, 17.9841, 17.91618, 17.84328, 
    17.76548, 17.68288, 17.5956, 17.50373, 17.4074, 17.30672, 17.20181, 
    17.09279, 16.97978, 16.86292, 16.74232, 16.61812, 16.49044, 16.35942, 
    16.22518, 16.08784, 15.94755, 15.80442, 15.65857, 15.51014, 15.35924, 
    15.20599, 15.05052, 14.89293, 14.73334, 14.57185, 14.40859, 14.24364, 
    14.07711, 13.90911, 13.73972, 13.56903, 13.39715, 13.22415,
  13.95882, 14.14067, 14.32132, 14.50067, 14.67863, 14.85512, 15.03002, 
    15.20323, 15.37465, 15.54417, 15.71168, 15.87706, 16.0402, 16.20097, 
    16.35925, 16.51492, 16.66785, 16.81791, 16.96498, 17.10892, 17.2496, 
    17.38689, 17.52065, 17.65075, 17.77705, 17.89944, 18.01776, 18.1319, 
    18.24172, 18.34711, 18.44792, 18.54405, 18.63538, 18.7218, 18.80319, 
    18.87945, 18.95048, 19.0162, 19.0765, 19.13132, 19.18058, 19.2242, 
    19.26213, 19.29432, 19.32071, 19.34128, 19.356, 19.36483, 19.36778, 
    19.36483, 19.356, 19.34128, 19.32071, 19.29432, 19.26213, 19.2242, 
    19.18058, 19.13132, 19.0765, 19.0162, 18.95048, 18.87945, 18.80319, 
    18.7218, 18.63538, 18.54405, 18.44792, 18.34711, 18.24172, 18.1319, 
    18.01776, 17.89944, 17.77705, 17.65075, 17.52065, 17.38689, 17.2496, 
    17.10892, 16.96498, 16.81791, 16.66785, 16.51492, 16.35925, 16.20097, 
    16.0402, 15.87706, 15.71168, 15.54417, 15.37465, 15.20323, 15.03002, 
    14.85512, 14.67863, 14.50067, 14.32132, 14.14067, 13.95882,
  14.6935, 14.88407, 15.07335, 15.26124, 15.44765, 15.63248, 15.81561, 
    15.99695, 16.17639, 16.3538, 16.52908, 16.7021, 16.87274, 17.04088, 
    17.20639, 17.36914, 17.52901, 17.68585, 17.83953, 17.98992, 18.13688, 
    18.28028, 18.41997, 18.55582, 18.68769, 18.81544, 18.93895, 19.05806, 
    19.17266, 19.28261, 19.38778, 19.48806, 19.58331, 19.67343, 19.7583, 
    19.83782, 19.91188, 19.98038, 20.04325, 20.10039, 20.15172, 20.19719, 
    20.23672, 20.27026, 20.29777, 20.3192, 20.33454, 20.34374, 20.34682, 
    20.34374, 20.33454, 20.3192, 20.29777, 20.27026, 20.23672, 20.19719, 
    20.15172, 20.10039, 20.04325, 19.98038, 19.91188, 19.83782, 19.7583, 
    19.67343, 19.58331, 19.48806, 19.38778, 19.28261, 19.17266, 19.05806, 
    18.93895, 18.81544, 18.68769, 18.55582, 18.41997, 18.28028, 18.13688, 
    17.98992, 17.83953, 17.68585, 17.52901, 17.36914, 17.20639, 17.04088, 
    16.87274, 16.7021, 16.52908, 16.3538, 16.17639, 15.99695, 15.81561, 
    15.63248, 15.44765, 15.26124, 15.07335, 14.88407, 14.6935,
  15.42817, 15.62734, 15.82513, 16.02143, 16.21614, 16.40917, 16.6004, 
    16.78971, 16.97701, 17.16216, 17.34505, 17.52556, 17.70355, 17.8789, 
    18.05148, 18.22116, 18.38779, 18.55125, 18.71139, 18.86807, 19.02115, 
    19.1705, 19.31597, 19.45741, 19.59469, 19.72766, 19.85619, 19.98014, 
    20.09937, 20.21375, 20.32315, 20.42744, 20.5265, 20.6202, 20.70844, 
    20.79111, 20.8681, 20.9393, 21.00464, 21.06402, 21.11737, 21.16462, 
    21.20569, 21.24054, 21.26912, 21.29139, 21.30732, 21.31689, 21.32008, 
    21.31689, 21.30732, 21.29139, 21.26912, 21.24054, 21.20569, 21.16462, 
    21.11737, 21.06402, 21.00464, 20.9393, 20.8681, 20.79111, 20.70844, 
    20.6202, 20.5265, 20.42744, 20.32315, 20.21375, 20.09937, 19.98014, 
    19.85619, 19.72766, 19.59469, 19.45741, 19.31597, 19.1705, 19.02115, 
    18.86807, 18.71139, 18.55125, 18.38779, 18.22116, 18.05148, 17.8789, 
    17.70355, 17.52556, 17.34505, 17.16216, 16.97701, 16.78971, 16.6004, 
    16.40917, 16.21614, 16.02143, 15.82513, 15.62734, 15.42817,
  16.16285, 16.37048, 16.57663, 16.7812, 16.98408, 17.18516, 17.38433, 
    17.58147, 17.77647, 17.96921, 18.15956, 18.34738, 18.53256, 18.71496, 
    18.89445, 19.07088, 19.24412, 19.41402, 19.58045, 19.74325, 19.9023, 
    20.05743, 20.20851, 20.35538, 20.49791, 20.63595, 20.76936, 20.89799, 
    21.02171, 21.14038, 21.25386, 21.36204, 21.46477, 21.56195, 21.65344, 
    21.73915, 21.81896, 21.89278, 21.9605, 22.02205, 22.07734, 22.1263, 
    22.16886, 22.20498, 22.23459, 22.25766, 22.27417, 22.28408, 22.28739, 
    22.28408, 22.27417, 22.25766, 22.23459, 22.20498, 22.16886, 22.1263, 
    22.07734, 22.02205, 21.9605, 21.89278, 21.81896, 21.73915, 21.65344, 
    21.56195, 21.46477, 21.36204, 21.25386, 21.14038, 21.02171, 20.89799, 
    20.76936, 20.63595, 20.49791, 20.35538, 20.20851, 20.05743, 19.9023, 
    19.74325, 19.58045, 19.41402, 19.24412, 19.07088, 18.89445, 18.71496, 
    18.53256, 18.34738, 18.15956, 17.96921, 17.77647, 17.58147, 17.38433, 
    17.18516, 16.98408, 16.7812, 16.57663, 16.37048, 16.16285,
  16.89752, 17.11348, 17.32786, 17.54054, 17.75143, 17.96042, 18.16737, 
    18.37219, 18.57473, 18.77489, 18.97252, 19.16751, 19.35971, 19.54898, 
    19.7352, 19.91821, 20.09789, 20.27407, 20.44661, 20.61537, 20.7802, 
    20.94095, 21.09747, 21.24961, 21.39723, 21.54018, 21.6783, 21.81147, 
    21.93953, 22.06234, 22.17978, 22.2917, 22.39799, 22.49851, 22.59314, 
    22.68178, 22.76431, 22.84064, 22.91066, 22.97429, 23.03145, 23.08206, 
    23.12605, 23.16338, 23.19399, 23.21784, 23.2349, 23.24514, 23.24856, 
    23.24514, 23.2349, 23.21784, 23.19399, 23.16338, 23.12605, 23.08206, 
    23.03145, 22.97429, 22.91066, 22.84064, 22.76431, 22.68178, 22.59314, 
    22.49851, 22.39799, 22.2917, 22.17978, 22.06234, 21.93953, 21.81147, 
    21.6783, 21.54018, 21.39723, 21.24961, 21.09747, 20.94095, 20.7802, 
    20.61537, 20.44661, 20.27407, 20.09789, 19.91821, 19.7352, 19.54898, 
    19.35971, 19.16751, 18.97252, 18.77489, 18.57473, 18.37219, 18.16737, 
    17.96042, 17.75143, 17.54054, 17.32786, 17.11348, 16.89752,
  17.63219, 17.85633, 18.07879, 18.29944, 18.51819, 18.73492, 18.9495, 
    19.16182, 19.37174, 19.57915, 19.7839, 19.98587, 20.18491, 20.38089, 
    20.57367, 20.76309, 20.94901, 21.13129, 21.30978, 21.48432, 21.65476, 
    21.82095, 21.98275, 22.13999, 22.29253, 22.44022, 22.5829, 22.72045, 
    22.85269, 22.97951, 23.10075, 23.21629, 23.32599, 23.42973, 23.52739, 
    23.61885, 23.704, 23.78273, 23.85496, 23.92059, 23.97954, 24.03174, 
    24.07711, 24.1156, 24.14717, 24.17175, 24.18934, 24.19991, 24.20343, 
    24.19991, 24.18934, 24.17175, 24.14717, 24.1156, 24.07711, 24.03174, 
    23.97954, 23.92059, 23.85496, 23.78273, 23.704, 23.61885, 23.52739, 
    23.42973, 23.32599, 23.21629, 23.10075, 22.97951, 22.85269, 22.72045, 
    22.5829, 22.44022, 22.29253, 22.13999, 21.98275, 21.82095, 21.65476, 
    21.48432, 21.30978, 21.13129, 20.94901, 20.76309, 20.57367, 20.38089, 
    20.18491, 19.98587, 19.7839, 19.57915, 19.37174, 19.16182, 18.9495, 
    18.73492, 18.51819, 18.29944, 18.07879, 17.85633, 17.63219,
  18.36687, 18.59904, 18.82941, 19.05788, 19.28433, 19.50863, 19.73068, 
    19.95033, 20.16746, 20.38194, 20.59364, 20.80241, 21.00812, 21.21062, 
    21.40977, 21.60542, 21.79742, 21.98561, 22.16986, 22.35, 22.52588, 
    22.69734, 22.86423, 23.0264, 23.18369, 23.33596, 23.48304, 23.6248, 
    23.76108, 23.89175, 24.01665, 24.13567, 24.24865, 24.35549, 24.45604, 
    24.55021, 24.63787, 24.71892, 24.79326, 24.86081, 24.92148, 24.97519, 
    25.02188, 25.06149, 25.09396, 25.11926, 25.13736, 25.14822, 25.15185, 
    25.14822, 25.13736, 25.11926, 25.09396, 25.06149, 25.02188, 24.97519, 
    24.92148, 24.86081, 24.79326, 24.71892, 24.63787, 24.55021, 24.45604, 
    24.35549, 24.24865, 24.13567, 24.01665, 23.89175, 23.76108, 23.6248, 
    23.48304, 23.33596, 23.18369, 23.0264, 22.86423, 22.69734, 22.52588, 
    22.35, 22.16986, 21.98561, 21.79742, 21.60542, 21.40977, 21.21062, 
    21.00812, 20.80241, 20.59364, 20.38194, 20.16746, 19.95033, 19.73068, 
    19.50863, 19.28433, 19.05788, 18.82941, 18.59904, 18.36687,
  19.10155, 19.34159, 19.57973, 19.81585, 20.04982, 20.28154, 20.51087, 
    20.73768, 20.96184, 21.18322, 21.40168, 21.61708, 21.82927, 22.03811, 
    22.24345, 22.44514, 22.64302, 22.83695, 23.02677, 23.21232, 23.39345, 
    23.57, 23.74181, 23.90874, 24.07061, 24.22728, 24.3786, 24.52441, 
    24.66457, 24.79893, 24.92736, 25.0497, 25.16584, 25.27564, 25.37897, 
    25.47573, 25.56579, 25.64905, 25.72542, 25.7948, 25.85711, 25.91227, 
    25.96022, 26.00089, 26.03424, 26.06021, 26.0788, 26.08995, 26.09367, 
    26.08995, 26.0788, 26.06021, 26.03424, 26.00089, 25.96022, 25.91227, 
    25.85711, 25.7948, 25.72542, 25.64905, 25.56579, 25.47573, 25.37897, 
    25.27564, 25.16584, 25.0497, 24.92736, 24.79893, 24.66457, 24.52441, 
    24.3786, 24.22728, 24.07061, 23.90874, 23.74181, 23.57, 23.39345, 
    23.21232, 23.02677, 22.83695, 22.64302, 22.44514, 22.24345, 22.03811, 
    21.82927, 21.61708, 21.40168, 21.18322, 20.96184, 20.73768, 20.51087, 
    20.28154, 20.04982, 19.81585, 19.57973, 19.34159, 19.10155,
  19.83622, 20.08398, 20.32972, 20.57332, 20.81466, 21.05361, 21.29005, 
    21.52384, 21.75485, 21.98295, 22.20798, 22.42981, 22.6483, 22.86328, 
    23.07462, 23.28216, 23.48574, 23.68522, 23.88042, 24.0712, 24.2574, 
    24.43885, 24.6154, 24.7869, 24.95318, 25.11408, 25.26947, 25.41917, 
    25.56305, 25.70096, 25.83275, 25.95829, 26.07744, 26.19007, 26.29606, 
    26.39529, 26.48764, 26.57302, 26.65132, 26.72244, 26.78632, 26.84286, 
    26.892, 26.93369, 26.96786, 26.99449, 27.01353, 27.02497, 27.02878, 
    27.02497, 27.01353, 26.99449, 26.96786, 26.93369, 26.892, 26.84286, 
    26.78632, 26.72244, 26.65132, 26.57302, 26.48764, 26.39529, 26.29606, 
    26.19007, 26.07744, 25.95829, 25.83275, 25.70096, 25.56305, 25.41917, 
    25.26947, 25.11408, 24.95318, 24.7869, 24.6154, 24.43885, 24.2574, 
    24.0712, 23.88042, 23.68522, 23.48574, 23.28216, 23.07462, 22.86328, 
    22.6483, 22.42981, 22.20798, 21.98295, 21.75485, 21.52384, 21.29005, 
    21.05361, 20.81466, 20.57332, 20.32972, 20.08398, 19.83622,
  20.57089, 20.8262, 21.07937, 21.33028, 21.5788, 21.82482, 22.06818, 
    22.30877, 22.54645, 22.78106, 23.01249, 23.24056, 23.46515, 23.68609, 
    23.90323, 24.11643, 24.32551, 24.53034, 24.73074, 24.92656, 25.11763, 
    25.3038, 25.48491, 25.6608, 25.8313, 25.99627, 26.15555, 26.30898, 
    26.45642, 26.59771, 26.73272, 26.86131, 26.98333, 27.09867, 27.20719, 
    27.30877, 27.40331, 27.4907, 27.57083, 27.64362, 27.70898, 27.76684, 
    27.81712, 27.85977, 27.89473, 27.92197, 27.94145, 27.95315, 27.95705, 
    27.95315, 27.94145, 27.92197, 27.89473, 27.85977, 27.81712, 27.76684, 
    27.70898, 27.64362, 27.57083, 27.4907, 27.40331, 27.30877, 27.20719, 
    27.09867, 26.98333, 26.86131, 26.73272, 26.59771, 26.45642, 26.30898, 
    26.15555, 25.99627, 25.8313, 25.6608, 25.48491, 25.3038, 25.11763, 
    24.92656, 24.73074, 24.53034, 24.32551, 24.11643, 23.90323, 23.68609, 
    23.46515, 23.24056, 23.01249, 22.78106, 22.54645, 22.30877, 22.06818, 
    21.82482, 21.5788, 21.33028, 21.07937, 20.8262, 20.57089,
  21.30557, 21.56826, 21.82868, 22.08672, 22.34225, 22.59513, 22.84524, 
    23.09244, 23.33659, 23.57754, 23.81515, 24.04927, 24.27976, 24.50646, 
    24.72922, 24.94787, 25.16227, 25.37224, 25.57764, 25.77831, 25.97407, 
    26.16477, 26.35024, 26.53034, 26.70489, 26.87375, 27.03675, 27.19374, 
    27.34457, 27.4891, 27.62718, 27.75867, 27.88343, 28.00133, 28.11226, 
    28.21608, 28.3127, 28.40199, 28.48387, 28.55823, 28.625, 28.6841, 
    28.73546, 28.77902, 28.81473, 28.84255, 28.86244, 28.87439, 28.87837, 
    28.87439, 28.86244, 28.84255, 28.81473, 28.77902, 28.73546, 28.6841, 
    28.625, 28.55823, 28.48387, 28.40199, 28.3127, 28.21608, 28.11226, 
    28.00133, 27.88343, 27.75867, 27.62718, 27.4891, 27.34457, 27.19374, 
    27.03675, 26.87375, 26.70489, 26.53034, 26.35024, 26.16477, 25.97407, 
    25.77831, 25.57764, 25.37224, 25.16227, 24.94787, 24.72922, 24.50646, 
    24.27976, 24.04927, 23.81515, 23.57754, 23.33659, 23.09244, 22.84524, 
    22.59513, 22.34225, 22.08672, 21.82868, 21.56826, 21.30557,
  22.04024, 22.31014, 22.57764, 22.84263, 23.10497, 23.36455, 23.6212, 
    23.87482, 24.12524, 24.37232, 24.61593, 24.85591, 25.0921, 25.32435, 
    25.55252, 25.77643, 25.99593, 26.21087, 26.42107, 26.62638, 26.82663, 
    27.02167, 27.21133, 27.39545, 27.57387, 27.74643, 27.91298, 28.07337, 
    28.22743, 28.37503, 28.51603, 28.65027, 28.77763, 28.89797, 29.01118, 
    29.11712, 29.2157, 29.3068, 29.39032, 29.46618, 29.53428, 29.59455, 
    29.64693, 29.69135, 29.72776, 29.75613, 29.77641, 29.78859, 29.79265, 
    29.78859, 29.77641, 29.75613, 29.72776, 29.69135, 29.64693, 29.59455, 
    29.53428, 29.46618, 29.39032, 29.3068, 29.2157, 29.11712, 29.01118, 
    28.89797, 28.77763, 28.65027, 28.51603, 28.37503, 28.22743, 28.07337, 
    27.91298, 27.74643, 27.57387, 27.39545, 27.21133, 27.02167, 26.82663, 
    26.62638, 26.42107, 26.21087, 25.99593, 25.77643, 25.55252, 25.32435, 
    25.0921, 24.85591, 24.61593, 24.37232, 24.12524, 23.87482, 23.6212, 
    23.36455, 23.10497, 22.84263, 22.57764, 22.31014, 22.04024,
  22.77492, 23.05183, 23.32623, 23.59798, 23.86696, 24.13302, 24.39604, 
    24.65587, 24.91236, 25.16539, 25.41478, 25.6604, 25.9021, 26.13971, 
    26.37307, 26.60204, 26.82645, 27.04614, 27.26094, 27.47071, 27.67526, 
    27.87444, 28.06809, 28.25605, 28.43815, 28.61425, 28.78417, 28.94778, 
    29.10491, 29.25543, 29.39919, 29.53604, 29.66586, 29.78851, 29.90387, 
    30.01182, 30.11224, 30.20505, 30.29012, 30.36738, 30.43673, 30.49811, 
    30.55145, 30.59668, 30.63375, 30.66263, 30.68328, 30.69568, 30.69982, 
    30.69568, 30.68328, 30.66263, 30.63375, 30.59668, 30.55145, 30.49811, 
    30.43673, 30.36738, 30.29012, 30.20505, 30.11224, 30.01182, 29.90387, 
    29.78851, 29.66586, 29.53604, 29.39919, 29.25543, 29.10491, 28.94778, 
    28.78417, 28.61425, 28.43815, 28.25605, 28.06809, 27.87444, 27.67526, 
    27.47071, 27.26094, 27.04614, 26.82645, 26.60204, 26.37307, 26.13971, 
    25.9021, 25.6604, 25.41478, 25.16539, 24.91236, 24.65587, 24.39604, 
    24.13302, 23.86696, 23.59798, 23.32623, 23.05183, 22.77492,
  23.50959, 23.79335, 24.07445, 24.35277, 24.62818, 24.90054, 25.16972, 
    25.43556, 25.69794, 25.95669, 26.21167, 26.46273, 26.70972, 26.95247, 
    27.19084, 27.42466, 27.65377, 27.87801, 28.09721, 28.31122, 28.51988, 
    28.72301, 28.92046, 29.11207, 29.29767, 29.47712, 29.65025, 29.8169, 
    29.97694, 30.13022, 30.27658, 30.4159, 30.54803, 30.67286, 30.79025, 
    30.90008, 31.00225, 31.09665, 31.18319, 31.26176, 31.33229, 31.39471, 
    31.44894, 31.49493, 31.53263, 31.56199, 31.58298, 31.59559, 31.59979, 
    31.59559, 31.58298, 31.56199, 31.53263, 31.49493, 31.44894, 31.39471, 
    31.33229, 31.26176, 31.18319, 31.09665, 31.00225, 30.90008, 30.79025, 
    30.67286, 30.54803, 30.4159, 30.27658, 30.13022, 29.97694, 29.8169, 
    29.65025, 29.47712, 29.29767, 29.11207, 28.92046, 28.72301, 28.51988, 
    28.31122, 28.09721, 27.87801, 27.65377, 27.42466, 27.19084, 26.95247, 
    26.70972, 26.46273, 26.21167, 25.95669, 25.69794, 25.43556, 25.16972, 
    24.90054, 24.62818, 24.35277, 24.07445, 23.79335, 23.50959,
  24.24427, 24.53467, 24.82229, 25.10699, 25.38863, 25.66709, 25.94222, 
    26.21387, 26.48191, 26.74619, 27.00655, 27.26284, 27.51491, 27.76261, 
    28.00576, 28.24422, 28.47782, 28.70641, 28.92981, 29.14787, 29.36043, 
    29.56732, 29.76838, 29.96344, 30.15236, 30.33498, 30.51114, 30.68068, 
    30.84346, 30.99933, 31.14815, 31.28979, 31.4241, 31.55096, 31.67025, 
    31.78186, 31.88566, 31.98156, 32.06945, 32.14926, 32.22089, 32.28428, 
    32.33934, 32.38604, 32.42432, 32.45413, 32.47544, 32.48825, 32.49251, 
    32.48825, 32.47544, 32.45413, 32.42432, 32.38604, 32.33934, 32.28428, 
    32.22089, 32.14926, 32.06945, 31.98156, 31.88566, 31.78186, 31.67025, 
    31.55096, 31.4241, 31.28979, 31.14815, 30.99933, 30.84346, 30.68068, 
    30.51114, 30.33498, 30.15236, 29.96344, 29.76838, 29.56732, 29.36043, 
    29.14787, 28.92981, 28.70641, 28.47782, 28.24422, 28.00576, 27.76261, 
    27.51491, 27.26284, 27.00655, 26.74619, 26.48191, 26.21387, 25.94222, 
    25.66709, 25.38863, 25.10699, 24.82229, 24.53467, 24.24427,
  24.97894, 25.2758, 25.56974, 25.86061, 26.14829, 26.43264, 26.71351, 
    26.99077, 27.26427, 27.53386, 27.79938, 28.0607, 28.31764, 28.57006, 
    28.81779, 29.06068, 29.29857, 29.5313, 29.75869, 29.9806, 30.19686, 
    30.4073, 30.61178, 30.81012, 31.00217, 31.18778, 31.36679, 31.53904, 
    31.7044, 31.86271, 32.01384, 32.15764, 32.29399, 32.42276, 32.54383, 
    32.65709, 32.76241, 32.85971, 32.94887, 33.02983, 33.10248, 33.16676, 
    33.22261, 33.26997, 33.30878, 33.33901, 33.36062, 33.3736, 33.37793, 
    33.3736, 33.36062, 33.33901, 33.30878, 33.26997, 33.22261, 33.16676, 
    33.10248, 33.02983, 32.94887, 32.85971, 32.76241, 32.65709, 32.54383, 
    32.42276, 32.29399, 32.15764, 32.01384, 31.86271, 31.7044, 31.53904, 
    31.36679, 31.18778, 31.00217, 30.81012, 30.61178, 30.4073, 30.19686, 
    29.9806, 29.75869, 29.5313, 29.29857, 29.06068, 28.81779, 28.57006, 
    28.31764, 28.0607, 27.79938, 27.53386, 27.26427, 26.99077, 26.71351, 
    26.43264, 26.14829, 25.86061, 25.56974, 25.2758, 24.97894,
  25.71362, 26.01674, 26.31679, 26.61363, 26.90714, 27.19717, 27.48358, 
    27.76624, 28.04498, 28.31966, 28.59014, 28.85626, 29.11786, 29.37479, 
    29.62689, 29.874, 30.11596, 30.35262, 30.5838, 30.80936, 31.02912, 
    31.24292, 31.45062, 31.65205, 31.84704, 32.03546, 32.21714, 32.39194, 
    32.55971, 32.7203, 32.87358, 33.01942, 33.15767, 33.28822, 33.41094, 
    33.52573, 33.63246, 33.73105, 33.8214, 33.90341, 33.97701, 34.04213, 
    34.0987, 34.14666, 34.18597, 34.21658, 34.23848, 34.25162, 34.256, 
    34.25162, 34.23848, 34.21658, 34.18597, 34.14666, 34.0987, 34.04213, 
    33.97701, 33.90341, 33.8214, 33.73105, 33.63246, 33.52573, 33.41094, 
    33.28822, 33.15767, 33.01942, 32.87358, 32.7203, 32.55971, 32.39194, 
    32.21714, 32.03546, 31.84704, 31.65205, 31.45062, 31.24292, 31.02912, 
    30.80936, 30.5838, 30.35262, 30.11596, 29.874, 29.62689, 29.37479, 
    29.11786, 28.85626, 28.59014, 28.31966, 28.04498, 27.76624, 27.48358, 
    27.19717, 26.90714, 26.61363, 26.31679, 26.01674, 25.71362,
  26.44829, 26.75747, 27.06343, 27.36604, 27.66517, 27.96067, 28.25241, 
    28.54023, 28.82401, 29.10357, 29.37879, 29.64949, 29.91554, 30.17676, 
    30.43301, 30.68413, 30.92996, 31.17034, 31.4051, 31.63409, 31.85715, 
    32.07413, 32.28485, 32.48917, 32.68693, 32.87798, 33.06216, 33.23934, 
    33.40936, 33.57207, 33.72735, 33.87507, 34.01508, 34.14728, 34.27153, 
    34.38773, 34.49578, 34.59556, 34.68699, 34.76999, 34.84446, 34.91034, 
    34.96757, 35.01609, 35.05586, 35.08683, 35.10897, 35.12226, 35.12669, 
    35.12226, 35.10897, 35.08683, 35.05586, 35.01609, 34.96757, 34.91034, 
    34.84446, 34.76999, 34.68699, 34.59556, 34.49578, 34.38773, 34.27153, 
    34.14728, 34.01508, 33.87507, 33.72735, 33.57207, 33.40936, 33.23934, 
    33.06216, 32.87798, 32.68693, 32.48917, 32.28485, 32.07413, 31.85715, 
    31.63409, 31.4051, 31.17034, 30.92996, 30.68413, 30.43301, 30.17676, 
    29.91554, 29.64949, 29.37879, 29.10357, 28.82401, 28.54023, 28.25241, 
    27.96067, 27.66517, 27.36604, 27.06343, 26.75747, 26.44829,
  27.18297, 27.49799, 27.80966, 28.11782, 28.42235, 28.72311, 29.01996, 
    29.31275, 29.60133, 29.88556, 30.16529, 30.44036, 30.71063, 30.97594, 
    31.23613, 31.49104, 31.74052, 31.98441, 32.22254, 32.45477, 32.68093, 
    32.90088, 33.11443, 33.32146, 33.5218, 33.7153, 33.90181, 34.08119, 
    34.25329, 34.41798, 34.57511, 34.72456, 34.8662, 34.99992, 35.12558, 
    35.24308, 35.35233, 35.45321, 35.54563, 35.62952, 35.70479, 35.77137, 
    35.8292, 35.87823, 35.91842, 35.94971, 35.97208, 35.98551, 35.98999, 
    35.98551, 35.97208, 35.94971, 35.91842, 35.87823, 35.8292, 35.77137, 
    35.70479, 35.62952, 35.54563, 35.45321, 35.35233, 35.24308, 35.12558, 
    34.99992, 34.8662, 34.72456, 34.57511, 34.41798, 34.25329, 34.08119, 
    33.90181, 33.7153, 33.5218, 33.32146, 33.11443, 32.90088, 32.68093, 
    32.45477, 32.22254, 31.98441, 31.74052, 31.49104, 31.23613, 30.97594, 
    30.71063, 30.44036, 30.16529, 29.88556, 29.60133, 29.31275, 29.01996, 
    28.72311, 28.42235, 28.11782, 27.80966, 27.49799, 27.18297,
  27.91764, 28.23831, 28.55546, 28.86897, 29.17869, 29.48449, 29.78622, 
    30.08375, 30.37692, 30.6656, 30.94962, 31.22885, 31.50312, 31.77229, 
    32.03619, 32.29469, 32.5476, 32.79479, 33.03609, 33.27135, 33.50042, 
    33.72313, 33.93933, 34.14888, 34.35161, 34.54738, 34.73605, 34.91746, 
    35.09149, 35.25799, 35.41682, 35.56787, 35.71101, 35.8461, 35.97306, 
    36.09175, 36.20208, 36.30396, 36.39729, 36.48199, 36.55799, 36.62521, 
    36.68359, 36.73308, 36.77364, 36.80522, 36.8278, 36.84136, 36.84588, 
    36.84136, 36.8278, 36.80522, 36.77364, 36.73308, 36.68359, 36.62521, 
    36.55799, 36.48199, 36.39729, 36.30396, 36.20208, 36.09175, 35.97306, 
    35.8461, 35.71101, 35.56787, 35.41682, 35.25799, 35.09149, 34.91746, 
    34.73605, 34.54738, 34.35161, 34.14888, 33.93933, 33.72313, 33.50042, 
    33.27135, 33.03609, 32.79479, 32.5476, 32.29469, 32.03619, 31.77229, 
    31.50312, 31.22885, 30.94962, 30.6656, 30.37692, 30.08375, 29.78622, 
    29.48449, 29.17869, 28.86897, 28.55546, 28.23831, 27.91764,
  28.65232, 28.97841, 29.30084, 29.61947, 29.93416, 30.24478, 30.55118, 
    30.85322, 31.15076, 31.44366, 31.73176, 32.01491, 32.29297, 32.56578, 
    32.83318, 33.09504, 33.35118, 33.60146, 33.84572, 34.08381, 34.31557, 
    34.54086, 34.75951, 34.97139, 35.17633, 35.3742, 35.56485, 35.74813, 
    35.92393, 36.09208, 36.25248, 36.40498, 36.54947, 36.68583, 36.81395, 
    36.93372, 37.04504, 37.14782, 37.24197, 37.3274, 37.40405, 37.47184, 
    37.53071, 37.58062, 37.62151, 37.65335, 37.67612, 37.68979, 37.69435, 
    37.68979, 37.67612, 37.65335, 37.62151, 37.58062, 37.53071, 37.47184, 
    37.40405, 37.3274, 37.24197, 37.14782, 37.04504, 36.93372, 36.81395, 
    36.68583, 36.54947, 36.40498, 36.25248, 36.09208, 35.92393, 35.74813, 
    35.56485, 35.3742, 35.17633, 34.97139, 34.75951, 34.54086, 34.31557, 
    34.08381, 33.84572, 33.60146, 33.35118, 33.09504, 32.83318, 32.56578, 
    32.29297, 32.01491, 31.73176, 31.44366, 31.15076, 30.85322, 30.55118, 
    30.24478, 29.93416, 29.61947, 29.30084, 28.97841, 28.65232,
  29.38699, 29.7183, 30.04578, 30.36931, 30.68875, 31.00396, 31.31481, 
    31.62114, 31.92283, 32.21972, 32.51167, 32.79853, 33.08015, 33.35638, 
    33.62707, 33.89207, 34.15122, 34.40438, 34.6514, 34.89211, 35.12637, 
    35.35404, 35.57495, 35.78897, 35.99594, 36.19573, 36.38819, 36.57319, 
    36.75058, 36.92025, 37.08205, 37.23587, 37.38158, 37.51908, 37.64825, 
    37.76899, 37.8812, 37.98478, 38.07965, 38.16574, 38.24297, 38.31126, 
    38.37057, 38.42085, 38.46204, 38.49412, 38.51705, 38.53082, 38.53541, 
    38.53082, 38.51705, 38.49412, 38.46204, 38.42085, 38.37057, 38.31126, 
    38.24297, 38.16574, 38.07965, 37.98478, 37.8812, 37.76899, 37.64825, 
    37.51908, 37.38158, 37.23587, 37.08205, 36.92025, 36.75058, 36.57319, 
    36.38819, 36.19573, 35.99594, 35.78897, 35.57495, 35.35404, 35.12637, 
    34.89211, 34.6514, 34.40438, 34.15122, 33.89207, 33.62707, 33.35638, 
    33.08015, 32.79853, 32.51167, 32.21972, 31.92283, 31.62114, 31.31481, 
    31.00396, 30.68875, 30.36931, 30.04578, 29.7183, 29.38699,
  30.12167, 30.45796, 30.79028, 31.11849, 31.44245, 31.76203, 32.0771, 
    32.3875, 32.6931, 32.99376, 33.28933, 33.57967, 33.86464, 34.14407, 
    34.41782, 34.68575, 34.94771, 35.20354, 35.45309, 35.69623, 35.9328, 
    36.16264, 36.38563, 36.6016, 36.81043, 37.01196, 37.20607, 37.39261, 
    37.57145, 37.74247, 37.90554, 38.06054, 38.20735, 38.34586, 38.47596, 
    38.59755, 38.71054, 38.81484, 38.91036, 38.99702, 39.07475, 39.1435, 
    39.20319, 39.25378, 39.29524, 39.32752, 39.3506, 39.36445, 39.36907, 
    39.36445, 39.3506, 39.32752, 39.29524, 39.25378, 39.20319, 39.1435, 
    39.07475, 38.99702, 38.91036, 38.81484, 38.71054, 38.59755, 38.47596, 
    38.34586, 38.20735, 38.06054, 37.90554, 37.74247, 37.57145, 37.39261, 
    37.20607, 37.01196, 36.81043, 36.6016, 36.38563, 36.16264, 35.9328, 
    35.69623, 35.45309, 35.20354, 34.94771, 34.68575, 34.41782, 34.14407, 
    33.86464, 33.57967, 33.28933, 32.99376, 32.6931, 32.3875, 32.0771, 
    31.76203, 31.44245, 31.11849, 30.79028, 30.45796, 30.12167,
  30.85634, 31.19741, 31.53433, 31.86699, 32.19525, 32.51897, 32.83802, 
    33.15226, 33.46156, 33.76576, 34.06473, 34.35833, 34.64641, 34.92882, 
    35.20542, 35.47607, 35.74061, 35.9989, 36.2508, 36.49615, 36.73482, 
    36.96666, 37.19153, 37.40928, 37.61977, 37.82288, 38.01846, 38.20639, 
    38.38652, 38.55875, 38.72294, 38.87898, 39.02676, 39.16616, 39.29708, 
    39.41943, 39.5331, 39.63801, 39.73409, 39.82125, 39.89942, 39.96855, 
    40.02857, 40.07944, 40.12112, 40.15358, 40.17678, 40.1907, 40.19535, 
    40.1907, 40.17678, 40.15358, 40.12112, 40.07944, 40.02857, 39.96855, 
    39.89942, 39.82125, 39.73409, 39.63801, 39.5331, 39.41943, 39.29708, 
    39.16616, 39.02676, 38.87898, 38.72294, 38.55875, 38.38652, 38.20639, 
    38.01846, 37.82288, 37.61977, 37.40928, 37.19153, 36.96666, 36.73482, 
    36.49615, 36.2508, 35.9989, 35.74061, 35.47607, 35.20542, 34.92882, 
    34.64641, 34.35833, 34.06473, 33.76576, 33.46156, 33.15226, 32.83802, 
    32.51897, 32.19525, 31.86699, 31.53433, 31.19741, 30.85634,
  31.59101, 31.93662, 32.27793, 32.61481, 32.94714, 33.27477, 33.59758, 
    33.91543, 34.22818, 34.5357, 34.83784, 35.13448, 35.42545, 35.71062, 
    35.98985, 36.26299, 36.52991, 36.79046, 37.04449, 37.29186, 37.53244, 
    37.76608, 37.99264, 38.21198, 38.42397, 38.62848, 38.82537, 39.01452, 
    39.1958, 39.36908, 39.53426, 39.69121, 39.83982, 39.97999, 40.11162, 
    40.23461, 40.34887, 40.45432, 40.55087, 40.63845, 40.717, 40.78645, 
    40.84675, 40.89785, 40.93972, 40.97232, 40.99562, 41.00961, 41.01428, 
    41.00961, 40.99562, 40.97232, 40.93972, 40.89785, 40.84675, 40.78645, 
    40.717, 40.63845, 40.55087, 40.45432, 40.34887, 40.23461, 40.11162, 
    39.97999, 39.83982, 39.69121, 39.53426, 39.36908, 39.1958, 39.01452, 
    38.82537, 38.62848, 38.42397, 38.21198, 37.99264, 37.76608, 37.53244, 
    37.29186, 37.04449, 36.79046, 36.52991, 36.26299, 35.98985, 35.71062, 
    35.42545, 35.13448, 34.83784, 34.5357, 34.22818, 33.91543, 33.59758, 
    33.27477, 32.94714, 32.61481, 32.27793, 31.93662, 31.59101,
  32.32569, 32.67561, 33.02107, 33.36194, 33.6981, 34.02942, 34.35575, 
    34.67698, 34.99296, 35.30357, 35.60866, 35.90809, 36.20173, 36.48944, 
    36.77109, 37.04652, 37.3156, 37.57819, 37.83415, 38.08334, 38.32563, 
    38.56088, 38.78895, 39.00971, 39.22302, 39.42876, 39.6268, 39.81702, 
    39.99928, 40.17348, 40.3395, 40.49723, 40.64656, 40.78738, 40.91961, 
    41.04314, 41.15789, 41.26377, 41.36071, 41.44865, 41.5275, 41.59722, 
    41.65775, 41.70904, 41.75106, 41.78378, 41.80717, 41.82121, 41.82589, 
    41.82121, 41.80717, 41.78378, 41.75106, 41.70904, 41.65775, 41.59722, 
    41.5275, 41.44865, 41.36071, 41.26377, 41.15789, 41.04314, 40.91961, 
    40.78738, 40.64656, 40.49723, 40.3395, 40.17348, 39.99928, 39.81702, 
    39.6268, 39.42876, 39.22302, 39.00971, 38.78895, 38.56088, 38.32563, 
    38.08334, 37.83415, 37.57819, 37.3156, 37.04652, 36.77109, 36.48944, 
    36.20173, 35.90809, 35.60866, 35.30357, 34.99296, 34.67698, 34.35575, 
    34.02942, 33.6981, 33.36194, 33.02107, 32.67561, 32.32569,
  33.06036, 33.41436, 33.76374, 34.10837, 34.44813, 34.78289, 35.11252, 
    35.4369, 35.75588, 36.06934, 36.37715, 36.67916, 36.97525, 37.26529, 
    37.54912, 37.82662, 38.09766, 38.36209, 38.61978, 38.87059, 39.1144, 
    39.35107, 39.58046, 39.80246, 40.01692, 40.22372, 40.42275, 40.61388, 
    40.79699, 40.97196, 41.13869, 41.29707, 41.44698, 41.58834, 41.72106, 
    41.84503, 41.96017, 42.06641, 42.16367, 42.25187, 42.33097, 42.40089, 
    42.4616, 42.51304, 42.55518, 42.58799, 42.61144, 42.62552, 42.63021, 
    42.62552, 42.61144, 42.58799, 42.55518, 42.51304, 42.4616, 42.40089, 
    42.33097, 42.25187, 42.16367, 42.06641, 41.96017, 41.84503, 41.72106, 
    41.58834, 41.44698, 41.29707, 41.13869, 40.97196, 40.79699, 40.61388, 
    40.42275, 40.22372, 40.01692, 39.80246, 39.58046, 39.35107, 39.1144, 
    38.87059, 38.61978, 38.36209, 38.09766, 37.82662, 37.54912, 37.26529, 
    36.97525, 36.67916, 36.37715, 36.06934, 35.75588, 35.4369, 35.11252, 
    34.78289, 34.44813, 34.10837, 33.76374, 33.41436, 33.06036,
  33.79504, 34.15289, 34.50594, 34.8541, 35.19722, 35.53519, 35.86789, 
    36.19517, 36.51693, 36.83301, 37.14331, 37.44768, 37.746, 38.03813, 
    38.32394, 38.6033, 38.87608, 39.14214, 39.40136, 39.6536, 39.89874, 
    40.13664, 40.36718, 40.59023, 40.80568, 41.01338, 41.21324, 41.40512, 
    41.58892, 41.76453, 41.93184, 42.09073, 42.24112, 42.38291, 42.516, 
    42.64032, 42.75576, 42.86227, 42.95976, 43.04817, 43.12745, 43.19752, 
    43.25835, 43.3099, 43.35213, 43.385, 43.4085, 43.4226, 43.42731, 43.4226, 
    43.4085, 43.385, 43.35213, 43.3099, 43.25835, 43.19752, 43.12745, 
    43.04817, 42.95976, 42.86227, 42.75576, 42.64032, 42.516, 42.38291, 
    42.24112, 42.09073, 41.93184, 41.76453, 41.58892, 41.40512, 41.21324, 
    41.01338, 40.80568, 40.59023, 40.36718, 40.13664, 39.89874, 39.6536, 
    39.40136, 39.14214, 38.87608, 38.6033, 38.32394, 38.03813, 37.746, 
    37.44768, 37.14331, 36.83301, 36.51693, 36.19517, 35.86789, 35.53519, 
    35.19722, 34.8541, 34.50594, 34.15289, 33.79504,
  34.52972, 34.89117, 35.24767, 35.59911, 35.94537, 36.28631, 36.62183, 
    36.95179, 37.27608, 37.59457, 37.90713, 38.21363, 38.51395, 38.80796, 
    39.09554, 39.37654, 39.65086, 39.91835, 40.1789, 40.43238, 40.67865, 
    40.9176, 41.14911, 41.37305, 41.5893, 41.79774, 41.99827, 42.19077, 
    42.37512, 42.55122, 42.71897, 42.87827, 43.02901, 43.17111, 43.30448, 
    43.42903, 43.54469, 43.65138, 43.74903, 43.83758, 43.91697, 43.98714, 
    44.04806, 44.09967, 44.14195, 44.17486, 44.19839, 44.21251, 44.21722, 
    44.21251, 44.19839, 44.17486, 44.14195, 44.09967, 44.04806, 43.98714, 
    43.91697, 43.83758, 43.74903, 43.65138, 43.54469, 43.42903, 43.30448, 
    43.17111, 43.02901, 42.87827, 42.71897, 42.55122, 42.37512, 42.19077, 
    41.99827, 41.79774, 41.5893, 41.37305, 41.14911, 40.9176, 40.67865, 
    40.43238, 40.1789, 39.91835, 39.65086, 39.37654, 39.09554, 38.80796, 
    38.51395, 38.21363, 37.90713, 37.59457, 37.27608, 36.95179, 36.62183, 
    36.28631, 35.94537, 35.59911, 35.24767, 34.89117, 34.52972,
  35.26439, 35.62921, 35.98892, 36.34341, 36.69255, 37.03624, 37.37434, 
    37.70675, 38.03334, 38.354, 38.66859, 38.977, 39.27911, 39.57478, 
    39.8639, 40.14635, 40.42199, 40.69072, 40.9524, 41.20691, 41.45414, 
    41.69396, 41.92625, 42.15091, 42.36781, 42.57683, 42.77788, 42.97084, 
    43.1556, 43.33206, 43.50012, 43.65969, 43.81068, 43.95298, 44.08652, 
    44.21122, 44.32701, 44.4338, 44.53154, 44.62016, 44.6996, 44.76982, 
    44.83077, 44.88241, 44.9247, 44.95763, 44.98116, 44.99529, 45, 44.99529, 
    44.98116, 44.95763, 44.9247, 44.88241, 44.83077, 44.76982, 44.6996, 
    44.62016, 44.53154, 44.4338, 44.32701, 44.21122, 44.08652, 43.95298, 
    43.81068, 43.65969, 43.50012, 43.33206, 43.1556, 42.97084, 42.77788, 
    42.57683, 42.36781, 42.15091, 41.92625, 41.69396, 41.45414, 41.20691, 
    40.9524, 40.69072, 40.42199, 40.14635, 39.8639, 39.57478, 39.27911, 
    38.977, 38.66859, 38.354, 38.03334, 37.70675, 37.37434, 37.03624, 
    36.69255, 36.34341, 35.98892, 35.62921, 35.26439 ;

 grid_lont =
  35.39052, 36.17686, 36.97036, 37.77106, 38.57902, 39.39428, 40.21688, 
    41.04685, 41.88421, 42.72898, 43.58115, 44.44075, 45.30774, 46.18213, 
    47.06388, 47.95295, 48.8493, 49.75288, 50.66362, 51.58143, 52.50624, 
    53.43794, 54.37642, 55.32156, 56.27322, 57.23126, 58.19552, 59.16583, 
    60.142, 61.12385, 62.11116, 63.10371, 64.10129, 65.10364, 66.11051, 
    67.12165, 68.13678, 69.15562, 70.17788, 71.20325, 72.23145, 73.26214, 
    74.29501, 75.32973, 76.36598, 77.40342, 78.44171, 79.48051, 80.51949, 
    81.55829, 82.59658, 83.63402, 84.67027, 85.70499, 86.73786, 87.76855, 
    88.79675, 89.82212, 90.84438, 91.86322, 92.87835, 93.88949, 94.89636, 
    95.89871, 96.89629, 97.88884, 98.87615, 99.85799, 100.8342, 101.8045, 
    102.7687, 103.7268, 104.6784, 105.6236, 106.5621, 107.4938, 108.4186, 
    109.3364, 110.2471, 111.1507, 112.0471, 112.9361, 113.8179, 114.6923, 
    115.5592, 116.4188, 117.271, 118.1158, 118.9531, 119.7831, 120.6057, 
    121.421, 122.2289, 123.0296, 123.8231, 124.6095,
  35.39055, 36.17689, 36.97039, 37.77109, 38.57905, 39.39432, 40.21692, 
    41.04689, 41.88424, 42.72901, 43.58118, 44.44078, 45.30777, 46.18216, 
    47.06391, 47.95298, 48.84933, 49.75291, 50.66364, 51.58146, 52.50626, 
    53.43797, 54.37645, 55.32158, 56.27325, 57.23129, 58.19555, 59.16585, 
    60.14202, 61.12387, 62.11118, 63.10373, 64.1013, 65.10365, 66.11053, 
    67.12167, 68.1368, 69.15563, 70.17789, 71.20326, 72.23145, 73.26215, 
    74.29501, 75.32974, 76.36599, 77.40343, 78.44171, 79.48051, 80.51949, 
    81.55829, 82.59657, 83.63401, 84.67026, 85.70499, 86.73785, 87.76855, 
    88.79674, 89.82211, 90.84437, 91.8632, 92.87833, 93.88947, 94.89635, 
    95.8987, 96.89627, 97.88882, 98.87613, 99.85798, 100.8342, 101.8045, 
    102.7687, 103.7268, 104.6784, 105.6236, 106.562, 107.4937, 108.4185, 
    109.3364, 110.2471, 111.1507, 112.047, 112.9361, 113.8178, 114.6922, 
    115.5592, 116.4188, 117.271, 118.1158, 118.9531, 119.7831, 120.6057, 
    121.4209, 122.2289, 123.0296, 123.8231, 124.6095,
  35.39058, 36.17692, 36.97042, 37.77112, 38.57908, 39.39435, 40.21695, 
    41.04692, 41.88427, 42.72904, 43.58121, 44.44081, 45.3078, 46.18219, 
    47.06393, 47.95301, 48.84936, 49.75294, 50.66367, 51.58149, 52.50629, 
    53.43799, 54.37647, 55.32161, 56.27327, 57.23131, 58.19557, 59.16587, 
    60.14204, 61.12389, 62.11119, 63.10375, 64.10132, 65.10367, 66.11054, 
    67.12168, 68.1368, 69.15564, 70.1779, 71.20328, 72.23147, 73.26215, 
    74.29502, 75.32975, 76.36599, 77.40343, 78.44172, 79.48051, 80.51949, 
    81.55828, 82.59657, 83.63401, 84.67025, 85.70498, 86.73785, 87.76853, 
    88.79672, 89.8221, 90.84436, 91.8632, 92.87832, 93.88946, 94.89633, 
    95.89868, 96.89625, 97.8888, 98.87611, 99.85796, 100.8341, 101.8044, 
    102.7687, 103.7267, 104.6784, 105.6235, 106.562, 107.4937, 108.4185, 
    109.3363, 110.2471, 111.1506, 112.047, 112.9361, 113.8178, 114.6922, 
    115.5592, 116.4188, 117.271, 118.1157, 118.9531, 119.7831, 120.6057, 
    121.4209, 122.2289, 123.0296, 123.8231, 124.6094,
  35.39061, 36.17695, 36.97045, 37.77115, 38.57912, 39.39438, 40.21698, 
    41.04695, 41.8843, 42.72907, 43.58125, 44.44084, 45.30783, 46.18222, 
    47.06396, 47.95304, 48.84939, 49.75296, 50.6637, 51.58151, 52.50632, 
    53.43801, 54.3765, 55.32163, 56.27329, 57.23133, 58.19559, 59.16589, 
    60.14207, 61.12391, 62.11121, 63.10377, 64.10134, 65.10368, 66.11056, 
    67.1217, 68.13682, 69.15565, 70.17791, 71.20329, 72.23148, 73.26216, 
    74.29503, 75.32975, 76.366, 77.40343, 78.44172, 79.48051, 80.51949, 
    81.55828, 82.59657, 83.634, 84.67025, 85.70497, 86.73784, 87.76852, 
    88.79671, 89.82209, 90.84435, 91.86318, 92.8783, 93.88944, 94.89632, 
    95.89866, 96.89623, 97.88879, 98.87609, 99.85793, 100.8341, 101.8044, 
    102.7687, 103.7267, 104.6784, 105.6235, 106.562, 107.4937, 108.4185, 
    109.3363, 110.247, 111.1506, 112.047, 112.936, 113.8178, 114.6922, 
    115.5592, 116.4188, 117.2709, 118.1157, 118.9531, 119.783, 120.6056, 
    121.4209, 122.2288, 123.0295, 123.823, 124.6094,
  35.39064, 36.17699, 36.97048, 37.77118, 38.57915, 39.39441, 40.21701, 
    41.04698, 41.88433, 42.7291, 43.58128, 44.44087, 45.30787, 46.18225, 
    47.064, 47.95307, 48.84942, 49.75299, 50.66373, 51.58154, 52.50634, 
    53.43804, 54.37652, 55.32166, 56.27332, 57.23135, 58.19561, 59.16592, 
    60.14209, 61.12393, 62.11123, 63.10379, 64.10136, 65.1037, 66.11057, 
    67.1217, 68.13683, 69.15567, 70.17793, 71.20329, 72.23148, 73.26217, 
    74.29504, 75.32976, 76.366, 77.40343, 78.44172, 79.48051, 80.51949, 
    81.55828, 82.59657, 83.634, 84.67024, 85.70496, 86.73783, 87.76852, 
    88.79671, 89.82207, 90.84433, 91.86317, 92.8783, 93.88943, 94.8963, 
    95.89864, 96.89622, 97.88876, 98.87608, 99.85791, 100.8341, 101.8044, 
    102.7686, 103.7267, 104.6783, 105.6235, 106.562, 107.4937, 108.4185, 
    109.3363, 110.247, 111.1506, 112.0469, 112.936, 113.8177, 114.6921, 
    115.5591, 116.4187, 117.2709, 118.1157, 118.953, 119.783, 120.6056, 
    121.4209, 122.2288, 123.0295, 123.823, 124.6094,
  35.39067, 36.17702, 36.97051, 37.77121, 38.57918, 39.39444, 40.21704, 
    41.04701, 41.88437, 42.72913, 43.58131, 44.4409, 45.30789, 46.18228, 
    47.06402, 47.95309, 48.84945, 49.75302, 50.66375, 51.58157, 52.50637, 
    53.43807, 54.37654, 55.32168, 56.27334, 57.23138, 58.19563, 59.16594, 
    60.14211, 61.12395, 62.11125, 63.10381, 64.10137, 65.10372, 66.11059, 
    67.12172, 68.13685, 69.15568, 70.17793, 71.20331, 72.23149, 73.26218, 
    74.29504, 75.32977, 76.366, 77.40343, 78.44172, 79.48051, 80.51949, 
    81.55828, 82.59657, 83.634, 84.67023, 85.70496, 86.73782, 87.76851, 
    88.79669, 89.82207, 90.84432, 91.86315, 92.87828, 93.88941, 94.89628, 
    95.89863, 96.89619, 97.88875, 98.87605, 99.85789, 100.8341, 101.8044, 
    102.7686, 103.7267, 104.6783, 105.6235, 106.5619, 107.4936, 108.4184, 
    109.3362, 110.247, 111.1506, 112.0469, 112.936, 113.8177, 114.6921, 
    115.5591, 116.4187, 117.2709, 118.1156, 118.953, 119.783, 120.6056, 
    121.4208, 122.2288, 123.0295, 123.823, 124.6093,
  35.39071, 36.17704, 36.97054, 37.77124, 38.57921, 39.39447, 40.21707, 
    41.04704, 41.8844, 42.72916, 43.58134, 44.44093, 45.30792, 46.1823, 
    47.06405, 47.95312, 48.84948, 49.75305, 50.66378, 51.58159, 52.5064, 
    53.43809, 54.37657, 55.3217, 56.27337, 57.2314, 58.19566, 59.16596, 
    60.14213, 61.12397, 62.11127, 63.10382, 64.10139, 65.10374, 66.1106, 
    67.12173, 68.13686, 69.15569, 70.17794, 71.20332, 72.2315, 73.26218, 
    74.29505, 75.32977, 76.36601, 77.40344, 78.44173, 79.48051, 80.51949, 
    81.55827, 82.59656, 83.63399, 84.67023, 85.70495, 86.73782, 87.7685, 
    88.79668, 89.82206, 90.84431, 91.86314, 92.87827, 93.8894, 94.89626, 
    95.89861, 96.89618, 97.88873, 98.87603, 99.85787, 100.834, 101.8043, 
    102.7686, 103.7266, 104.6783, 105.6234, 106.5619, 107.4936, 108.4184, 
    109.3362, 110.2469, 111.1505, 112.0469, 112.936, 113.8177, 114.6921, 
    115.5591, 116.4187, 117.2708, 118.1156, 118.953, 119.7829, 120.6055, 
    121.4208, 122.2288, 123.0295, 123.823, 124.6093,
  35.39074, 36.17707, 36.97057, 37.77127, 38.57924, 39.3945, 40.2171, 
    41.04707, 41.88443, 42.72919, 43.58136, 44.44096, 45.30795, 46.18233, 
    47.06408, 47.95315, 48.8495, 49.75307, 50.66381, 51.58162, 52.50642, 
    53.43812, 54.37659, 55.32173, 56.27339, 57.23142, 58.19568, 59.16598, 
    60.14215, 61.12399, 62.11129, 63.10384, 64.10141, 65.10375, 66.11062, 
    67.12175, 68.13687, 69.1557, 70.17796, 71.20332, 72.23151, 73.26219, 
    74.29506, 75.32977, 76.36601, 77.40344, 78.44173, 79.48051, 80.51949, 
    81.55827, 82.59656, 83.63399, 84.67023, 85.70494, 86.73781, 87.76849, 
    88.79668, 89.82204, 90.8443, 91.86313, 92.87825, 93.88938, 94.89625, 
    95.89859, 96.89616, 97.88871, 98.87601, 99.85785, 100.834, 101.8043, 
    102.7686, 103.7266, 104.6783, 105.6234, 106.5619, 107.4936, 108.4184, 
    109.3362, 110.2469, 111.1505, 112.0469, 112.9359, 113.8177, 114.692, 
    115.559, 116.4186, 117.2708, 118.1156, 118.9529, 119.7829, 120.6055, 
    121.4208, 122.2287, 123.0294, 123.8229, 124.6093,
  35.39077, 36.1771, 36.9706, 37.77131, 38.57927, 39.39453, 40.21713, 
    41.0471, 41.88445, 42.72922, 43.58139, 44.44098, 45.30798, 46.18237, 
    47.06411, 47.95318, 48.84953, 49.75311, 50.66383, 51.58165, 52.50645, 
    53.43814, 54.37662, 55.32175, 56.27341, 57.23145, 58.1957, 59.166, 
    60.14217, 61.12401, 62.11131, 63.10386, 64.10143, 65.10377, 66.11063, 
    67.12177, 68.13689, 69.15572, 70.17796, 71.20334, 72.23152, 73.2622, 
    74.29506, 75.32978, 76.36602, 77.40345, 78.44173, 79.48052, 80.51948, 
    81.55827, 82.59655, 83.63398, 84.67022, 85.70494, 86.7378, 87.76848, 
    88.79666, 89.82204, 90.84428, 91.86311, 92.87823, 93.88937, 94.89623, 
    95.89857, 96.89614, 97.88869, 98.87599, 99.85783, 100.834, 101.8043, 
    102.7686, 103.7266, 104.6782, 105.6234, 106.5619, 107.4936, 108.4184, 
    109.3362, 110.2469, 111.1505, 112.0468, 112.9359, 113.8176, 114.692, 
    115.559, 116.4186, 117.2708, 118.1155, 118.9529, 119.7829, 120.6055, 
    121.4207, 122.2287, 123.0294, 123.8229, 124.6092,
  35.39079, 36.17713, 36.97063, 37.77133, 38.5793, 39.39456, 40.21716, 
    41.04713, 41.88448, 42.72924, 43.58142, 44.44101, 45.30801, 46.18239, 
    47.06414, 47.95321, 48.84956, 49.75313, 50.66386, 51.58167, 52.50647, 
    53.43817, 54.37664, 55.32178, 56.27344, 57.23147, 58.19572, 59.16602, 
    60.14219, 61.12403, 62.11133, 63.10388, 64.10144, 65.10378, 66.11065, 
    67.12178, 68.1369, 69.15573, 70.17798, 71.20335, 72.23153, 73.26221, 
    74.29507, 75.32978, 76.36602, 77.40345, 78.44173, 79.48052, 80.51948, 
    81.55827, 82.59655, 83.63398, 84.67022, 85.70493, 86.73779, 87.76847, 
    88.79665, 89.82202, 90.84427, 91.8631, 92.87822, 93.88935, 94.89622, 
    95.89856, 96.89613, 97.88867, 98.87597, 99.85781, 100.834, 101.8043, 
    102.7685, 103.7266, 104.6782, 105.6234, 106.5618, 107.4935, 108.4183, 
    109.3361, 110.2469, 111.1504, 112.0468, 112.9359, 113.8176, 114.692, 
    115.559, 116.4186, 117.2708, 118.1155, 118.9529, 119.7828, 120.6054, 
    121.4207, 122.2287, 123.0294, 123.8229, 124.6092,
  35.39082, 36.17716, 36.97066, 37.77136, 38.57932, 39.39459, 40.21719, 
    41.04715, 41.88451, 42.72927, 43.58145, 44.44104, 45.30804, 46.18242, 
    47.06416, 47.95324, 48.84959, 49.75316, 50.66389, 51.5817, 52.5065, 
    53.43819, 54.37667, 55.3218, 56.27346, 57.23149, 58.19575, 59.16605, 
    60.14221, 61.12405, 62.11135, 63.1039, 64.10146, 65.1038, 66.11066, 
    67.1218, 68.13691, 69.15574, 70.17799, 71.20335, 72.23154, 73.26221, 
    74.29507, 75.32979, 76.36603, 77.40345, 78.44173, 79.48052, 80.51948, 
    81.55827, 82.59655, 83.63397, 84.67021, 85.70493, 86.73779, 87.76846, 
    88.79665, 89.82201, 90.84426, 91.86309, 92.8782, 93.88934, 94.8962, 
    95.89854, 96.8961, 97.88865, 98.87595, 99.85779, 100.834, 101.8043, 
    102.7685, 103.7265, 104.6782, 105.6233, 106.5618, 107.4935, 108.4183, 
    109.3361, 110.2468, 111.1504, 112.0468, 112.9358, 113.8176, 114.692, 
    115.559, 116.4185, 117.2707, 118.1155, 118.9528, 119.7828, 120.6054, 
    121.4207, 122.2286, 123.0293, 123.8228, 124.6092,
  35.39085, 36.17719, 36.97068, 37.77139, 38.57935, 39.39462, 40.21722, 
    41.04718, 41.88454, 42.7293, 43.58148, 44.44107, 45.30806, 46.18245, 
    47.06419, 47.95326, 48.84961, 49.75319, 50.66391, 51.58173, 52.50653, 
    53.43822, 54.37669, 55.32183, 56.27348, 57.23152, 58.19577, 59.16607, 
    60.14223, 61.12407, 62.11137, 63.10391, 64.10148, 65.10381, 66.11068, 
    67.12181, 68.13692, 69.15575, 70.178, 71.20337, 72.23154, 73.26222, 
    74.29508, 75.3298, 76.36603, 77.40346, 78.44173, 79.48052, 80.51948, 
    81.55827, 82.59654, 83.63397, 84.6702, 85.70492, 86.73778, 87.76846, 
    88.79663, 89.822, 90.84425, 91.86308, 92.87819, 93.88932, 94.89619, 
    95.89852, 96.89609, 97.88863, 98.87593, 99.85777, 100.8339, 101.8042, 
    102.7685, 103.7265, 104.6782, 105.6233, 106.5618, 107.4935, 108.4183, 
    109.3361, 110.2468, 111.1504, 112.0467, 112.9358, 113.8176, 114.6919, 
    115.5589, 116.4185, 117.2707, 118.1155, 118.9528, 119.7828, 120.6054, 
    121.4206, 122.2286, 123.0293, 123.8228, 124.6092,
  35.39088, 36.17722, 36.97071, 37.77142, 38.57938, 39.39464, 40.21724, 
    41.04721, 41.88457, 42.72933, 43.58151, 44.4411, 45.30809, 46.18248, 
    47.06422, 47.95329, 48.84964, 49.75321, 50.66394, 51.58175, 52.50655, 
    53.43824, 54.37672, 55.32185, 56.27351, 57.23154, 58.19579, 59.16609, 
    60.14225, 61.12409, 62.11139, 63.10393, 64.10149, 65.10384, 66.11069, 
    67.12183, 68.13694, 69.15577, 70.17801, 71.20338, 72.23155, 73.26223, 
    74.29509, 75.3298, 76.36604, 77.40346, 78.44173, 79.48052, 80.51948, 
    81.55827, 82.59654, 83.63396, 84.6702, 85.70491, 86.73777, 87.76845, 
    88.79662, 89.82199, 90.84423, 91.86306, 92.87817, 93.88931, 94.89616, 
    95.89851, 96.89606, 97.88861, 98.87592, 99.85775, 100.8339, 101.8042, 
    102.7685, 103.7265, 104.6781, 105.6233, 106.5618, 107.4934, 108.4183, 
    109.3361, 110.2468, 111.1504, 112.0467, 112.9358, 113.8175, 114.6919, 
    115.5589, 116.4185, 117.2707, 118.1154, 118.9528, 119.7828, 120.6054, 
    121.4206, 122.2286, 123.0293, 123.8228, 124.6091,
  35.3909, 36.17724, 36.97074, 37.77145, 38.57941, 39.39467, 40.21727, 
    41.04724, 41.88459, 42.72936, 43.58154, 44.44112, 45.30812, 46.1825, 
    47.06425, 47.95332, 48.84967, 49.75324, 50.66397, 51.58178, 52.50658, 
    53.43827, 54.37674, 55.32187, 56.27353, 57.23156, 58.19581, 59.16611, 
    60.14227, 61.12411, 62.1114, 63.10395, 64.10151, 65.10385, 66.11071, 
    67.12183, 68.13696, 69.15578, 70.17802, 71.20338, 72.23156, 73.26224, 
    74.2951, 75.3298, 76.36604, 77.40347, 78.44173, 79.48052, 80.51948, 
    81.55827, 82.59653, 83.63396, 84.6702, 85.7049, 86.73776, 87.76844, 
    88.79662, 89.82198, 90.84422, 91.86304, 92.87817, 93.88929, 94.89615, 
    95.89849, 96.89605, 97.8886, 98.87589, 99.85773, 100.8339, 101.8042, 
    102.7684, 103.7265, 104.6781, 105.6233, 106.5617, 107.4934, 108.4182, 
    109.336, 110.2468, 111.1503, 112.0467, 112.9358, 113.8175, 114.6919, 
    115.5589, 116.4185, 117.2706, 118.1154, 118.9528, 119.7827, 120.6053, 
    121.4206, 122.2286, 123.0293, 123.8228, 124.6091,
  35.39093, 36.17727, 36.97076, 37.77147, 38.57943, 39.3947, 40.2173, 
    41.04726, 41.88462, 42.72939, 43.58156, 44.44115, 45.30815, 46.18253, 
    47.06427, 47.95334, 48.84969, 49.75326, 50.66399, 51.5818, 52.5066, 
    53.43829, 54.37677, 55.3219, 56.27355, 57.23158, 58.19584, 59.16613, 
    60.14229, 61.12413, 62.11142, 63.10397, 64.10153, 65.10387, 66.11073, 
    67.12185, 68.13696, 69.15579, 70.17803, 71.20339, 72.23158, 73.26225, 
    74.2951, 75.32981, 76.36604, 77.40347, 78.44173, 79.48052, 80.51948, 
    81.55827, 82.59653, 83.63396, 84.67019, 85.7049, 86.73775, 87.76842, 
    88.79661, 89.82197, 90.84421, 91.86304, 92.87815, 93.88927, 94.89613, 
    95.89847, 96.89603, 97.88857, 98.87587, 99.8577, 100.8339, 101.8042, 
    102.7684, 103.7264, 104.6781, 105.6232, 106.5617, 107.4934, 108.4182, 
    109.336, 110.2467, 111.1503, 112.0467, 112.9357, 113.8175, 114.6919, 
    115.5588, 116.4184, 117.2706, 118.1154, 118.9527, 119.7827, 120.6053, 
    121.4206, 122.2285, 123.0292, 123.8227, 124.6091,
  35.39095, 36.1773, 36.97079, 37.7715, 38.57946, 39.39472, 40.21732, 
    41.04729, 41.88465, 42.72941, 43.58159, 44.44118, 45.30817, 46.18256, 
    47.0643, 47.95337, 48.84972, 49.75329, 50.66402, 51.58183, 52.50663, 
    53.43832, 54.37679, 55.32192, 56.27357, 57.23161, 58.19585, 59.16615, 
    60.14231, 61.12415, 62.11144, 63.10398, 64.10155, 65.10388, 66.11074, 
    67.12186, 68.13698, 69.1558, 70.17805, 71.20341, 72.23158, 73.26225, 
    74.29511, 75.32982, 76.36605, 77.40347, 78.44174, 79.48052, 80.51948, 
    81.55826, 82.59653, 83.63395, 84.67018, 85.70489, 86.73775, 87.76842, 
    88.79659, 89.82195, 90.8442, 91.86302, 92.87814, 93.88926, 94.89612, 
    95.89845, 96.89601, 97.88856, 98.87585, 99.85769, 100.8338, 101.8041, 
    102.7684, 103.7264, 104.6781, 105.6232, 106.5617, 107.4934, 108.4182, 
    109.336, 110.2467, 111.1503, 112.0466, 112.9357, 113.8174, 114.6918, 
    115.5588, 116.4184, 117.2706, 118.1153, 118.9527, 119.7827, 120.6053, 
    121.4205, 122.2285, 123.0292, 123.8227, 124.609,
  35.39098, 36.17732, 36.97082, 37.77152, 38.57949, 39.39475, 40.21735, 
    41.04732, 41.88467, 42.72944, 43.58162, 44.4412, 45.3082, 46.18258, 
    47.06433, 47.9534, 48.84974, 49.75331, 50.66404, 51.58185, 52.50665, 
    53.43834, 54.37682, 55.32195, 56.2736, 57.23163, 58.19588, 59.16617, 
    60.14233, 61.12416, 62.11146, 63.104, 64.10156, 65.1039, 66.11076, 
    67.12188, 68.13699, 69.15582, 70.17805, 71.20341, 72.23159, 73.26226, 
    74.29511, 75.32982, 76.36605, 77.40347, 78.44174, 79.48052, 80.51948, 
    81.55826, 82.59653, 83.63395, 84.67018, 85.70489, 86.73774, 87.76841, 
    88.79659, 89.82195, 90.84418, 91.86301, 92.87812, 93.88924, 94.8961, 
    95.89844, 96.896, 97.88854, 98.87583, 99.85767, 100.8338, 101.8041, 
    102.7684, 103.7264, 104.6781, 105.6232, 106.5617, 107.4933, 108.4182, 
    109.336, 110.2467, 111.1503, 112.0466, 112.9357, 113.8174, 114.6918, 
    115.5588, 116.4184, 117.2706, 118.1153, 118.9527, 119.7826, 120.6052, 
    121.4205, 122.2285, 123.0292, 123.8227, 124.609,
  35.391, 36.17735, 36.97084, 37.77155, 38.57951, 39.39478, 40.21738, 
    41.04734, 41.8847, 42.72947, 43.58164, 44.44123, 45.30822, 46.18261, 
    47.06435, 47.95342, 48.84977, 49.75334, 50.66407, 51.58187, 52.50668, 
    53.43837, 54.37684, 55.32197, 56.27362, 57.23165, 58.1959, 59.16619, 
    60.14235, 61.12418, 62.11148, 63.10402, 64.10158, 65.10391, 66.11077, 
    67.12189, 68.137, 69.15582, 70.17806, 71.20342, 72.2316, 73.26227, 
    74.29512, 75.32983, 76.36606, 77.40347, 78.44174, 79.48052, 80.51948, 
    81.55826, 82.59653, 83.63394, 84.67017, 85.70488, 86.73773, 87.7684, 
    88.79658, 89.82194, 90.84418, 91.863, 92.87811, 93.88923, 94.89609, 
    95.89842, 96.89598, 97.88852, 98.87582, 99.85765, 100.8338, 101.8041, 
    102.7683, 103.7264, 104.678, 105.6232, 106.5616, 107.4933, 108.4181, 
    109.3359, 110.2467, 111.1502, 112.0466, 112.9356, 113.8174, 114.6918, 
    115.5588, 116.4184, 117.2705, 118.1153, 118.9527, 119.7826, 120.6052, 
    121.4205, 122.2285, 123.0292, 123.8227, 124.609,
  35.39103, 36.17737, 36.97087, 37.77157, 38.57954, 39.3948, 40.2174, 
    41.04737, 41.88473, 42.72949, 43.58167, 44.44125, 45.30825, 46.18263, 
    47.06438, 47.95345, 48.84979, 49.75336, 50.66409, 51.5819, 52.5067, 
    53.43839, 54.37686, 55.32199, 56.27364, 57.23167, 58.19592, 59.16621, 
    60.14237, 61.1242, 62.1115, 63.10404, 64.10159, 65.10393, 66.11079, 
    67.12191, 68.13702, 69.15584, 70.17808, 71.20344, 72.23161, 73.26228, 
    74.29513, 75.32983, 76.36606, 77.40348, 78.44174, 79.48052, 80.51948, 
    81.55826, 82.59652, 83.63394, 84.67017, 85.70487, 86.73772, 87.76839, 
    88.79656, 89.82192, 90.84416, 91.86298, 92.87809, 93.88921, 94.89607, 
    95.89841, 96.89597, 97.8885, 98.8758, 99.85763, 100.8338, 101.8041, 
    102.7683, 103.7264, 104.678, 105.6231, 106.5616, 107.4933, 108.4181, 
    109.3359, 110.2466, 111.1502, 112.0466, 112.9356, 113.8174, 114.6917, 
    115.5587, 116.4183, 117.2705, 118.1153, 118.9526, 119.7826, 120.6052, 
    121.4205, 122.2284, 123.0291, 123.8226, 124.609,
  35.39105, 36.17739, 36.97089, 37.7716, 38.57956, 39.39482, 40.21743, 
    41.04739, 41.88475, 42.72952, 43.58169, 44.44128, 45.30827, 46.18266, 
    47.0644, 47.95347, 48.84982, 49.75339, 50.66412, 51.58192, 52.50672, 
    53.43841, 54.37688, 55.32201, 56.27366, 57.23169, 58.19594, 59.16623, 
    60.14239, 61.12422, 62.11152, 63.10405, 64.10161, 65.10394, 66.1108, 
    67.12192, 68.13703, 69.15585, 70.17809, 71.20345, 72.23161, 73.26228, 
    74.29514, 75.32983, 76.36607, 77.40348, 78.44175, 79.48052, 80.51948, 
    81.55825, 82.59652, 83.63393, 84.67017, 85.70486, 86.73772, 87.76839, 
    88.79655, 89.82191, 90.84415, 91.86297, 92.87808, 93.8892, 94.89606, 
    95.89839, 96.89594, 97.88849, 98.87578, 99.8576, 100.8338, 101.8041, 
    102.7683, 103.7263, 104.678, 105.6231, 106.5616, 107.4933, 108.4181, 
    109.3359, 110.2466, 111.1502, 112.0465, 112.9356, 113.8173, 114.6917, 
    115.5587, 116.4183, 117.2705, 118.1152, 118.9526, 119.7826, 120.6052, 
    121.4204, 122.2284, 123.0291, 123.8226, 124.6089,
  35.39108, 36.17741, 36.97091, 37.77162, 38.57958, 39.39485, 40.21745, 
    41.04742, 41.88477, 42.72954, 43.58171, 44.4413, 45.3083, 46.18268, 
    47.06442, 47.95349, 48.84984, 49.75341, 50.66414, 51.58195, 52.50674, 
    53.43843, 54.3769, 55.32203, 56.27369, 57.23171, 58.19596, 59.16625, 
    60.14241, 61.12424, 62.11153, 63.10407, 64.10162, 65.10396, 66.11082, 
    67.12193, 68.13704, 69.15586, 70.1781, 71.20345, 72.23162, 73.26229, 
    74.29514, 75.32984, 76.36607, 77.40348, 78.44175, 79.48052, 80.51948, 
    81.55825, 82.59652, 83.63393, 84.67016, 85.70486, 86.73771, 87.76838, 
    88.79655, 89.8219, 90.84414, 91.86296, 92.87807, 93.88918, 94.89604, 
    95.89838, 96.89593, 97.88847, 98.87576, 99.85759, 100.8337, 101.804, 
    102.7683, 103.7263, 104.678, 105.6231, 106.5616, 107.4933, 108.4181, 
    109.3359, 110.2466, 111.1502, 112.0465, 112.9356, 113.8173, 114.6917, 
    115.5587, 116.4183, 117.2705, 118.1152, 118.9526, 119.7826, 120.6052, 
    121.4204, 122.2284, 123.0291, 123.8226, 124.6089,
  35.39109, 36.17744, 36.97094, 37.77164, 38.57961, 39.39487, 40.21747, 
    41.04744, 41.8848, 42.72956, 43.58174, 44.44133, 45.30832, 46.1827, 
    47.06445, 47.95351, 48.84986, 49.75343, 50.66416, 51.58197, 52.50677, 
    53.43846, 54.37693, 55.32205, 56.2737, 57.23173, 58.19598, 59.16627, 
    60.14243, 61.12426, 62.11155, 63.10409, 64.10165, 65.10397, 66.11083, 
    67.12195, 68.13705, 69.15587, 70.17811, 71.20346, 72.23163, 73.2623, 
    74.29514, 75.32985, 76.36607, 77.40349, 78.44175, 79.48053, 80.51947, 
    81.55825, 82.59651, 83.63393, 84.67015, 85.70486, 86.7377, 87.76837, 
    88.79654, 89.82189, 90.84413, 91.86295, 92.87805, 93.88917, 94.89603, 
    95.89835, 96.89591, 97.88845, 98.87574, 99.85757, 100.8337, 101.804, 
    102.7683, 103.7263, 104.6779, 105.6231, 106.5615, 107.4932, 108.418, 
    109.3358, 110.2466, 111.1501, 112.0465, 112.9356, 113.8173, 114.6917, 
    115.5587, 116.4183, 117.2704, 118.1152, 118.9526, 119.7825, 120.6051, 
    121.4204, 122.2284, 123.0291, 123.8226, 124.6089,
  35.39112, 36.17746, 36.97095, 37.77166, 38.57963, 39.39489, 40.21749, 
    41.04746, 41.88482, 42.72958, 43.58176, 44.44135, 45.30835, 46.18273, 
    47.06447, 47.95354, 48.84988, 49.75346, 50.66418, 51.58199, 52.50679, 
    53.43848, 54.37695, 55.32207, 56.27372, 57.23175, 58.196, 59.16629, 
    60.14245, 61.12428, 62.11156, 63.1041, 64.10166, 65.10399, 66.11084, 
    67.12196, 68.13707, 69.15588, 70.17812, 71.20347, 72.23164, 73.26231, 
    74.29515, 75.32985, 76.36607, 77.40349, 78.44175, 79.48053, 80.51947, 
    81.55825, 82.59651, 83.63393, 84.67015, 85.70485, 86.73769, 87.76836, 
    88.79653, 89.82188, 90.84412, 91.86293, 92.87804, 93.88916, 94.89601, 
    95.89834, 96.8959, 97.88844, 98.87572, 99.85755, 100.8337, 101.804, 
    102.7682, 103.7263, 104.6779, 105.6231, 106.5615, 107.4932, 108.418, 
    109.3358, 110.2465, 111.1501, 112.0465, 112.9355, 113.8173, 114.6917, 
    115.5586, 116.4182, 117.2704, 118.1152, 118.9525, 119.7825, 120.6051, 
    121.4204, 122.2283, 123.029, 123.8225, 124.6089,
  35.39114, 36.17748, 36.97098, 37.77168, 38.57965, 39.39491, 40.21751, 
    41.04749, 41.88484, 42.72961, 43.58178, 44.44137, 45.30836, 46.18275, 
    47.06449, 47.95356, 48.84991, 49.75348, 50.6642, 51.58201, 52.50681, 
    53.4385, 54.37697, 55.32209, 56.27374, 57.23177, 58.19601, 59.16631, 
    60.14246, 61.12429, 62.11158, 63.10412, 64.10167, 65.104, 66.11086, 
    67.12197, 68.13708, 69.15589, 70.17813, 71.20348, 72.23165, 73.26231, 
    74.29516, 75.32986, 76.36608, 77.40349, 78.44175, 79.48053, 80.51947, 
    81.55825, 82.59651, 83.63392, 84.67014, 85.70484, 86.73769, 87.76835, 
    88.79652, 89.82187, 90.84411, 91.86292, 92.87803, 93.88914, 94.896, 
    95.89833, 96.89588, 97.88842, 98.87571, 99.85754, 100.8337, 101.804, 
    102.7682, 103.7263, 104.6779, 105.623, 106.5615, 107.4932, 108.418, 
    109.3358, 110.2465, 111.1501, 112.0464, 112.9355, 113.8173, 114.6916, 
    115.5586, 116.4182, 117.2704, 118.1152, 118.9525, 119.7825, 120.6051, 
    121.4203, 122.2283, 123.029, 123.8225, 124.6089,
  35.39116, 36.1775, 36.971, 37.77171, 38.57967, 39.39494, 40.21754, 41.0475, 
    41.88486, 42.72963, 43.5818, 44.44139, 45.30839, 46.18277, 47.06451, 
    47.95358, 48.84993, 49.7535, 50.66423, 51.58203, 52.50683, 53.43852, 
    54.37699, 55.32211, 56.27377, 57.23179, 58.19603, 59.16632, 60.14248, 
    61.12431, 62.1116, 63.10413, 64.10168, 65.10402, 66.11087, 67.12199, 
    68.13709, 69.15591, 70.17814, 71.20349, 72.23166, 73.26232, 74.29517, 
    75.32986, 76.36608, 77.4035, 78.44176, 79.48053, 80.51947, 81.55824, 
    82.5965, 83.63392, 84.67014, 85.70483, 86.73768, 87.76834, 88.79651, 
    89.82186, 90.84409, 91.86291, 92.87801, 93.88913, 94.89598, 95.89832, 
    96.89587, 97.8884, 98.87569, 99.85752, 100.8337, 101.804, 102.7682, 
    103.7262, 104.6779, 105.623, 106.5615, 107.4932, 108.418, 109.3358, 
    110.2465, 111.1501, 112.0464, 112.9355, 113.8172, 114.6916, 115.5586, 
    116.4182, 117.2704, 118.1151, 118.9525, 119.7825, 120.6051, 121.4203, 
    122.2283, 123.029, 123.8225, 124.6088,
  35.39117, 36.17752, 36.97102, 37.77172, 38.57969, 39.39495, 40.21756, 
    41.04753, 41.88488, 42.72965, 43.58183, 44.44141, 45.30841, 46.18279, 
    47.06453, 47.9536, 48.84995, 49.75352, 50.66425, 51.58205, 52.50685, 
    53.43854, 54.37701, 55.32213, 56.27378, 57.23181, 58.19605, 59.16634, 
    60.1425, 61.12432, 62.11161, 63.10415, 64.1017, 65.10403, 66.11088, 
    67.12199, 68.1371, 69.15591, 70.17815, 71.2035, 72.23167, 73.26233, 
    74.29517, 75.32986, 76.36609, 77.4035, 78.44176, 79.48053, 80.51947, 
    81.55824, 82.5965, 83.63391, 84.67014, 85.70483, 86.73767, 87.76833, 
    88.7965, 89.82185, 90.84409, 91.8629, 92.87801, 93.88912, 94.89597, 
    95.8983, 96.89585, 97.88838, 98.87568, 99.8575, 100.8337, 101.8039, 
    102.7682, 103.7262, 104.6779, 105.623, 106.5615, 107.4931, 108.4179, 
    109.3358, 110.2465, 111.15, 112.0464, 112.9355, 113.8172, 114.6916, 
    115.5586, 116.4182, 117.2704, 118.1151, 118.9525, 119.7824, 120.605, 
    121.4203, 122.2283, 123.029, 123.8225, 124.6088,
  35.39119, 36.17754, 36.97104, 37.77174, 38.57971, 39.39497, 40.21758, 
    41.04755, 41.8849, 42.72967, 43.58184, 44.44143, 45.30843, 46.18281, 
    47.06456, 47.95362, 48.84997, 49.75354, 50.66426, 51.58207, 52.50687, 
    53.43856, 54.37703, 55.32215, 56.2738, 57.23183, 58.19607, 59.16636, 
    60.14251, 61.12434, 62.11163, 63.10416, 64.10172, 65.10404, 66.11089, 
    67.12201, 68.13711, 69.15592, 70.17815, 71.20351, 72.23167, 73.26234, 
    74.29517, 75.32987, 76.36609, 77.4035, 78.44176, 79.48053, 80.51947, 
    81.55824, 82.5965, 83.63391, 84.67013, 85.70483, 86.73766, 87.76833, 
    88.79649, 89.82185, 90.84408, 91.86289, 92.87799, 93.88911, 94.89596, 
    95.89828, 96.89584, 97.88837, 98.87566, 99.85748, 100.8336, 101.8039, 
    102.7682, 103.7262, 104.6778, 105.623, 106.5614, 107.4931, 108.4179, 
    109.3357, 110.2465, 111.15, 112.0464, 112.9354, 113.8172, 114.6916, 
    115.5586, 116.4182, 117.2703, 118.1151, 118.9525, 119.7824, 120.605, 
    121.4203, 122.2283, 123.029, 123.8225, 124.6088,
  35.39121, 36.17756, 36.97105, 37.77176, 38.57973, 39.39499, 40.21759, 
    41.04757, 41.88492, 42.72969, 43.58186, 44.44145, 45.30845, 46.18283, 
    47.06458, 47.95364, 48.84999, 49.75356, 50.66428, 51.58209, 52.50689, 
    53.43858, 54.37704, 55.32217, 56.27382, 57.23184, 58.19609, 59.16637, 
    60.14253, 61.12436, 62.11164, 63.10418, 64.10173, 65.10406, 66.11091, 
    67.12202, 68.13712, 69.15594, 70.17816, 71.20351, 72.23167, 73.26234, 
    74.29518, 75.32987, 76.3661, 77.4035, 78.44176, 79.48053, 80.51947, 
    81.55824, 82.5965, 83.6339, 84.67013, 85.70482, 86.73766, 87.76833, 
    88.79649, 89.82184, 90.84406, 91.86288, 92.87798, 93.88909, 94.89594, 
    95.89827, 96.89582, 97.88836, 98.87564, 99.85747, 100.8336, 101.8039, 
    102.7682, 103.7262, 104.6778, 105.623, 106.5614, 107.4931, 108.4179, 
    109.3357, 110.2464, 111.15, 112.0464, 112.9354, 113.8172, 114.6916, 
    115.5585, 116.4181, 117.2703, 118.1151, 118.9524, 119.7824, 120.605, 
    121.4203, 122.2282, 123.0289, 123.8224, 124.6088,
  35.39123, 36.17757, 36.97107, 37.77178, 38.57975, 39.39501, 40.21761, 
    41.04758, 41.88494, 42.72971, 43.58188, 44.44147, 45.30847, 46.18285, 
    47.06459, 47.95366, 48.85001, 49.75358, 50.6643, 51.58211, 52.5069, 
    53.43859, 54.37706, 55.32219, 56.27383, 57.23186, 58.1961, 59.16639, 
    60.14255, 61.12437, 62.11166, 63.10419, 64.10175, 65.10406, 66.11092, 
    67.12203, 68.13713, 69.15594, 70.17818, 71.20352, 72.23168, 73.26234, 
    74.29519, 75.32988, 76.3661, 77.4035, 78.44176, 79.48053, 80.51947, 
    81.55824, 82.5965, 83.6339, 84.67012, 85.70481, 86.73766, 87.76832, 
    88.79648, 89.82182, 90.84406, 91.86287, 92.87797, 93.88908, 94.89594, 
    95.89825, 96.89581, 97.88834, 98.87563, 99.85745, 100.8336, 101.8039, 
    102.7681, 103.7262, 104.6778, 105.6229, 106.5614, 107.4931, 108.4179, 
    109.3357, 110.2464, 111.15, 112.0463, 112.9354, 113.8172, 114.6915, 
    115.5585, 116.4181, 117.2703, 118.1151, 118.9524, 119.7824, 120.605, 
    121.4203, 122.2282, 123.0289, 123.8224, 124.6088,
  35.39124, 36.17759, 36.97109, 37.7718, 38.57976, 39.39503, 40.21763, 
    41.0476, 41.88496, 42.72972, 43.5819, 44.44149, 45.30849, 46.18287, 
    47.06461, 47.95368, 48.85003, 49.75359, 50.66432, 51.58213, 52.50692, 
    53.43861, 54.37708, 55.3222, 56.27385, 57.23188, 58.19612, 59.16641, 
    60.14256, 61.12439, 62.11167, 63.10421, 64.10175, 65.10408, 66.11093, 
    67.12204, 68.13714, 69.15595, 70.17818, 71.20353, 72.23169, 73.26235, 
    74.29519, 75.32989, 76.3661, 77.4035, 78.44176, 79.48053, 80.51947, 
    81.55824, 82.5965, 83.6339, 84.67011, 85.70481, 86.73765, 87.76831, 
    88.79647, 89.82182, 90.84405, 91.86286, 92.87796, 93.88907, 94.89592, 
    95.89825, 96.8958, 97.88833, 98.87562, 99.85744, 100.8336, 101.8039, 
    102.7681, 103.7262, 104.6778, 105.6229, 106.5614, 107.4931, 108.4179, 
    109.3357, 110.2464, 111.15, 112.0463, 112.9354, 113.8171, 114.6915, 
    115.5585, 116.4181, 117.2703, 118.115, 118.9524, 119.7824, 120.605, 
    121.4202, 122.2282, 123.0289, 123.8224, 124.6088,
  35.39126, 36.1776, 36.9711, 37.77181, 38.57978, 39.39504, 40.21765, 
    41.04762, 41.88498, 42.72974, 43.58192, 44.44151, 45.3085, 46.18288, 
    47.06463, 47.95369, 48.85004, 49.75361, 50.66434, 51.58214, 52.50694, 
    53.43863, 54.37709, 55.32222, 56.27387, 57.23189, 58.19613, 59.16642, 
    60.14257, 61.1244, 62.11169, 63.10422, 64.10177, 65.10409, 66.11094, 
    67.12205, 68.13715, 69.15596, 70.17819, 71.20354, 72.2317, 73.26236, 
    74.2952, 75.32989, 76.3661, 77.40351, 78.44176, 79.48053, 80.51947, 
    81.55824, 82.59649, 83.6339, 84.67011, 85.7048, 86.73764, 87.7683, 
    88.79646, 89.82181, 90.84404, 91.86285, 92.87795, 93.88906, 94.89591, 
    95.89823, 96.89578, 97.88831, 98.8756, 99.85742, 100.8336, 101.8039, 
    102.7681, 103.7261, 104.6778, 105.6229, 106.5614, 107.4931, 108.4179, 
    109.3357, 110.2464, 111.15, 112.0463, 112.9354, 113.8171, 114.6915, 
    115.5585, 116.4181, 117.2703, 118.115, 118.9524, 119.7824, 120.605, 
    121.4202, 122.2282, 123.0289, 123.8224, 124.6087,
  35.39127, 36.17762, 36.97112, 37.77183, 38.57979, 39.39506, 40.21766, 
    41.04763, 41.88499, 42.72976, 43.58193, 44.44152, 45.30852, 46.1829, 
    47.06464, 47.95371, 48.85006, 49.75363, 50.66435, 51.58216, 52.50695, 
    53.43864, 54.37711, 55.32224, 56.27388, 57.23191, 58.19615, 59.16644, 
    60.14259, 61.12441, 62.1117, 63.10423, 64.10178, 65.1041, 66.11095, 
    67.12206, 68.13716, 69.15597, 70.1782, 71.20354, 72.2317, 73.26236, 
    74.2952, 75.3299, 76.3661, 77.40351, 78.44176, 79.48053, 80.51947, 
    81.55824, 82.59649, 83.6339, 84.6701, 85.7048, 86.73764, 87.7683, 
    88.79646, 89.8218, 90.84403, 91.86284, 92.87794, 93.88905, 94.8959, 
    95.89822, 96.89577, 97.88831, 98.87559, 99.85741, 100.8336, 101.8039, 
    102.7681, 103.7261, 104.6778, 105.6229, 106.5614, 107.493, 108.4178, 
    109.3356, 110.2464, 111.1499, 112.0463, 112.9354, 113.8171, 114.6915, 
    115.5585, 116.4181, 117.2702, 118.115, 118.9524, 119.7823, 120.6049, 
    121.4202, 122.2282, 123.0289, 123.8224, 124.6087,
  35.39129, 36.17763, 36.97113, 37.77184, 38.57981, 39.39507, 40.21768, 
    41.04765, 41.88501, 42.72977, 43.58195, 44.44154, 45.30853, 46.18291, 
    47.06466, 47.95373, 48.85007, 49.75364, 50.66437, 51.58217, 52.50697, 
    53.43866, 54.37712, 55.32225, 56.2739, 57.23192, 58.19616, 59.16645, 
    60.1426, 61.12442, 62.11171, 63.10424, 64.10179, 65.10411, 66.11096, 
    67.12207, 68.13717, 69.15598, 70.17821, 71.20355, 72.23171, 73.26237, 
    74.2952, 75.3299, 76.36611, 77.40351, 78.44176, 79.48053, 80.51947, 
    81.55824, 82.59649, 83.63389, 84.6701, 85.7048, 86.73763, 87.76829, 
    88.79645, 89.82179, 90.84402, 91.86283, 92.87793, 93.88904, 94.89589, 
    95.89821, 96.89576, 97.88829, 98.87558, 99.8574, 100.8335, 101.8038, 
    102.7681, 103.7261, 104.6777, 105.6229, 106.5613, 107.493, 108.4178, 
    109.3356, 110.2464, 111.1499, 112.0463, 112.9353, 113.8171, 114.6915, 
    115.5585, 116.4181, 117.2702, 118.115, 118.9524, 119.7823, 120.6049, 
    121.4202, 122.2282, 123.0289, 123.8224, 124.6087,
  35.3913, 36.17765, 36.97115, 37.77185, 38.57982, 39.39509, 40.21769, 
    41.04766, 41.88502, 42.72979, 43.58196, 44.44155, 45.30855, 46.18293, 
    47.06467, 47.95374, 48.85009, 49.75366, 50.66438, 51.58219, 52.50698, 
    53.43867, 54.37714, 55.32226, 56.27391, 57.23193, 58.19617, 59.16646, 
    60.14261, 61.12444, 62.11172, 63.10425, 64.1018, 65.10413, 66.11097, 
    67.12208, 68.13718, 69.15598, 70.17822, 71.20356, 72.23171, 73.26237, 
    74.29521, 75.3299, 76.36611, 77.40351, 78.44176, 79.48053, 80.51947, 
    81.55824, 82.59649, 83.63389, 84.6701, 85.70479, 86.73763, 87.76829, 
    88.79644, 89.82178, 90.84402, 91.86282, 92.87792, 93.88903, 94.89587, 
    95.8982, 96.89574, 97.88828, 98.87556, 99.85738, 100.8335, 101.8038, 
    102.7681, 103.7261, 104.6777, 105.6229, 106.5613, 107.493, 108.4178, 
    109.3356, 110.2463, 111.1499, 112.0463, 112.9353, 113.8171, 114.6915, 
    115.5584, 116.418, 117.2702, 118.115, 118.9523, 119.7823, 120.6049, 
    121.4202, 122.2281, 123.0289, 123.8224, 124.6087,
  35.39131, 36.17766, 36.97116, 37.77187, 38.57983, 39.3951, 40.2177, 
    41.04767, 41.88503, 42.7298, 43.58197, 44.44157, 45.30856, 46.18295, 
    47.06469, 47.95375, 48.8501, 49.75367, 50.6644, 51.5822, 52.507, 
    53.43868, 54.37715, 55.32228, 56.27392, 57.23195, 58.19619, 59.16647, 
    60.14262, 61.12445, 62.11173, 63.10426, 64.10181, 65.10413, 66.11098, 
    67.12209, 68.13718, 69.15599, 70.17822, 71.20356, 72.23172, 73.26237, 
    74.29521, 75.3299, 76.36611, 77.40352, 78.44176, 79.48053, 80.51947, 
    81.55824, 82.59648, 83.63389, 84.6701, 85.70479, 86.73763, 87.76828, 
    88.79644, 89.82178, 90.84401, 91.86282, 92.87791, 93.88902, 94.89587, 
    95.89819, 96.89574, 97.88827, 98.87556, 99.85738, 100.8335, 101.8038, 
    102.7681, 103.7261, 104.6777, 105.6228, 106.5613, 107.493, 108.4178, 
    109.3356, 110.2463, 111.1499, 112.0462, 112.9353, 113.8171, 114.6914, 
    115.5584, 116.418, 117.2702, 118.115, 118.9523, 119.7823, 120.6049, 
    121.4202, 122.2281, 123.0288, 123.8223, 124.6087,
  35.39132, 36.17767, 36.97117, 37.77188, 38.57985, 39.39511, 40.21772, 
    41.04769, 41.88504, 42.72981, 43.58199, 44.44158, 45.30857, 46.18296, 
    47.0647, 47.95377, 48.85011, 49.75368, 50.66441, 51.58221, 52.50701, 
    53.4387, 54.37716, 55.32229, 56.27393, 57.23196, 58.1962, 59.16648, 
    60.14264, 61.12446, 62.11174, 63.10427, 64.10182, 65.10414, 66.11098, 
    67.12209, 68.13719, 69.156, 70.17822, 71.20357, 72.23173, 73.26238, 
    74.29522, 75.3299, 76.36612, 77.40352, 78.44177, 79.48053, 80.51947, 
    81.55823, 82.59648, 83.63388, 84.6701, 85.70478, 86.73762, 87.76827, 
    88.79643, 89.82178, 90.844, 91.86281, 92.87791, 93.88902, 94.89586, 
    95.89818, 96.89573, 97.88826, 98.87554, 99.85736, 100.8335, 101.8038, 
    102.768, 103.7261, 104.6777, 105.6228, 106.5613, 107.493, 108.4178, 
    109.3356, 110.2463, 111.1499, 112.0462, 112.9353, 113.817, 114.6914, 
    115.5584, 116.418, 117.2702, 118.115, 118.9523, 119.7823, 120.6049, 
    121.4202, 122.2281, 123.0288, 123.8223, 124.6087,
  35.39133, 36.17768, 36.97118, 37.77189, 38.57986, 39.39512, 40.21773, 
    41.0477, 41.88506, 42.72982, 43.582, 44.44159, 45.30859, 46.18297, 
    47.06471, 47.95378, 48.85013, 49.7537, 50.66442, 51.58223, 52.50702, 
    53.43871, 54.37717, 55.3223, 56.27394, 57.23197, 58.19621, 59.16649, 
    60.14265, 61.12447, 62.11175, 63.10428, 64.10183, 65.10415, 66.11099, 
    67.1221, 68.1372, 69.15601, 70.17823, 71.20358, 72.23173, 73.26238, 
    74.29522, 75.32991, 76.36612, 77.40352, 78.44177, 79.48053, 80.51947, 
    81.55823, 82.59648, 83.63388, 84.67009, 85.70478, 86.73762, 87.76827, 
    88.79642, 89.82177, 90.84399, 91.8628, 92.8779, 93.88901, 94.89585, 
    95.89817, 96.89572, 97.88825, 98.87553, 99.85735, 100.8335, 101.8038, 
    102.768, 103.7261, 104.6777, 105.6228, 106.5613, 107.493, 108.4178, 
    109.3356, 110.2463, 111.1499, 112.0462, 112.9353, 113.817, 114.6914, 
    115.5584, 116.418, 117.2702, 118.1149, 118.9523, 119.7823, 120.6049, 
    121.4201, 122.2281, 123.0288, 123.8223, 124.6087,
  35.39134, 36.17769, 36.97119, 37.7719, 38.57987, 39.39513, 40.21774, 
    41.04771, 41.88507, 42.72983, 43.58201, 44.4416, 45.3086, 46.18298, 
    47.06472, 47.95379, 48.85014, 49.75371, 50.66443, 51.58224, 52.50703, 
    53.43872, 54.37719, 55.32231, 56.27396, 57.23198, 58.19622, 59.1665, 
    60.14265, 61.12447, 62.11176, 63.10429, 64.10184, 65.10416, 66.111, 
    67.12211, 68.13721, 69.15601, 70.17824, 71.20358, 72.23174, 73.26239, 
    74.29522, 75.32991, 76.36612, 77.40352, 78.44177, 79.48053, 80.51947, 
    81.55823, 82.59648, 83.63388, 84.67009, 85.70478, 86.73761, 87.76826, 
    88.79642, 89.82176, 90.84399, 91.86279, 92.87789, 93.889, 94.89584, 
    95.89816, 96.89571, 97.88824, 98.87553, 99.85735, 100.8335, 101.8038, 
    102.768, 103.726, 104.6777, 105.6228, 106.5613, 107.493, 108.4178, 
    109.3356, 110.2463, 111.1499, 112.0462, 112.9353, 113.817, 114.6914, 
    115.5584, 116.418, 117.2702, 118.1149, 118.9523, 119.7823, 120.6049, 
    121.4201, 122.2281, 123.0288, 123.8223, 124.6087,
  35.39135, 36.1777, 36.9712, 37.77191, 38.57988, 39.39514, 40.21775, 
    41.04772, 41.88508, 42.72984, 43.58202, 44.44161, 45.30861, 46.18299, 
    47.06473, 47.9538, 48.85015, 49.75372, 50.66444, 51.58225, 52.50704, 
    53.43873, 54.37719, 55.32232, 56.27396, 57.23199, 58.19622, 59.16651, 
    60.14266, 61.12449, 62.11177, 63.1043, 64.10184, 65.10416, 66.11101, 
    67.12212, 68.13721, 69.15601, 70.17824, 71.20358, 72.23174, 73.26239, 
    74.29523, 75.32991, 76.36612, 77.40352, 78.44177, 79.48054, 80.51946, 
    81.55823, 82.59648, 83.63388, 84.67009, 85.70477, 86.73761, 87.76826, 
    88.79642, 89.82176, 90.84399, 91.86279, 92.87788, 93.88899, 94.89584, 
    95.89816, 96.89571, 97.88823, 98.87552, 99.85734, 100.8335, 101.8038, 
    102.768, 103.726, 104.6777, 105.6228, 106.5613, 107.493, 108.4178, 
    109.3356, 110.2463, 111.1498, 112.0462, 112.9353, 113.817, 114.6914, 
    115.5584, 116.418, 117.2702, 118.1149, 118.9523, 119.7822, 120.6049, 
    121.4201, 122.2281, 123.0288, 123.8223, 124.6087,
  35.39136, 36.17771, 36.97121, 37.77192, 38.57988, 39.39515, 40.21775, 
    41.04773, 41.88509, 42.72985, 43.58203, 44.44162, 45.30862, 46.183, 
    47.06474, 47.95381, 48.85015, 49.75373, 50.66445, 51.58226, 52.50705, 
    53.43874, 54.3772, 55.32233, 56.27397, 57.23199, 58.19624, 59.16652, 
    60.14267, 61.12449, 62.11177, 63.10431, 64.10185, 65.10417, 66.11102, 
    67.12212, 68.13721, 69.15602, 70.17825, 71.20358, 72.23174, 73.2624, 
    74.29523, 75.32992, 76.36613, 77.40353, 78.44177, 79.48054, 80.51946, 
    81.55823, 82.59647, 83.63387, 84.67008, 85.70477, 86.7376, 87.76826, 
    88.79642, 89.82175, 90.84398, 91.86279, 92.87788, 93.88898, 94.89583, 
    95.89815, 96.8957, 97.88822, 98.87551, 99.85733, 100.8335, 101.8038, 
    102.768, 103.726, 104.6777, 105.6228, 106.5613, 107.493, 108.4177, 
    109.3355, 110.2463, 111.1498, 112.0462, 112.9353, 113.817, 114.6914, 
    115.5584, 116.418, 117.2701, 118.1149, 118.9523, 119.7822, 120.6049, 
    121.4201, 122.2281, 123.0288, 123.8223, 124.6086,
  35.39137, 36.17771, 36.97121, 37.77192, 38.57989, 39.39516, 40.21776, 
    41.04773, 41.88509, 42.72986, 43.58204, 44.44163, 45.30862, 46.18301, 
    47.06475, 47.95382, 48.85017, 49.75373, 50.66446, 51.58226, 52.50706, 
    53.43874, 54.37721, 55.32233, 56.27398, 57.232, 58.19624, 59.16653, 
    60.14268, 61.1245, 62.11178, 63.10431, 64.10185, 65.10417, 66.11102, 
    67.12212, 68.13722, 69.15603, 70.17825, 71.20359, 72.23174, 73.2624, 
    74.29523, 75.32992, 76.36613, 77.40353, 78.44177, 79.48054, 80.51946, 
    81.55823, 82.59647, 83.63387, 84.67008, 85.70477, 86.7376, 87.76826, 
    88.79641, 89.82175, 90.84397, 91.86278, 92.87788, 93.88898, 94.89583, 
    95.89815, 96.89569, 97.88822, 98.8755, 99.85732, 100.8335, 101.8038, 
    102.768, 103.726, 104.6777, 105.6228, 106.5613, 107.4929, 108.4177, 
    109.3355, 110.2463, 111.1498, 112.0462, 112.9352, 113.817, 114.6914, 
    115.5584, 116.418, 117.2701, 118.1149, 118.9523, 119.7822, 120.6048, 
    121.4201, 122.2281, 123.0288, 123.8223, 124.6086,
  35.39137, 36.17772, 36.97122, 37.77193, 38.5799, 39.39516, 40.21777, 
    41.04774, 41.8851, 42.72987, 43.58204, 44.44164, 45.30863, 46.18301, 
    47.06476, 47.95383, 48.85017, 49.75374, 50.66447, 51.58227, 52.50706, 
    53.43875, 54.37722, 55.32234, 56.27399, 57.23201, 58.19625, 59.16653, 
    60.14268, 61.1245, 62.11179, 63.10432, 64.10186, 65.10418, 66.11102, 
    67.12213, 68.13722, 69.15603, 70.17825, 71.20359, 72.23175, 73.2624, 
    74.29523, 75.32992, 76.36613, 77.40353, 78.44177, 79.48054, 80.51946, 
    81.55823, 82.59647, 83.63387, 84.67008, 85.70477, 86.7376, 87.76825, 
    88.79641, 89.82175, 90.84397, 91.86278, 92.87787, 93.88898, 94.89582, 
    95.89814, 96.89568, 97.88821, 98.8755, 99.85732, 100.8335, 101.8037, 
    102.768, 103.726, 104.6777, 105.6228, 106.5612, 107.4929, 108.4177, 
    109.3355, 110.2463, 111.1498, 112.0462, 112.9352, 113.817, 114.6914, 
    115.5584, 116.418, 117.2701, 118.1149, 118.9523, 119.7822, 120.6048, 
    121.4201, 122.2281, 123.0288, 123.8223, 124.6086,
  35.39138, 36.17772, 36.97123, 37.77193, 38.5799, 39.39517, 40.21778, 
    41.04775, 41.88511, 42.72987, 43.58205, 44.44164, 45.30864, 46.18302, 
    47.06476, 47.95383, 48.85018, 49.75375, 50.66447, 51.58228, 52.50707, 
    53.43876, 54.37722, 55.32235, 56.27399, 57.23201, 58.19625, 59.16654, 
    60.14269, 61.12451, 62.11179, 63.10432, 64.10187, 65.10419, 66.11103, 
    67.12213, 68.13723, 69.15603, 70.17825, 71.2036, 72.23175, 73.26241, 
    74.29523, 75.32992, 76.36613, 77.40353, 78.44177, 79.48054, 80.51946, 
    81.55823, 82.59647, 83.63387, 84.67008, 85.70477, 86.73759, 87.76825, 
    88.7964, 89.82175, 90.84397, 91.86277, 92.87787, 93.88897, 94.89581, 
    95.89813, 96.89568, 97.88821, 98.87549, 99.85731, 100.8335, 101.8037, 
    102.768, 103.726, 104.6777, 105.6228, 106.5612, 107.4929, 108.4177, 
    109.3355, 110.2463, 111.1498, 112.0462, 112.9352, 113.817, 114.6914, 
    115.5584, 116.4179, 117.2701, 118.1149, 118.9523, 119.7822, 120.6048, 
    121.4201, 122.2281, 123.0288, 123.8223, 124.6086,
  35.39138, 36.17773, 36.97123, 37.77194, 38.57991, 39.39518, 40.21778, 
    41.04775, 41.88511, 42.72988, 43.58205, 44.44165, 45.30864, 46.18303, 
    47.06477, 47.95383, 48.85018, 49.75375, 50.66448, 51.58228, 52.50708, 
    53.43876, 54.37723, 55.32235, 56.274, 57.23202, 58.19626, 59.16654, 
    60.14269, 61.12451, 62.1118, 63.10432, 64.10187, 65.10419, 66.11103, 
    67.12214, 68.13723, 69.15604, 70.17826, 71.2036, 72.23175, 73.26241, 
    74.29523, 75.32992, 76.36613, 77.40353, 78.44177, 79.48054, 80.51946, 
    81.55823, 82.59647, 83.63387, 84.67008, 85.70477, 86.73759, 87.76825, 
    88.7964, 89.82174, 90.84396, 91.86277, 92.87786, 93.88897, 94.89581, 
    95.89813, 96.89568, 97.88821, 98.87549, 99.85731, 100.8335, 101.8037, 
    102.768, 103.726, 104.6777, 105.6228, 106.5612, 107.4929, 108.4177, 
    109.3355, 110.2462, 111.1498, 112.0462, 112.9352, 113.817, 114.6914, 
    115.5583, 116.4179, 117.2701, 118.1149, 118.9522, 119.7822, 120.6048, 
    121.4201, 122.2281, 123.0288, 123.8223, 124.6086,
  35.39139, 36.17773, 36.97123, 37.77195, 38.57991, 39.39518, 40.21778, 
    41.04776, 41.88512, 42.72988, 43.58206, 44.44165, 45.30865, 46.18303, 
    47.06477, 47.95384, 48.85019, 49.75376, 50.66448, 51.58229, 52.50708, 
    53.43877, 54.37723, 55.32236, 56.274, 57.23202, 58.19626, 59.16655, 
    60.1427, 61.12452, 62.1118, 63.10433, 64.10187, 65.10419, 66.11103, 
    67.12214, 68.13724, 69.15604, 70.17826, 71.2036, 72.23175, 73.26241, 
    74.29523, 75.32993, 76.36613, 77.40353, 78.44177, 79.48054, 80.51946, 
    81.55823, 82.59647, 83.63387, 84.67007, 85.70477, 86.73759, 87.76825, 
    88.7964, 89.82174, 90.84396, 91.86276, 92.87786, 93.88897, 94.89581, 
    95.89813, 96.89568, 97.8882, 98.87548, 99.8573, 100.8335, 101.8037, 
    102.768, 103.726, 104.6776, 105.6228, 106.5612, 107.4929, 108.4177, 
    109.3355, 110.2462, 111.1498, 112.0462, 112.9352, 113.817, 114.6914, 
    115.5583, 116.4179, 117.2701, 118.1149, 118.9522, 119.7822, 120.6048, 
    121.4201, 122.2281, 123.0288, 123.8223, 124.6086,
  35.39139, 36.17773, 36.97124, 37.77195, 38.57991, 39.39518, 40.21779, 
    41.04776, 41.88512, 42.72989, 43.58206, 44.44165, 45.30865, 46.18303, 
    47.06478, 47.95384, 48.85019, 49.75376, 50.66449, 51.58229, 52.50708, 
    53.43877, 54.37724, 55.32236, 56.27401, 57.23203, 58.19626, 59.16655, 
    60.1427, 61.12452, 62.1118, 63.10433, 64.10188, 65.10419, 66.11104, 
    67.12214, 68.13724, 69.15604, 70.17826, 71.2036, 72.23176, 73.26241, 
    74.29523, 75.32993, 76.36613, 77.40353, 78.44177, 79.48054, 80.51946, 
    81.55823, 82.59647, 83.63387, 84.67007, 85.70477, 86.73759, 87.76824, 
    88.7964, 89.82174, 90.84396, 91.86276, 92.87786, 93.88896, 94.89581, 
    95.89812, 96.89567, 97.8882, 98.87548, 99.8573, 100.8335, 101.8037, 
    102.768, 103.726, 104.6776, 105.6228, 106.5612, 107.4929, 108.4177, 
    109.3355, 110.2462, 111.1498, 112.0462, 112.9352, 113.817, 114.6914, 
    115.5583, 116.4179, 117.2701, 118.1149, 118.9522, 119.7822, 120.6048, 
    121.4201, 122.2281, 123.0288, 123.8223, 124.6086,
  35.39139, 36.17774, 36.97124, 37.77195, 38.57992, 39.39518, 40.21779, 
    41.04776, 41.88512, 42.72989, 43.58207, 44.44165, 45.30865, 46.18303, 
    47.06478, 47.95385, 48.85019, 49.75376, 50.66449, 51.58229, 52.50709, 
    53.43877, 54.37724, 55.32236, 56.27401, 57.23203, 58.19627, 59.16655, 
    60.1427, 61.12452, 62.1118, 63.10433, 64.10188, 65.10419, 66.11104, 
    67.12214, 68.13724, 69.15604, 70.17826, 71.20361, 72.23176, 73.26241, 
    74.29524, 75.32993, 76.36613, 77.40353, 78.44177, 79.48054, 80.51946, 
    81.55823, 82.59647, 83.63387, 84.67007, 85.70476, 86.73759, 87.76824, 
    88.79639, 89.82174, 90.84396, 91.86276, 92.87786, 93.88896, 94.89581, 
    95.89812, 96.89567, 97.8882, 98.87548, 99.8573, 100.8335, 101.8037, 
    102.768, 103.726, 104.6776, 105.6228, 106.5612, 107.4929, 108.4177, 
    109.3355, 110.2462, 111.1498, 112.0462, 112.9352, 113.817, 114.6913, 
    115.5583, 116.4179, 117.2701, 118.1149, 118.9522, 119.7822, 120.6048, 
    121.4201, 122.2281, 123.0288, 123.8223, 124.6086,
  35.39139, 36.17774, 36.97124, 37.77195, 38.57992, 39.39519, 40.21779, 
    41.04776, 41.88512, 42.72989, 43.58207, 44.44166, 45.30865, 46.18304, 
    47.06478, 47.95385, 48.85019, 49.75376, 50.66449, 51.58229, 52.50709, 
    53.43877, 54.37724, 55.32236, 56.27401, 57.23203, 58.19627, 59.16655, 
    60.1427, 61.12452, 62.1118, 63.10433, 64.10188, 65.10419, 66.11104, 
    67.12214, 68.13724, 69.15604, 70.17826, 71.20361, 72.23176, 73.26241, 
    74.29524, 75.32993, 76.36613, 77.40353, 78.44177, 79.48054, 80.51946, 
    81.55823, 82.59647, 83.63387, 84.67007, 85.70476, 86.73759, 87.76824, 
    88.79639, 89.82174, 90.84396, 91.86276, 92.87786, 93.88896, 94.89581, 
    95.89812, 96.89567, 97.8882, 98.87548, 99.8573, 100.8335, 101.8037, 
    102.768, 103.726, 104.6776, 105.6228, 106.5612, 107.4929, 108.4177, 
    109.3355, 110.2462, 111.1498, 112.0462, 112.9352, 113.817, 114.6913, 
    115.5583, 116.4179, 117.2701, 118.1149, 118.9522, 119.7822, 120.6048, 
    121.4201, 122.2281, 123.0288, 123.8223, 124.6086,
  35.39139, 36.17774, 36.97124, 37.77195, 38.57992, 39.39519, 40.21779, 
    41.04776, 41.88512, 42.72989, 43.58207, 44.44166, 45.30865, 46.18304, 
    47.06478, 47.95385, 48.85019, 49.75376, 50.66449, 51.58229, 52.50709, 
    53.43877, 54.37724, 55.32236, 56.27401, 57.23203, 58.19627, 59.16655, 
    60.1427, 61.12452, 62.1118, 63.10433, 64.10188, 65.10419, 66.11104, 
    67.12214, 68.13724, 69.15604, 70.17826, 71.20361, 72.23176, 73.26241, 
    74.29524, 75.32993, 76.36613, 77.40353, 78.44177, 79.48054, 80.51946, 
    81.55823, 82.59647, 83.63387, 84.67007, 85.70476, 86.73759, 87.76824, 
    88.79639, 89.82174, 90.84396, 91.86276, 92.87786, 93.88896, 94.89581, 
    95.89812, 96.89567, 97.8882, 98.87548, 99.8573, 100.8335, 101.8037, 
    102.768, 103.726, 104.6776, 105.6228, 106.5612, 107.4929, 108.4177, 
    109.3355, 110.2462, 111.1498, 112.0462, 112.9352, 113.817, 114.6913, 
    115.5583, 116.4179, 117.2701, 118.1149, 118.9522, 119.7822, 120.6048, 
    121.4201, 122.2281, 123.0288, 123.8223, 124.6086,
  35.39139, 36.17774, 36.97124, 37.77195, 38.57992, 39.39518, 40.21779, 
    41.04776, 41.88512, 42.72989, 43.58207, 44.44165, 45.30865, 46.18303, 
    47.06478, 47.95385, 48.85019, 49.75376, 50.66449, 51.58229, 52.50709, 
    53.43877, 54.37724, 55.32236, 56.27401, 57.23203, 58.19627, 59.16655, 
    60.1427, 61.12452, 62.1118, 63.10433, 64.10188, 65.10419, 66.11104, 
    67.12214, 68.13724, 69.15604, 70.17826, 71.20361, 72.23176, 73.26241, 
    74.29524, 75.32993, 76.36613, 77.40353, 78.44177, 79.48054, 80.51946, 
    81.55823, 82.59647, 83.63387, 84.67007, 85.70476, 86.73759, 87.76824, 
    88.79639, 89.82174, 90.84396, 91.86276, 92.87786, 93.88896, 94.89581, 
    95.89812, 96.89567, 97.8882, 98.87548, 99.8573, 100.8335, 101.8037, 
    102.768, 103.726, 104.6776, 105.6228, 106.5612, 107.4929, 108.4177, 
    109.3355, 110.2462, 111.1498, 112.0462, 112.9352, 113.817, 114.6913, 
    115.5583, 116.4179, 117.2701, 118.1149, 118.9522, 119.7822, 120.6048, 
    121.4201, 122.2281, 123.0288, 123.8223, 124.6086,
  35.39139, 36.17773, 36.97124, 37.77195, 38.57991, 39.39518, 40.21779, 
    41.04776, 41.88512, 42.72989, 43.58206, 44.44165, 45.30865, 46.18303, 
    47.06478, 47.95384, 48.85019, 49.75376, 50.66449, 51.58229, 52.50708, 
    53.43877, 54.37724, 55.32236, 56.27401, 57.23203, 58.19626, 59.16655, 
    60.1427, 61.12452, 62.1118, 63.10433, 64.10188, 65.10419, 66.11104, 
    67.12214, 68.13724, 69.15604, 70.17826, 71.2036, 72.23176, 73.26241, 
    74.29523, 75.32993, 76.36613, 77.40353, 78.44177, 79.48054, 80.51946, 
    81.55823, 82.59647, 83.63387, 84.67007, 85.70477, 86.73759, 87.76824, 
    88.7964, 89.82174, 90.84396, 91.86276, 92.87786, 93.88896, 94.89581, 
    95.89812, 96.89567, 97.8882, 98.87548, 99.8573, 100.8335, 101.8037, 
    102.768, 103.726, 104.6776, 105.6228, 106.5612, 107.4929, 108.4177, 
    109.3355, 110.2462, 111.1498, 112.0462, 112.9352, 113.817, 114.6914, 
    115.5583, 116.4179, 117.2701, 118.1149, 118.9522, 119.7822, 120.6048, 
    121.4201, 122.2281, 123.0288, 123.8223, 124.6086,
  35.39139, 36.17773, 36.97123, 37.77195, 38.57991, 39.39518, 40.21778, 
    41.04776, 41.88512, 42.72988, 43.58206, 44.44165, 45.30865, 46.18303, 
    47.06477, 47.95384, 48.85019, 49.75376, 50.66448, 51.58229, 52.50708, 
    53.43877, 54.37723, 55.32236, 56.274, 57.23202, 58.19626, 59.16655, 
    60.1427, 61.12452, 62.1118, 63.10433, 64.10187, 65.10419, 66.11103, 
    67.12214, 68.13724, 69.15604, 70.17826, 71.2036, 72.23175, 73.26241, 
    74.29523, 75.32993, 76.36613, 77.40353, 78.44177, 79.48054, 80.51946, 
    81.55823, 82.59647, 83.63387, 84.67007, 85.70477, 86.73759, 87.76825, 
    88.7964, 89.82174, 90.84396, 91.86276, 92.87786, 93.88897, 94.89581, 
    95.89813, 96.89568, 97.8882, 98.87548, 99.8573, 100.8335, 101.8037, 
    102.768, 103.726, 104.6776, 105.6228, 106.5612, 107.4929, 108.4177, 
    109.3355, 110.2462, 111.1498, 112.0462, 112.9352, 113.817, 114.6914, 
    115.5583, 116.4179, 117.2701, 118.1149, 118.9522, 119.7822, 120.6048, 
    121.4201, 122.2281, 123.0288, 123.8223, 124.6086,
  35.39138, 36.17773, 36.97123, 37.77194, 38.57991, 39.39518, 40.21778, 
    41.04775, 41.88511, 42.72988, 43.58205, 44.44165, 45.30864, 46.18303, 
    47.06477, 47.95383, 48.85018, 49.75375, 50.66448, 51.58228, 52.50708, 
    53.43876, 54.37723, 55.32235, 56.274, 57.23202, 58.19626, 59.16654, 
    60.14269, 61.12451, 62.1118, 63.10432, 64.10187, 65.10419, 66.11103, 
    67.12214, 68.13723, 69.15604, 70.17826, 71.2036, 72.23175, 73.26241, 
    74.29523, 75.32992, 76.36613, 77.40353, 78.44177, 79.48054, 80.51946, 
    81.55823, 82.59647, 83.63387, 84.67008, 85.70477, 86.73759, 87.76825, 
    88.7964, 89.82174, 90.84396, 91.86277, 92.87786, 93.88897, 94.89581, 
    95.89813, 96.89568, 97.88821, 98.87549, 99.85731, 100.8335, 101.8037, 
    102.768, 103.726, 104.6777, 105.6228, 106.5612, 107.4929, 108.4177, 
    109.3355, 110.2462, 111.1498, 112.0462, 112.9352, 113.817, 114.6914, 
    115.5583, 116.4179, 117.2701, 118.1149, 118.9522, 119.7822, 120.6048, 
    121.4201, 122.2281, 123.0288, 123.8223, 124.6086,
  35.39138, 36.17772, 36.97123, 37.77193, 38.5799, 39.39517, 40.21778, 
    41.04775, 41.88511, 42.72987, 43.58205, 44.44164, 45.30864, 46.18302, 
    47.06476, 47.95383, 48.85018, 49.75375, 50.66447, 51.58228, 52.50707, 
    53.43876, 54.37722, 55.32235, 56.27399, 57.23201, 58.19625, 59.16654, 
    60.14269, 61.12451, 62.11179, 63.10432, 64.10187, 65.10419, 66.11103, 
    67.12213, 68.13723, 69.15603, 70.17825, 71.2036, 72.23175, 73.26241, 
    74.29523, 75.32992, 76.36613, 77.40353, 78.44177, 79.48054, 80.51946, 
    81.55823, 82.59647, 83.63387, 84.67008, 85.70477, 86.73759, 87.76825, 
    88.7964, 89.82175, 90.84397, 91.86277, 92.87787, 93.88897, 94.89581, 
    95.89813, 96.89568, 97.88821, 98.87549, 99.85731, 100.8335, 101.8037, 
    102.768, 103.726, 104.6777, 105.6228, 106.5612, 107.4929, 108.4177, 
    109.3355, 110.2463, 111.1498, 112.0462, 112.9352, 113.817, 114.6914, 
    115.5584, 116.4179, 117.2701, 118.1149, 118.9523, 119.7822, 120.6048, 
    121.4201, 122.2281, 123.0288, 123.8223, 124.6086,
  35.39137, 36.17772, 36.97122, 37.77193, 38.5799, 39.39516, 40.21777, 
    41.04774, 41.8851, 42.72987, 43.58204, 44.44164, 45.30863, 46.18301, 
    47.06476, 47.95383, 48.85017, 49.75374, 50.66447, 51.58227, 52.50706, 
    53.43875, 54.37722, 55.32234, 56.27399, 57.23201, 58.19625, 59.16653, 
    60.14268, 61.1245, 62.11179, 63.10432, 64.10186, 65.10418, 66.11102, 
    67.12213, 68.13722, 69.15603, 70.17825, 71.20359, 72.23175, 73.2624, 
    74.29523, 75.32992, 76.36613, 77.40353, 78.44177, 79.48054, 80.51946, 
    81.55823, 82.59647, 83.63387, 84.67008, 85.70477, 86.7376, 87.76825, 
    88.79641, 89.82175, 90.84397, 91.86278, 92.87787, 93.88898, 94.89582, 
    95.89814, 96.89568, 97.88821, 98.8755, 99.85732, 100.8335, 101.8037, 
    102.768, 103.726, 104.6777, 105.6228, 106.5612, 107.4929, 108.4177, 
    109.3355, 110.2463, 111.1498, 112.0462, 112.9352, 113.817, 114.6914, 
    115.5584, 116.418, 117.2701, 118.1149, 118.9523, 119.7822, 120.6048, 
    121.4201, 122.2281, 123.0288, 123.8223, 124.6086,
  35.39137, 36.17771, 36.97121, 37.77192, 38.57989, 39.39516, 40.21776, 
    41.04773, 41.88509, 42.72986, 43.58204, 44.44163, 45.30862, 46.18301, 
    47.06475, 47.95382, 48.85017, 49.75373, 50.66446, 51.58226, 52.50706, 
    53.43874, 54.37721, 55.32233, 56.27398, 57.232, 58.19624, 59.16653, 
    60.14268, 61.1245, 62.11178, 63.10431, 64.10185, 65.10417, 66.11102, 
    67.12212, 68.13722, 69.15603, 70.17825, 71.20359, 72.23174, 73.2624, 
    74.29523, 75.32992, 76.36613, 77.40353, 78.44177, 79.48054, 80.51946, 
    81.55823, 82.59647, 83.63387, 84.67008, 85.70477, 86.7376, 87.76826, 
    88.79641, 89.82175, 90.84397, 91.86278, 92.87788, 93.88898, 94.89583, 
    95.89815, 96.89569, 97.88822, 98.8755, 99.85732, 100.8335, 101.8038, 
    102.768, 103.726, 104.6777, 105.6228, 106.5613, 107.4929, 108.4177, 
    109.3355, 110.2463, 111.1498, 112.0462, 112.9352, 113.817, 114.6914, 
    115.5584, 116.418, 117.2701, 118.1149, 118.9523, 119.7822, 120.6048, 
    121.4201, 122.2281, 123.0288, 123.8223, 124.6086,
  35.39136, 36.17771, 36.97121, 37.77192, 38.57988, 39.39515, 40.21775, 
    41.04773, 41.88509, 42.72985, 43.58203, 44.44162, 45.30862, 46.183, 
    47.06474, 47.95381, 48.85015, 49.75373, 50.66445, 51.58226, 52.50705, 
    53.43874, 54.3772, 55.32233, 56.27397, 57.23199, 58.19624, 59.16652, 
    60.14267, 61.12449, 62.11177, 63.10431, 64.10185, 65.10417, 66.11102, 
    67.12212, 68.13721, 69.15602, 70.17825, 71.20358, 72.23174, 73.2624, 
    74.29523, 75.32992, 76.36613, 77.40353, 78.44177, 79.48054, 80.51946, 
    81.55823, 82.59647, 83.63387, 84.67008, 85.70477, 86.7376, 87.76826, 
    88.79642, 89.82175, 90.84398, 91.86279, 92.87788, 93.88898, 94.89583, 
    95.89815, 96.8957, 97.88822, 98.87551, 99.85733, 100.8335, 101.8038, 
    102.768, 103.726, 104.6777, 105.6228, 106.5613, 107.493, 108.4177, 
    109.3355, 110.2463, 111.1498, 112.0462, 112.9353, 113.817, 114.6914, 
    115.5584, 116.418, 117.2701, 118.1149, 118.9523, 119.7822, 120.6049, 
    121.4201, 122.2281, 123.0288, 123.8223, 124.6086,
  35.39135, 36.1777, 36.9712, 37.77191, 38.57988, 39.39514, 40.21775, 
    41.04772, 41.88508, 42.72984, 43.58202, 44.44161, 45.30861, 46.18299, 
    47.06473, 47.9538, 48.85015, 49.75372, 50.66444, 51.58225, 52.50704, 
    53.43873, 54.37719, 55.32232, 56.27396, 57.23199, 58.19622, 59.16651, 
    60.14266, 61.12449, 62.11177, 63.1043, 64.10184, 65.10416, 66.11101, 
    67.12212, 68.13721, 69.15601, 70.17824, 71.20358, 72.23174, 73.26239, 
    74.29523, 75.32991, 76.36612, 77.40352, 78.44177, 79.48054, 80.51946, 
    81.55823, 82.59648, 83.63388, 84.67009, 85.70477, 86.73761, 87.76826, 
    88.79642, 89.82176, 90.84399, 91.86279, 92.87788, 93.88899, 94.89584, 
    95.89816, 96.89571, 97.88823, 98.87552, 99.85734, 100.8335, 101.8038, 
    102.768, 103.726, 104.6777, 105.6228, 106.5613, 107.493, 108.4178, 
    109.3356, 110.2463, 111.1498, 112.0462, 112.9353, 113.817, 114.6914, 
    115.5584, 116.418, 117.2702, 118.1149, 118.9523, 119.7822, 120.6049, 
    121.4201, 122.2281, 123.0288, 123.8223, 124.6087,
  35.39134, 36.17769, 36.97119, 37.7719, 38.57987, 39.39513, 40.21774, 
    41.04771, 41.88507, 42.72983, 43.58201, 44.4416, 45.3086, 46.18298, 
    47.06472, 47.95379, 48.85014, 49.75371, 50.66443, 51.58224, 52.50703, 
    53.43872, 54.37719, 55.32231, 56.27396, 57.23198, 58.19622, 59.1665, 
    60.14265, 61.12447, 62.11176, 63.10429, 64.10184, 65.10416, 66.111, 
    67.12211, 68.13721, 69.15601, 70.17824, 71.20358, 72.23174, 73.26239, 
    74.29522, 75.32991, 76.36612, 77.40352, 78.44177, 79.48053, 80.51947, 
    81.55823, 82.59648, 83.63388, 84.67009, 85.70478, 86.73761, 87.76826, 
    88.79642, 89.82176, 90.84399, 91.86279, 92.87789, 93.889, 94.89584, 
    95.89816, 96.89571, 97.88824, 98.87553, 99.85735, 100.8335, 101.8038, 
    102.768, 103.726, 104.6777, 105.6228, 106.5613, 107.493, 108.4178, 
    109.3356, 110.2463, 111.1499, 112.0462, 112.9353, 113.817, 114.6914, 
    115.5584, 116.418, 117.2702, 118.1149, 118.9523, 119.7823, 120.6049, 
    121.4201, 122.2281, 123.0288, 123.8223, 124.6087,
  35.39133, 36.17768, 36.97118, 37.77189, 38.57986, 39.39512, 40.21773, 
    41.0477, 41.88506, 42.72982, 43.582, 44.44159, 45.30859, 46.18297, 
    47.06471, 47.95378, 48.85013, 49.7537, 50.66442, 51.58223, 52.50702, 
    53.43871, 54.37717, 55.3223, 56.27394, 57.23197, 58.19621, 59.16649, 
    60.14265, 61.12447, 62.11175, 63.10428, 64.10183, 65.10415, 66.11099, 
    67.1221, 68.1372, 69.15601, 70.17823, 71.20358, 72.23173, 73.26238, 
    74.29522, 75.32991, 76.36612, 77.40352, 78.44177, 79.48053, 80.51947, 
    81.55823, 82.59648, 83.63388, 84.67009, 85.70478, 86.73762, 87.76827, 
    88.79642, 89.82177, 90.84399, 91.8628, 92.8779, 93.88901, 94.89585, 
    95.89817, 96.89572, 97.88825, 98.87553, 99.85735, 100.8335, 101.8038, 
    102.768, 103.7261, 104.6777, 105.6228, 106.5613, 107.493, 108.4178, 
    109.3356, 110.2463, 111.1499, 112.0462, 112.9353, 113.817, 114.6914, 
    115.5584, 116.418, 117.2702, 118.1149, 118.9523, 119.7823, 120.6049, 
    121.4201, 122.2281, 123.0288, 123.8223, 124.6087,
  35.39132, 36.17767, 36.97117, 37.77188, 38.57985, 39.39511, 40.21772, 
    41.04769, 41.88504, 42.72981, 43.58199, 44.44158, 45.30857, 46.18296, 
    47.0647, 47.95377, 48.85011, 49.75368, 50.66441, 51.58221, 52.50701, 
    53.4387, 54.37716, 55.32229, 56.27393, 57.23196, 58.1962, 59.16648, 
    60.14264, 61.12446, 62.11174, 63.10427, 64.10182, 65.10414, 66.11098, 
    67.12209, 68.13719, 69.156, 70.17822, 71.20357, 72.23173, 73.26238, 
    74.29522, 75.3299, 76.36612, 77.40352, 78.44177, 79.48053, 80.51947, 
    81.55823, 82.59648, 83.63388, 84.6701, 85.70478, 86.73762, 87.76827, 
    88.79643, 89.82178, 90.844, 91.86281, 92.87791, 93.88902, 94.89586, 
    95.89818, 96.89573, 97.88826, 98.87554, 99.85736, 100.8335, 101.8038, 
    102.768, 103.7261, 104.6777, 105.6228, 106.5613, 107.493, 108.4178, 
    109.3356, 110.2463, 111.1499, 112.0462, 112.9353, 113.817, 114.6914, 
    115.5584, 116.418, 117.2702, 118.115, 118.9523, 119.7823, 120.6049, 
    121.4202, 122.2281, 123.0288, 123.8223, 124.6087,
  35.39131, 36.17766, 36.97116, 37.77187, 38.57983, 39.3951, 40.2177, 
    41.04767, 41.88503, 42.7298, 43.58197, 44.44157, 45.30856, 46.18295, 
    47.06469, 47.95375, 48.8501, 49.75367, 50.6644, 51.5822, 52.507, 
    53.43868, 54.37715, 55.32228, 56.27392, 57.23195, 58.19619, 59.16647, 
    60.14262, 61.12445, 62.11173, 63.10426, 64.10181, 65.10413, 66.11098, 
    67.12209, 68.13718, 69.15599, 70.17822, 71.20356, 72.23172, 73.26237, 
    74.29521, 75.3299, 76.36611, 77.40352, 78.44176, 79.48053, 80.51947, 
    81.55824, 82.59648, 83.63389, 84.6701, 85.70479, 86.73763, 87.76828, 
    88.79644, 89.82178, 90.84401, 91.86282, 92.87791, 93.88902, 94.89587, 
    95.89819, 96.89574, 97.88827, 98.87556, 99.85738, 100.8335, 101.8038, 
    102.7681, 103.7261, 104.6777, 105.6228, 106.5613, 107.493, 108.4178, 
    109.3356, 110.2463, 111.1499, 112.0462, 112.9353, 113.8171, 114.6914, 
    115.5584, 116.418, 117.2702, 118.115, 118.9523, 119.7823, 120.6049, 
    121.4202, 122.2281, 123.0288, 123.8223, 124.6087,
  35.3913, 36.17765, 36.97115, 37.77185, 38.57982, 39.39509, 40.21769, 
    41.04766, 41.88502, 42.72979, 43.58196, 44.44155, 45.30855, 46.18293, 
    47.06467, 47.95374, 48.85009, 49.75366, 50.66438, 51.58219, 52.50698, 
    53.43867, 54.37714, 55.32226, 56.27391, 57.23193, 58.19617, 59.16646, 
    60.14261, 61.12444, 62.11172, 63.10425, 64.1018, 65.10413, 66.11097, 
    67.12208, 68.13718, 69.15598, 70.17822, 71.20356, 72.23171, 73.26237, 
    74.29521, 75.3299, 76.36611, 77.40351, 78.44176, 79.48053, 80.51947, 
    81.55824, 82.59649, 83.63389, 84.6701, 85.70479, 86.73763, 87.76829, 
    88.79644, 89.82178, 90.84402, 91.86282, 92.87792, 93.88903, 94.89587, 
    95.8982, 96.89574, 97.88828, 98.87556, 99.85738, 100.8335, 101.8038, 
    102.7681, 103.7261, 104.6777, 105.6229, 106.5613, 107.493, 108.4178, 
    109.3356, 110.2463, 111.1499, 112.0463, 112.9353, 113.8171, 114.6915, 
    115.5584, 116.418, 117.2702, 118.115, 118.9523, 119.7823, 120.6049, 
    121.4202, 122.2281, 123.0289, 123.8224, 124.6087,
  35.39129, 36.17763, 36.97113, 37.77184, 38.57981, 39.39507, 40.21768, 
    41.04765, 41.88501, 42.72977, 43.58195, 44.44154, 45.30853, 46.18291, 
    47.06466, 47.95373, 48.85007, 49.75364, 50.66437, 51.58217, 52.50697, 
    53.43866, 54.37712, 55.32225, 56.2739, 57.23192, 58.19616, 59.16645, 
    60.1426, 61.12442, 62.11171, 63.10424, 64.10179, 65.10411, 66.11096, 
    67.12207, 68.13717, 69.15598, 70.17821, 71.20355, 72.23171, 73.26237, 
    74.2952, 75.3299, 76.36611, 77.40351, 78.44176, 79.48053, 80.51947, 
    81.55824, 82.59649, 83.63389, 84.6701, 85.7048, 86.73763, 87.76829, 
    88.79645, 89.82179, 90.84402, 91.86283, 92.87793, 93.88904, 94.89589, 
    95.89821, 96.89576, 97.88829, 98.87558, 99.8574, 100.8335, 101.8038, 
    102.7681, 103.7261, 104.6777, 105.6229, 106.5613, 107.493, 108.4178, 
    109.3356, 110.2464, 111.1499, 112.0463, 112.9353, 113.8171, 114.6915, 
    115.5585, 116.4181, 117.2702, 118.115, 118.9524, 119.7823, 120.6049, 
    121.4202, 122.2282, 123.0289, 123.8224, 124.6087,
  35.39127, 36.17762, 36.97112, 37.77183, 38.57979, 39.39506, 40.21766, 
    41.04763, 41.88499, 42.72976, 43.58193, 44.44152, 45.30852, 46.1829, 
    47.06464, 47.95371, 48.85006, 49.75363, 50.66435, 51.58216, 52.50695, 
    53.43864, 54.37711, 55.32224, 56.27388, 57.23191, 58.19615, 59.16644, 
    60.14259, 61.12441, 62.1117, 63.10423, 64.10178, 65.1041, 66.11095, 
    67.12206, 68.13716, 69.15597, 70.1782, 71.20354, 72.2317, 73.26236, 
    74.2952, 75.3299, 76.3661, 77.40351, 78.44176, 79.48053, 80.51947, 
    81.55824, 82.59649, 83.6339, 84.6701, 85.7048, 86.73764, 87.7683, 
    88.79646, 89.8218, 90.84403, 91.86284, 92.87794, 93.88905, 94.8959, 
    95.89822, 96.89577, 97.88831, 98.87559, 99.85741, 100.8336, 101.8039, 
    102.7681, 103.7261, 104.6778, 105.6229, 106.5614, 107.493, 108.4178, 
    109.3356, 110.2464, 111.1499, 112.0463, 112.9354, 113.8171, 114.6915, 
    115.5585, 116.4181, 117.2702, 118.115, 118.9524, 119.7823, 120.6049, 
    121.4202, 122.2282, 123.0289, 123.8224, 124.6087,
  35.39126, 36.1776, 36.9711, 37.77181, 38.57978, 39.39504, 40.21765, 
    41.04762, 41.88498, 42.72974, 43.58192, 44.44151, 45.3085, 46.18288, 
    47.06463, 47.95369, 48.85004, 49.75361, 50.66434, 51.58214, 52.50694, 
    53.43863, 54.37709, 55.32222, 56.27387, 57.23189, 58.19613, 59.16642, 
    60.14257, 61.1244, 62.11169, 63.10422, 64.10177, 65.10409, 66.11094, 
    67.12205, 68.13715, 69.15596, 70.17819, 71.20354, 72.2317, 73.26236, 
    74.2952, 75.32989, 76.3661, 77.40351, 78.44176, 79.48053, 80.51947, 
    81.55824, 82.59649, 83.6339, 84.67011, 85.7048, 86.73764, 87.7683, 
    88.79646, 89.82181, 90.84404, 91.86285, 92.87795, 93.88906, 94.89591, 
    95.89823, 96.89578, 97.88831, 98.8756, 99.85742, 100.8336, 101.8039, 
    102.7681, 103.7261, 104.6778, 105.6229, 106.5614, 107.4931, 108.4179, 
    109.3357, 110.2464, 111.15, 112.0463, 112.9354, 113.8171, 114.6915, 
    115.5585, 116.4181, 117.2703, 118.115, 118.9524, 119.7824, 120.605, 
    121.4202, 122.2282, 123.0289, 123.8224, 124.6087,
  35.39124, 36.17759, 36.97109, 37.7718, 38.57976, 39.39503, 40.21763, 
    41.0476, 41.88496, 42.72972, 43.5819, 44.44149, 45.30849, 46.18287, 
    47.06461, 47.95368, 48.85003, 49.75359, 50.66432, 51.58213, 52.50692, 
    53.43861, 54.37708, 55.3222, 56.27385, 57.23188, 58.19612, 59.16641, 
    60.14256, 61.12439, 62.11167, 63.10421, 64.10175, 65.10408, 66.11093, 
    67.12204, 68.13714, 69.15595, 70.17818, 71.20353, 72.23169, 73.26235, 
    74.29519, 75.32989, 76.3661, 77.4035, 78.44176, 79.48053, 80.51947, 
    81.55824, 82.5965, 83.6339, 84.67011, 85.70481, 86.73765, 87.76831, 
    88.79647, 89.82182, 90.84405, 91.86286, 92.87796, 93.88907, 94.89592, 
    95.89825, 96.8958, 97.88833, 98.87562, 99.85744, 100.8336, 101.8039, 
    102.7681, 103.7262, 104.6778, 105.6229, 106.5614, 107.4931, 108.4179, 
    109.3357, 110.2464, 111.15, 112.0463, 112.9354, 113.8171, 114.6915, 
    115.5585, 116.4181, 117.2703, 118.115, 118.9524, 119.7824, 120.605, 
    121.4202, 122.2282, 123.0289, 123.8224, 124.6088,
  35.39123, 36.17757, 36.97107, 37.77178, 38.57975, 39.39501, 40.21761, 
    41.04758, 41.88494, 42.72971, 43.58188, 44.44147, 45.30847, 46.18285, 
    47.06459, 47.95366, 48.85001, 49.75358, 50.6643, 51.58211, 52.5069, 
    53.43859, 54.37706, 55.32219, 56.27383, 57.23186, 58.1961, 59.16639, 
    60.14255, 61.12437, 62.11166, 63.10419, 64.10175, 65.10406, 66.11092, 
    67.12203, 68.13713, 69.15594, 70.17818, 71.20352, 72.23168, 73.26234, 
    74.29519, 75.32988, 76.3661, 77.4035, 78.44176, 79.48053, 80.51947, 
    81.55824, 82.5965, 83.6339, 84.67012, 85.70481, 86.73766, 87.76832, 
    88.79648, 89.82182, 90.84406, 91.86287, 92.87797, 93.88908, 94.89594, 
    95.89825, 96.89581, 97.88834, 98.87563, 99.85745, 100.8336, 101.8039, 
    102.7681, 103.7262, 104.6778, 105.6229, 106.5614, 107.4931, 108.4179, 
    109.3357, 110.2464, 111.15, 112.0463, 112.9354, 113.8172, 114.6915, 
    115.5585, 116.4181, 117.2703, 118.1151, 118.9524, 119.7824, 120.605, 
    121.4203, 122.2282, 123.0289, 123.8224, 124.6088,
  35.39121, 36.17756, 36.97105, 37.77176, 38.57973, 39.39499, 40.21759, 
    41.04757, 41.88492, 42.72969, 43.58186, 44.44145, 45.30845, 46.18283, 
    47.06458, 47.95364, 48.84999, 49.75356, 50.66428, 51.58209, 52.50689, 
    53.43858, 54.37704, 55.32217, 56.27382, 57.23184, 58.19609, 59.16637, 
    60.14253, 61.12436, 62.11164, 63.10418, 64.10173, 65.10406, 66.11091, 
    67.12202, 68.13712, 69.15594, 70.17816, 71.20351, 72.23167, 73.26234, 
    74.29518, 75.32987, 76.3661, 77.4035, 78.44176, 79.48053, 80.51947, 
    81.55824, 82.5965, 83.6339, 84.67013, 85.70482, 86.73766, 87.76833, 
    88.79649, 89.82184, 90.84406, 91.86288, 92.87798, 93.88909, 94.89594, 
    95.89827, 96.89582, 97.88836, 98.87564, 99.85747, 100.8336, 101.8039, 
    102.7682, 103.7262, 104.6778, 105.623, 106.5614, 107.4931, 108.4179, 
    109.3357, 110.2464, 111.15, 112.0464, 112.9354, 113.8172, 114.6916, 
    115.5585, 116.4181, 117.2703, 118.1151, 118.9524, 119.7824, 120.605, 
    121.4203, 122.2282, 123.0289, 123.8224, 124.6088,
  35.39119, 36.17754, 36.97104, 37.77174, 38.57971, 39.39497, 40.21758, 
    41.04755, 41.8849, 42.72967, 43.58184, 44.44143, 45.30843, 46.18281, 
    47.06456, 47.95362, 48.84997, 49.75354, 50.66426, 51.58207, 52.50687, 
    53.43856, 54.37703, 55.32215, 56.2738, 57.23183, 58.19607, 59.16636, 
    60.14251, 61.12434, 62.11163, 63.10416, 64.10172, 65.10404, 66.11089, 
    67.12201, 68.13711, 69.15592, 70.17815, 71.20351, 72.23167, 73.26234, 
    74.29517, 75.32987, 76.36609, 77.4035, 78.44176, 79.48053, 80.51947, 
    81.55824, 82.5965, 83.63391, 84.67013, 85.70483, 86.73766, 87.76833, 
    88.79649, 89.82185, 90.84408, 91.86289, 92.87799, 93.88911, 94.89596, 
    95.89828, 96.89584, 97.88837, 98.87566, 99.85748, 100.8336, 101.8039, 
    102.7682, 103.7262, 104.6778, 105.623, 106.5614, 107.4931, 108.4179, 
    109.3357, 110.2465, 111.15, 112.0464, 112.9354, 113.8172, 114.6916, 
    115.5586, 116.4182, 117.2703, 118.1151, 118.9525, 119.7824, 120.605, 
    121.4203, 122.2283, 123.029, 123.8225, 124.6088,
  35.39117, 36.17752, 36.97102, 37.77172, 38.57969, 39.39495, 40.21756, 
    41.04753, 41.88488, 42.72965, 43.58183, 44.44141, 45.30841, 46.18279, 
    47.06453, 47.9536, 48.84995, 49.75352, 50.66425, 51.58205, 52.50685, 
    53.43854, 54.37701, 55.32213, 56.27378, 57.23181, 58.19605, 59.16634, 
    60.1425, 61.12432, 62.11161, 63.10415, 64.1017, 65.10403, 66.11088, 
    67.12199, 68.1371, 69.15591, 70.17815, 71.2035, 72.23167, 73.26233, 
    74.29517, 75.32986, 76.36609, 77.4035, 78.44176, 79.48053, 80.51947, 
    81.55824, 82.5965, 83.63391, 84.67014, 85.70483, 86.73767, 87.76833, 
    88.7965, 89.82185, 90.84409, 91.8629, 92.87801, 93.88912, 94.89597, 
    95.8983, 96.89585, 97.88838, 98.87568, 99.8575, 100.8337, 101.8039, 
    102.7682, 103.7262, 104.6779, 105.623, 106.5615, 107.4931, 108.4179, 
    109.3358, 110.2465, 111.15, 112.0464, 112.9355, 113.8172, 114.6916, 
    115.5586, 116.4182, 117.2704, 118.1151, 118.9525, 119.7824, 120.605, 
    121.4203, 122.2283, 123.029, 123.8225, 124.6088,
  35.39116, 36.1775, 36.971, 37.77171, 38.57967, 39.39494, 40.21754, 41.0475, 
    41.88486, 42.72963, 43.5818, 44.44139, 45.30839, 46.18277, 47.06451, 
    47.95358, 48.84993, 49.7535, 50.66423, 51.58203, 52.50683, 53.43852, 
    54.37699, 55.32211, 56.27377, 57.23179, 58.19603, 59.16632, 60.14248, 
    61.12431, 62.1116, 63.10413, 64.10168, 65.10402, 66.11087, 67.12199, 
    68.13709, 69.15591, 70.17814, 71.20349, 72.23166, 73.26232, 74.29517, 
    75.32986, 76.36608, 77.4035, 78.44176, 79.48053, 80.51947, 81.55824, 
    82.5965, 83.63392, 84.67014, 85.70483, 86.73768, 87.76834, 88.79651, 
    89.82186, 90.84409, 91.86291, 92.87801, 93.88913, 94.89598, 95.89832, 
    96.89587, 97.8884, 98.87569, 99.85752, 100.8337, 101.804, 102.7682, 
    103.7262, 104.6779, 105.623, 106.5615, 107.4932, 108.418, 109.3358, 
    110.2465, 111.1501, 112.0464, 112.9355, 113.8172, 114.6916, 115.5586, 
    116.4182, 117.2704, 118.1151, 118.9525, 119.7825, 120.6051, 121.4203, 
    122.2283, 123.029, 123.8225, 124.6088,
  35.39114, 36.17748, 36.97098, 37.77168, 38.57965, 39.39491, 40.21751, 
    41.04749, 41.88484, 42.72961, 43.58178, 44.44137, 45.30836, 46.18275, 
    47.06449, 47.95356, 48.84991, 49.75348, 50.6642, 51.58201, 52.50681, 
    53.4385, 54.37697, 55.32209, 56.27374, 57.23177, 58.19601, 59.16631, 
    60.14246, 61.12429, 62.11158, 63.10412, 64.10167, 65.104, 66.11086, 
    67.12197, 68.13708, 69.15589, 70.17813, 71.20348, 72.23165, 73.26231, 
    74.29516, 75.32986, 76.36608, 77.40349, 78.44175, 79.48053, 80.51947, 
    81.55825, 82.59651, 83.63392, 84.67014, 85.70484, 86.73769, 87.76835, 
    88.79652, 89.82187, 90.84411, 91.86292, 92.87803, 93.88914, 94.896, 
    95.89833, 96.89588, 97.88842, 98.87571, 99.85754, 100.8337, 101.804, 
    102.7682, 103.7263, 104.6779, 105.623, 106.5615, 107.4932, 108.418, 
    109.3358, 110.2465, 111.1501, 112.0464, 112.9355, 113.8173, 114.6916, 
    115.5586, 116.4182, 117.2704, 118.1152, 118.9525, 119.7825, 120.6051, 
    121.4203, 122.2283, 123.029, 123.8225, 124.6089,
  35.39112, 36.17746, 36.97095, 37.77166, 38.57963, 39.39489, 40.21749, 
    41.04746, 41.88482, 42.72958, 43.58176, 44.44135, 45.30835, 46.18273, 
    47.06447, 47.95354, 48.84988, 49.75346, 50.66418, 51.58199, 52.50679, 
    53.43848, 54.37695, 55.32207, 56.27372, 57.23175, 58.196, 59.16629, 
    60.14245, 61.12428, 62.11156, 63.1041, 64.10166, 65.10399, 66.11084, 
    67.12196, 68.13707, 69.15588, 70.17812, 71.20347, 72.23164, 73.26231, 
    74.29515, 75.32985, 76.36607, 77.40349, 78.44175, 79.48053, 80.51947, 
    81.55825, 82.59651, 83.63393, 84.67015, 85.70485, 86.73769, 87.76836, 
    88.79653, 89.82188, 90.84412, 91.86293, 92.87804, 93.88916, 94.89601, 
    95.89834, 96.8959, 97.88844, 98.87572, 99.85755, 100.8337, 101.804, 
    102.7682, 103.7263, 104.6779, 105.6231, 106.5615, 107.4932, 108.418, 
    109.3358, 110.2465, 111.1501, 112.0465, 112.9355, 113.8173, 114.6917, 
    115.5586, 116.4182, 117.2704, 118.1152, 118.9525, 119.7825, 120.6051, 
    121.4204, 122.2283, 123.029, 123.8225, 124.6089,
  35.39109, 36.17744, 36.97094, 37.77164, 38.57961, 39.39487, 40.21747, 
    41.04744, 41.8848, 42.72956, 43.58174, 44.44133, 45.30832, 46.1827, 
    47.06445, 47.95351, 48.84986, 49.75343, 50.66416, 51.58197, 52.50677, 
    53.43846, 54.37693, 55.32205, 56.2737, 57.23173, 58.19598, 59.16627, 
    60.14243, 61.12426, 62.11155, 63.10409, 64.10165, 65.10397, 66.11083, 
    67.12195, 68.13705, 69.15587, 70.17811, 71.20346, 72.23163, 73.2623, 
    74.29514, 75.32985, 76.36607, 77.40349, 78.44175, 79.48053, 80.51947, 
    81.55825, 82.59651, 83.63393, 84.67015, 85.70486, 86.7377, 87.76837, 
    88.79654, 89.82189, 90.84413, 91.86295, 92.87805, 93.88917, 94.89603, 
    95.89835, 96.89591, 97.88845, 98.87574, 99.85757, 100.8337, 101.804, 
    102.7683, 103.7263, 104.6779, 105.6231, 106.5615, 107.4932, 108.418, 
    109.3358, 110.2466, 111.1501, 112.0465, 112.9356, 113.8173, 114.6917, 
    115.5587, 116.4183, 117.2704, 118.1152, 118.9526, 119.7825, 120.6051, 
    121.4204, 122.2284, 123.0291, 123.8226, 124.6089,
  35.39108, 36.17741, 36.97091, 37.77162, 38.57958, 39.39485, 40.21745, 
    41.04742, 41.88477, 42.72954, 43.58171, 44.4413, 45.3083, 46.18268, 
    47.06442, 47.95349, 48.84984, 49.75341, 50.66414, 51.58195, 52.50674, 
    53.43843, 54.3769, 55.32203, 56.27369, 57.23171, 58.19596, 59.16625, 
    60.14241, 61.12424, 62.11153, 63.10407, 64.10162, 65.10396, 66.11082, 
    67.12193, 68.13704, 69.15586, 70.1781, 71.20345, 72.23162, 73.26229, 
    74.29514, 75.32984, 76.36607, 77.40348, 78.44175, 79.48052, 80.51948, 
    81.55825, 82.59652, 83.63393, 84.67016, 85.70486, 86.73771, 87.76838, 
    88.79655, 89.8219, 90.84414, 91.86296, 92.87807, 93.88918, 94.89604, 
    95.89838, 96.89593, 97.88847, 98.87576, 99.85759, 100.8337, 101.804, 
    102.7683, 103.7263, 104.678, 105.6231, 106.5616, 107.4933, 108.4181, 
    109.3359, 110.2466, 111.1502, 112.0465, 112.9356, 113.8173, 114.6917, 
    115.5587, 116.4183, 117.2705, 118.1152, 118.9526, 119.7826, 120.6052, 
    121.4204, 122.2284, 123.0291, 123.8226, 124.6089,
  35.39105, 36.17739, 36.97089, 37.7716, 38.57956, 39.39482, 40.21743, 
    41.04739, 41.88475, 42.72952, 43.58169, 44.44128, 45.30827, 46.18266, 
    47.0644, 47.95347, 48.84982, 49.75339, 50.66412, 51.58192, 52.50672, 
    53.43841, 54.37688, 55.32201, 56.27366, 57.23169, 58.19594, 59.16623, 
    60.14239, 61.12422, 62.11152, 63.10405, 64.10161, 65.10394, 66.1108, 
    67.12192, 68.13703, 69.15585, 70.17809, 71.20345, 72.23161, 73.26228, 
    74.29514, 75.32983, 76.36607, 77.40348, 78.44175, 79.48052, 80.51948, 
    81.55825, 82.59652, 83.63393, 84.67017, 85.70486, 86.73772, 87.76839, 
    88.79655, 89.82191, 90.84415, 91.86297, 92.87808, 93.8892, 94.89606, 
    95.89839, 96.89594, 97.88849, 98.87578, 99.8576, 100.8338, 101.8041, 
    102.7683, 103.7263, 104.678, 105.6231, 106.5616, 107.4933, 108.4181, 
    109.3359, 110.2466, 111.1502, 112.0465, 112.9356, 113.8173, 114.6917, 
    115.5587, 116.4183, 117.2705, 118.1152, 118.9526, 119.7826, 120.6052, 
    121.4204, 122.2284, 123.0291, 123.8226, 124.6089,
  35.39103, 36.17737, 36.97087, 37.77157, 38.57954, 39.3948, 40.2174, 
    41.04737, 41.88473, 42.72949, 43.58167, 44.44125, 45.30825, 46.18263, 
    47.06438, 47.95345, 48.84979, 49.75336, 50.66409, 51.5819, 52.5067, 
    53.43839, 54.37686, 55.32199, 56.27364, 57.23167, 58.19592, 59.16621, 
    60.14237, 61.1242, 62.1115, 63.10404, 64.10159, 65.10393, 66.11079, 
    67.12191, 68.13702, 69.15584, 70.17808, 71.20344, 72.23161, 73.26228, 
    74.29513, 75.32983, 76.36606, 77.40348, 78.44174, 79.48052, 80.51948, 
    81.55826, 82.59652, 83.63394, 84.67017, 85.70487, 86.73772, 87.76839, 
    88.79656, 89.82192, 90.84416, 91.86298, 92.87809, 93.88921, 94.89607, 
    95.89841, 96.89597, 97.8885, 98.8758, 99.85763, 100.8338, 101.8041, 
    102.7683, 103.7264, 104.678, 105.6231, 106.5616, 107.4933, 108.4181, 
    109.3359, 110.2466, 111.1502, 112.0466, 112.9356, 113.8174, 114.6917, 
    115.5587, 116.4183, 117.2705, 118.1153, 118.9526, 119.7826, 120.6052, 
    121.4205, 122.2284, 123.0291, 123.8226, 124.609,
  35.391, 36.17735, 36.97084, 37.77155, 38.57951, 39.39478, 40.21738, 
    41.04734, 41.8847, 42.72947, 43.58164, 44.44123, 45.30822, 46.18261, 
    47.06435, 47.95342, 48.84977, 49.75334, 50.66407, 51.58187, 52.50668, 
    53.43837, 54.37684, 55.32197, 56.27362, 57.23165, 58.1959, 59.16619, 
    60.14235, 61.12418, 62.11148, 63.10402, 64.10158, 65.10391, 66.11077, 
    67.12189, 68.137, 69.15582, 70.17806, 71.20342, 72.2316, 73.26227, 
    74.29512, 75.32983, 76.36606, 77.40347, 78.44174, 79.48052, 80.51948, 
    81.55826, 82.59653, 83.63394, 84.67017, 85.70488, 86.73773, 87.7684, 
    88.79658, 89.82194, 90.84418, 91.863, 92.87811, 93.88923, 94.89609, 
    95.89842, 96.89598, 97.88852, 98.87582, 99.85765, 100.8338, 101.8041, 
    102.7683, 103.7264, 104.678, 105.6232, 106.5616, 107.4933, 108.4181, 
    109.3359, 110.2467, 111.1502, 112.0466, 112.9356, 113.8174, 114.6918, 
    115.5588, 116.4184, 117.2705, 118.1153, 118.9527, 119.7826, 120.6052, 
    121.4205, 122.2285, 123.0292, 123.8227, 124.609,
  35.39098, 36.17732, 36.97082, 37.77152, 38.57949, 39.39475, 40.21735, 
    41.04732, 41.88467, 42.72944, 43.58162, 44.4412, 45.3082, 46.18258, 
    47.06433, 47.9534, 48.84974, 49.75331, 50.66404, 51.58185, 52.50665, 
    53.43834, 54.37682, 55.32195, 56.2736, 57.23163, 58.19588, 59.16617, 
    60.14233, 61.12416, 62.11146, 63.104, 64.10156, 65.1039, 66.11076, 
    67.12188, 68.13699, 69.15582, 70.17805, 71.20341, 72.23159, 73.26226, 
    74.29511, 75.32982, 76.36605, 77.40347, 78.44174, 79.48052, 80.51948, 
    81.55826, 82.59653, 83.63395, 84.67018, 85.70489, 86.73774, 87.76841, 
    88.79659, 89.82195, 90.84418, 91.86301, 92.87812, 93.88924, 94.8961, 
    95.89844, 96.896, 97.88854, 98.87583, 99.85767, 100.8338, 101.8041, 
    102.7684, 103.7264, 104.6781, 105.6232, 106.5617, 107.4933, 108.4182, 
    109.336, 110.2467, 111.1503, 112.0466, 112.9357, 113.8174, 114.6918, 
    115.5588, 116.4184, 117.2706, 118.1153, 118.9527, 119.7826, 120.6052, 
    121.4205, 122.2285, 123.0292, 123.8227, 124.609,
  35.39095, 36.1773, 36.97079, 37.7715, 38.57946, 39.39472, 40.21732, 
    41.04729, 41.88465, 42.72941, 43.58159, 44.44118, 45.30817, 46.18256, 
    47.0643, 47.95337, 48.84972, 49.75329, 50.66402, 51.58183, 52.50663, 
    53.43832, 54.37679, 55.32192, 56.27357, 57.23161, 58.19585, 59.16615, 
    60.14231, 61.12415, 62.11144, 63.10398, 64.10155, 65.10388, 66.11074, 
    67.12186, 68.13698, 69.1558, 70.17805, 71.20341, 72.23158, 73.26225, 
    74.29511, 75.32982, 76.36605, 77.40347, 78.44174, 79.48052, 80.51948, 
    81.55826, 82.59653, 83.63395, 84.67018, 85.70489, 86.73775, 87.76842, 
    88.79659, 89.82195, 90.8442, 91.86302, 92.87814, 93.88926, 94.89612, 
    95.89845, 96.89601, 97.88856, 98.87585, 99.85769, 100.8338, 101.8041, 
    102.7684, 103.7264, 104.6781, 105.6232, 106.5617, 107.4934, 108.4182, 
    109.336, 110.2467, 111.1503, 112.0466, 112.9357, 113.8174, 114.6918, 
    115.5588, 116.4184, 117.2706, 118.1153, 118.9527, 119.7827, 120.6053, 
    121.4205, 122.2285, 123.0292, 123.8227, 124.609,
  35.39093, 36.17727, 36.97076, 37.77147, 38.57943, 39.3947, 40.2173, 
    41.04726, 41.88462, 42.72939, 43.58156, 44.44115, 45.30815, 46.18253, 
    47.06427, 47.95334, 48.84969, 49.75326, 50.66399, 51.5818, 52.5066, 
    53.43829, 54.37677, 55.3219, 56.27355, 57.23158, 58.19584, 59.16613, 
    60.14229, 61.12413, 62.11142, 63.10397, 64.10153, 65.10387, 66.11073, 
    67.12185, 68.13696, 69.15579, 70.17803, 71.20339, 72.23158, 73.26225, 
    74.2951, 75.32981, 76.36604, 77.40347, 78.44173, 79.48052, 80.51948, 
    81.55827, 82.59653, 83.63396, 84.67019, 85.7049, 86.73775, 87.76842, 
    88.79661, 89.82197, 90.84421, 91.86304, 92.87815, 93.88927, 94.89613, 
    95.89847, 96.89603, 97.88857, 98.87587, 99.8577, 100.8339, 101.8042, 
    102.7684, 103.7264, 104.6781, 105.6232, 106.5617, 107.4934, 108.4182, 
    109.336, 110.2467, 111.1503, 112.0467, 112.9357, 113.8175, 114.6919, 
    115.5588, 116.4184, 117.2706, 118.1154, 118.9527, 119.7827, 120.6053, 
    121.4206, 122.2285, 123.0292, 123.8227, 124.6091,
  35.3909, 36.17724, 36.97074, 37.77145, 38.57941, 39.39467, 40.21727, 
    41.04724, 41.88459, 42.72936, 43.58154, 44.44112, 45.30812, 46.1825, 
    47.06425, 47.95332, 48.84967, 49.75324, 50.66397, 51.58178, 52.50658, 
    53.43827, 54.37674, 55.32187, 56.27353, 57.23156, 58.19581, 59.16611, 
    60.14227, 61.12411, 62.1114, 63.10395, 64.10151, 65.10385, 66.11071, 
    67.12183, 68.13696, 69.15578, 70.17802, 71.20338, 72.23156, 73.26224, 
    74.2951, 75.3298, 76.36604, 77.40347, 78.44173, 79.48052, 80.51948, 
    81.55827, 82.59653, 83.63396, 84.6702, 85.7049, 86.73776, 87.76844, 
    88.79662, 89.82198, 90.84422, 91.86304, 92.87817, 93.88929, 94.89615, 
    95.89849, 96.89605, 97.8886, 98.87589, 99.85773, 100.8339, 101.8042, 
    102.7684, 103.7265, 104.6781, 105.6233, 106.5617, 107.4934, 108.4182, 
    109.336, 110.2468, 111.1503, 112.0467, 112.9358, 113.8175, 114.6919, 
    115.5589, 116.4185, 117.2706, 118.1154, 118.9528, 119.7827, 120.6053, 
    121.4206, 122.2286, 123.0293, 123.8228, 124.6091,
  35.39088, 36.17722, 36.97071, 37.77142, 38.57938, 39.39464, 40.21724, 
    41.04721, 41.88457, 42.72933, 43.58151, 44.4411, 45.30809, 46.18248, 
    47.06422, 47.95329, 48.84964, 49.75321, 50.66394, 51.58175, 52.50655, 
    53.43824, 54.37672, 55.32185, 56.27351, 57.23154, 58.19579, 59.16609, 
    60.14225, 61.12409, 62.11139, 63.10393, 64.10149, 65.10384, 66.11069, 
    67.12183, 68.13694, 69.15577, 70.17801, 71.20338, 72.23155, 73.26223, 
    74.29509, 75.3298, 76.36604, 77.40346, 78.44173, 79.48052, 80.51948, 
    81.55827, 82.59654, 83.63396, 84.6702, 85.70491, 86.73777, 87.76845, 
    88.79662, 89.82199, 90.84423, 91.86306, 92.87817, 93.88931, 94.89616, 
    95.89851, 96.89606, 97.88861, 98.87592, 99.85775, 100.8339, 101.8042, 
    102.7685, 103.7265, 104.6781, 105.6233, 106.5618, 107.4934, 108.4183, 
    109.3361, 110.2468, 111.1504, 112.0467, 112.9358, 113.8175, 114.6919, 
    115.5589, 116.4185, 117.2707, 118.1154, 118.9528, 119.7828, 120.6054, 
    121.4206, 122.2286, 123.0293, 123.8228, 124.6091,
  35.39085, 36.17719, 36.97068, 37.77139, 38.57935, 39.39462, 40.21722, 
    41.04718, 41.88454, 42.7293, 43.58148, 44.44107, 45.30806, 46.18245, 
    47.06419, 47.95326, 48.84961, 49.75319, 50.66391, 51.58173, 52.50653, 
    53.43822, 54.37669, 55.32183, 56.27348, 57.23152, 58.19577, 59.16607, 
    60.14223, 61.12407, 62.11137, 63.10391, 64.10148, 65.10381, 66.11068, 
    67.12181, 68.13692, 69.15575, 70.178, 71.20337, 72.23154, 73.26222, 
    74.29508, 75.3298, 76.36603, 77.40346, 78.44173, 79.48052, 80.51948, 
    81.55827, 82.59654, 83.63397, 84.6702, 85.70492, 86.73778, 87.76846, 
    88.79663, 89.822, 90.84425, 91.86308, 92.87819, 93.88932, 94.89619, 
    95.89852, 96.89609, 97.88863, 98.87593, 99.85777, 100.8339, 101.8042, 
    102.7685, 103.7265, 104.6782, 105.6233, 106.5618, 107.4935, 108.4183, 
    109.3361, 110.2468, 111.1504, 112.0467, 112.9358, 113.8176, 114.6919, 
    115.5589, 116.4185, 117.2707, 118.1155, 118.9528, 119.7828, 120.6054, 
    121.4206, 122.2286, 123.0293, 123.8228, 124.6092,
  35.39082, 36.17716, 36.97066, 37.77136, 38.57932, 39.39459, 40.21719, 
    41.04715, 41.88451, 42.72927, 43.58145, 44.44104, 45.30804, 46.18242, 
    47.06416, 47.95324, 48.84959, 49.75316, 50.66389, 51.5817, 52.5065, 
    53.43819, 54.37667, 55.3218, 56.27346, 57.23149, 58.19575, 59.16605, 
    60.14221, 61.12405, 62.11135, 63.1039, 64.10146, 65.1038, 66.11066, 
    67.1218, 68.13691, 69.15574, 70.17799, 71.20335, 72.23154, 73.26221, 
    74.29507, 75.32979, 76.36603, 77.40345, 78.44173, 79.48052, 80.51948, 
    81.55827, 82.59655, 83.63397, 84.67021, 85.70493, 86.73779, 87.76846, 
    88.79665, 89.82201, 90.84426, 91.86309, 92.8782, 93.88934, 94.8962, 
    95.89854, 96.8961, 97.88865, 98.87595, 99.85779, 100.834, 101.8043, 
    102.7685, 103.7265, 104.6782, 105.6233, 106.5618, 107.4935, 108.4183, 
    109.3361, 110.2468, 111.1504, 112.0468, 112.9358, 113.8176, 114.692, 
    115.559, 116.4185, 117.2707, 118.1155, 118.9528, 119.7828, 120.6054, 
    121.4207, 122.2286, 123.0293, 123.8228, 124.6092,
  35.39079, 36.17713, 36.97063, 37.77133, 38.5793, 39.39456, 40.21716, 
    41.04713, 41.88448, 42.72924, 43.58142, 44.44101, 45.30801, 46.18239, 
    47.06414, 47.95321, 48.84956, 49.75313, 50.66386, 51.58167, 52.50647, 
    53.43817, 54.37664, 55.32178, 56.27344, 57.23147, 58.19572, 59.16602, 
    60.14219, 61.12403, 62.11133, 63.10388, 64.10144, 65.10378, 66.11065, 
    67.12178, 68.1369, 69.15573, 70.17798, 71.20335, 72.23153, 73.26221, 
    74.29507, 75.32978, 76.36602, 77.40345, 78.44173, 79.48052, 80.51948, 
    81.55827, 82.59655, 83.63398, 84.67022, 85.70493, 86.73779, 87.76847, 
    88.79665, 89.82202, 90.84427, 91.8631, 92.87822, 93.88935, 94.89622, 
    95.89856, 96.89613, 97.88867, 98.87597, 99.85781, 100.834, 101.8043, 
    102.7685, 103.7266, 104.6782, 105.6234, 106.5618, 107.4935, 108.4183, 
    109.3361, 110.2469, 111.1504, 112.0468, 112.9359, 113.8176, 114.692, 
    115.559, 116.4186, 117.2708, 118.1155, 118.9529, 119.7828, 120.6054, 
    121.4207, 122.2287, 123.0294, 123.8229, 124.6092,
  35.39077, 36.1771, 36.9706, 37.77131, 38.57927, 39.39453, 40.21713, 
    41.0471, 41.88445, 42.72922, 43.58139, 44.44098, 45.30798, 46.18237, 
    47.06411, 47.95318, 48.84953, 49.75311, 50.66383, 51.58165, 52.50645, 
    53.43814, 54.37662, 55.32175, 56.27341, 57.23145, 58.1957, 59.166, 
    60.14217, 61.12401, 62.11131, 63.10386, 64.10143, 65.10377, 66.11063, 
    67.12177, 68.13689, 69.15572, 70.17796, 71.20334, 72.23152, 73.2622, 
    74.29506, 75.32978, 76.36602, 77.40345, 78.44173, 79.48052, 80.51948, 
    81.55827, 82.59655, 83.63398, 84.67022, 85.70494, 86.7378, 87.76848, 
    88.79666, 89.82204, 90.84428, 91.86311, 92.87823, 93.88937, 94.89623, 
    95.89857, 96.89614, 97.88869, 98.87599, 99.85783, 100.834, 101.8043, 
    102.7686, 103.7266, 104.6782, 105.6234, 106.5619, 107.4936, 108.4184, 
    109.3362, 110.2469, 111.1505, 112.0468, 112.9359, 113.8176, 114.692, 
    115.559, 116.4186, 117.2708, 118.1155, 118.9529, 119.7829, 120.6055, 
    121.4207, 122.2287, 123.0294, 123.8229, 124.6092,
  35.39074, 36.17707, 36.97057, 37.77127, 38.57924, 39.3945, 40.2171, 
    41.04707, 41.88443, 42.72919, 43.58136, 44.44096, 45.30795, 46.18233, 
    47.06408, 47.95315, 48.8495, 49.75307, 50.66381, 51.58162, 52.50642, 
    53.43812, 54.37659, 55.32173, 56.27339, 57.23142, 58.19568, 59.16598, 
    60.14215, 61.12399, 62.11129, 63.10384, 64.10141, 65.10375, 66.11062, 
    67.12175, 68.13687, 69.1557, 70.17796, 71.20332, 72.23151, 73.26219, 
    74.29506, 75.32977, 76.36601, 77.40344, 78.44173, 79.48051, 80.51949, 
    81.55827, 82.59656, 83.63399, 84.67023, 85.70494, 86.73781, 87.76849, 
    88.79668, 89.82204, 90.8443, 91.86313, 92.87825, 93.88938, 94.89625, 
    95.89859, 96.89616, 97.88871, 98.87601, 99.85785, 100.834, 101.8043, 
    102.7686, 103.7266, 104.6783, 105.6234, 106.5619, 107.4936, 108.4184, 
    109.3362, 110.2469, 111.1505, 112.0469, 112.9359, 113.8177, 114.692, 
    115.559, 116.4186, 117.2708, 118.1156, 118.9529, 119.7829, 120.6055, 
    121.4208, 122.2287, 123.0294, 123.8229, 124.6093,
  35.39071, 36.17704, 36.97054, 37.77124, 38.57921, 39.39447, 40.21707, 
    41.04704, 41.8844, 42.72916, 43.58134, 44.44093, 45.30792, 46.1823, 
    47.06405, 47.95312, 48.84948, 49.75305, 50.66378, 51.58159, 52.5064, 
    53.43809, 54.37657, 55.3217, 56.27337, 57.2314, 58.19566, 59.16596, 
    60.14213, 61.12397, 62.11127, 63.10382, 64.10139, 65.10374, 66.1106, 
    67.12173, 68.13686, 69.15569, 70.17794, 71.20332, 72.2315, 73.26218, 
    74.29505, 75.32977, 76.36601, 77.40344, 78.44173, 79.48051, 80.51949, 
    81.55827, 82.59656, 83.63399, 84.67023, 85.70495, 86.73782, 87.7685, 
    88.79668, 89.82206, 90.84431, 91.86314, 92.87827, 93.8894, 94.89626, 
    95.89861, 96.89618, 97.88873, 98.87603, 99.85787, 100.834, 101.8043, 
    102.7686, 103.7266, 104.6783, 105.6234, 106.5619, 107.4936, 108.4184, 
    109.3362, 110.2469, 111.1505, 112.0469, 112.936, 113.8177, 114.6921, 
    115.5591, 116.4187, 117.2708, 118.1156, 118.953, 119.7829, 120.6055, 
    121.4208, 122.2288, 123.0295, 123.823, 124.6093,
  35.39067, 36.17702, 36.97051, 37.77121, 38.57918, 39.39444, 40.21704, 
    41.04701, 41.88437, 42.72913, 43.58131, 44.4409, 45.30789, 46.18228, 
    47.06402, 47.95309, 48.84945, 49.75302, 50.66375, 51.58157, 52.50637, 
    53.43807, 54.37654, 55.32168, 56.27334, 57.23138, 58.19563, 59.16594, 
    60.14211, 61.12395, 62.11125, 63.10381, 64.10137, 65.10372, 66.11059, 
    67.12172, 68.13685, 69.15568, 70.17793, 71.20331, 72.23149, 73.26218, 
    74.29504, 75.32977, 76.366, 77.40343, 78.44172, 79.48051, 80.51949, 
    81.55828, 82.59657, 83.634, 84.67023, 85.70496, 86.73782, 87.76851, 
    88.79669, 89.82207, 90.84432, 91.86315, 92.87828, 93.88941, 94.89628, 
    95.89863, 96.89619, 97.88875, 98.87605, 99.85789, 100.8341, 101.8044, 
    102.7686, 103.7267, 104.6783, 105.6235, 106.5619, 107.4936, 108.4184, 
    109.3362, 110.247, 111.1506, 112.0469, 112.936, 113.8177, 114.6921, 
    115.5591, 116.4187, 117.2709, 118.1156, 118.953, 119.783, 120.6056, 
    121.4208, 122.2288, 123.0295, 123.823, 124.6093,
  35.39064, 36.17699, 36.97048, 37.77118, 38.57915, 39.39441, 40.21701, 
    41.04698, 41.88433, 42.7291, 43.58128, 44.44087, 45.30787, 46.18225, 
    47.064, 47.95307, 48.84942, 49.75299, 50.66373, 51.58154, 52.50634, 
    53.43804, 54.37652, 55.32166, 56.27332, 57.23135, 58.19561, 59.16592, 
    60.14209, 61.12393, 62.11123, 63.10379, 64.10136, 65.1037, 66.11057, 
    67.1217, 68.13683, 69.15567, 70.17793, 71.20329, 72.23148, 73.26217, 
    74.29504, 75.32976, 76.366, 77.40343, 78.44172, 79.48051, 80.51949, 
    81.55828, 82.59657, 83.634, 84.67024, 85.70496, 86.73783, 87.76852, 
    88.79671, 89.82207, 90.84433, 91.86317, 92.8783, 93.88943, 94.8963, 
    95.89864, 96.89622, 97.88876, 98.87608, 99.85791, 100.8341, 101.8044, 
    102.7686, 103.7267, 104.6783, 105.6235, 106.562, 107.4937, 108.4185, 
    109.3363, 110.247, 111.1506, 112.0469, 112.936, 113.8177, 114.6921, 
    115.5591, 116.4187, 117.2709, 118.1157, 118.953, 119.783, 120.6056, 
    121.4209, 122.2288, 123.0295, 123.823, 124.6094,
  35.39061, 36.17695, 36.97045, 37.77115, 38.57912, 39.39438, 40.21698, 
    41.04695, 41.8843, 42.72907, 43.58125, 44.44084, 45.30783, 46.18222, 
    47.06396, 47.95304, 48.84939, 49.75296, 50.6637, 51.58151, 52.50632, 
    53.43801, 54.3765, 55.32163, 56.27329, 57.23133, 58.19559, 59.16589, 
    60.14207, 61.12391, 62.11121, 63.10377, 64.10134, 65.10368, 66.11056, 
    67.1217, 68.13682, 69.15565, 70.17791, 71.20329, 72.23148, 73.26216, 
    74.29503, 75.32975, 76.366, 77.40343, 78.44172, 79.48051, 80.51949, 
    81.55828, 82.59657, 83.634, 84.67025, 85.70497, 86.73784, 87.76852, 
    88.79671, 89.82209, 90.84435, 91.86318, 92.8783, 93.88944, 94.89632, 
    95.89866, 96.89623, 97.88879, 98.87609, 99.85793, 100.8341, 101.8044, 
    102.7687, 103.7267, 104.6784, 105.6235, 106.562, 107.4937, 108.4185, 
    109.3363, 110.247, 111.1506, 112.047, 112.936, 113.8178, 114.6922, 
    115.5592, 116.4188, 117.2709, 118.1157, 118.9531, 119.783, 120.6056, 
    121.4209, 122.2288, 123.0295, 123.823, 124.6094,
  35.39058, 36.17692, 36.97042, 37.77112, 38.57908, 39.39435, 40.21695, 
    41.04692, 41.88427, 42.72904, 43.58121, 44.44081, 45.3078, 46.18219, 
    47.06393, 47.95301, 48.84936, 49.75294, 50.66367, 51.58149, 52.50629, 
    53.43799, 54.37647, 55.32161, 56.27327, 57.23131, 58.19557, 59.16587, 
    60.14204, 61.12389, 62.11119, 63.10375, 64.10132, 65.10367, 66.11054, 
    67.12168, 68.1368, 69.15564, 70.1779, 71.20328, 72.23147, 73.26215, 
    74.29502, 75.32975, 76.36599, 77.40343, 78.44172, 79.48051, 80.51949, 
    81.55828, 82.59657, 83.63401, 84.67025, 85.70498, 86.73785, 87.76853, 
    88.79672, 89.8221, 90.84436, 91.8632, 92.87832, 93.88946, 94.89633, 
    95.89868, 96.89625, 97.8888, 98.87611, 99.85796, 100.8341, 101.8044, 
    102.7687, 103.7267, 104.6784, 105.6235, 106.562, 107.4937, 108.4185, 
    109.3363, 110.2471, 111.1506, 112.047, 112.9361, 113.8178, 114.6922, 
    115.5592, 116.4188, 117.271, 118.1157, 118.9531, 119.7831, 120.6057, 
    121.4209, 122.2289, 123.0296, 123.8231, 124.6094,
  35.39055, 36.17689, 36.97039, 37.77109, 38.57905, 39.39432, 40.21692, 
    41.04689, 41.88424, 42.72901, 43.58118, 44.44078, 45.30777, 46.18216, 
    47.06391, 47.95298, 48.84933, 49.75291, 50.66364, 51.58146, 52.50626, 
    53.43797, 54.37645, 55.32158, 56.27325, 57.23129, 58.19555, 59.16585, 
    60.14202, 61.12387, 62.11118, 63.10373, 64.1013, 65.10365, 66.11053, 
    67.12167, 68.1368, 69.15563, 70.17789, 71.20326, 72.23145, 73.26215, 
    74.29501, 75.32974, 76.36599, 77.40343, 78.44171, 79.48051, 80.51949, 
    81.55829, 82.59657, 83.63401, 84.67026, 85.70499, 86.73785, 87.76855, 
    88.79674, 89.82211, 90.84437, 91.8632, 92.87833, 93.88947, 94.89635, 
    95.8987, 96.89627, 97.88882, 98.87613, 99.85798, 100.8342, 101.8045, 
    102.7687, 103.7268, 104.6784, 105.6236, 106.562, 107.4937, 108.4185, 
    109.3364, 110.2471, 111.1507, 112.047, 112.9361, 113.8178, 114.6922, 
    115.5592, 116.4188, 117.271, 118.1158, 118.9531, 119.7831, 120.6057, 
    121.4209, 122.2289, 123.0296, 123.8231, 124.6095,
  35.39052, 36.17686, 36.97036, 37.77106, 38.57902, 39.39428, 40.21688, 
    41.04685, 41.88421, 42.72898, 43.58115, 44.44075, 45.30774, 46.18213, 
    47.06388, 47.95295, 48.8493, 49.75288, 50.66362, 51.58143, 52.50624, 
    53.43794, 54.37642, 55.32156, 56.27322, 57.23126, 58.19552, 59.16583, 
    60.142, 61.12385, 62.11116, 63.10371, 64.10129, 65.10364, 66.11051, 
    67.12165, 68.13678, 69.15562, 70.17788, 71.20325, 72.23145, 73.26214, 
    74.29501, 75.32973, 76.36598, 77.40342, 78.44171, 79.48051, 80.51949, 
    81.55829, 82.59658, 83.63402, 84.67027, 85.70499, 86.73786, 87.76855, 
    88.79675, 89.82212, 90.84438, 91.86322, 92.87835, 93.88949, 94.89636, 
    95.89871, 96.89629, 97.88884, 98.87615, 99.85799, 100.8342, 101.8045, 
    102.7687, 103.7268, 104.6784, 105.6236, 106.5621, 107.4938, 108.4186, 
    109.3364, 110.2471, 111.1507, 112.0471, 112.9361, 113.8179, 114.6923, 
    115.5592, 116.4188, 117.271, 118.1158, 118.9531, 119.7831, 120.6057, 
    121.421, 122.2289, 123.0296, 123.8231, 124.6095 ;

 grid_latt =
  -35.07925, -35.43988, -35.79544, -36.14578, -36.4908, -36.83038, -37.1644, 
    -37.49273, -37.81525, -38.13184, -38.44237, -38.74672, -39.04476, 
    -39.33637, -39.62142, -39.89979, -40.17135, -40.43598, -40.69355, 
    -40.94394, -41.18702, -41.42268, -41.65079, -41.87124, -42.08391, 
    -42.28868, -42.48545, -42.67411, -42.85454, -43.02665, -43.19033, 
    -43.34549, -43.49203, -43.62987, -43.75893, -43.87911, -43.99035, 
    -44.09258, -44.18572, -44.26973, -44.34454, -44.41011, -44.46639, 
    -44.51335, -44.55096, -44.57919, -44.59801, -44.60743, -44.60743, 
    -44.59801, -44.57919, -44.55096, -44.51335, -44.46639, -44.41011, 
    -44.34454, -44.26973, -44.18572, -44.09258, -43.99035, -43.87911, 
    -43.75893, -43.62987, -43.49203, -43.34549, -43.19033, -43.02665, 
    -42.85454, -42.67411, -42.48545, -42.28868, -42.08391, -41.87124, 
    -41.65079, -41.42268, -41.18702, -40.94394, -40.69355, -40.43598, 
    -40.17135, -39.89979, -39.62142, -39.33637, -39.04476, -38.74672, 
    -38.44237, -38.13184, -37.81525, -37.49273, -37.1644, -36.83038, 
    -36.4908, -36.14578, -35.79544, -35.43988, -35.07925,
  -34.34282, -34.70005, -35.05236, -35.39962, -35.7417, -36.0785, -36.40988, 
    -36.73572, -37.05589, -37.37026, -37.67871, -37.9811, -38.27731, 
    -38.56721, -38.85067, -39.12755, -39.39772, -39.66107, -39.91746, 
    -40.16676, -40.40884, -40.64358, -40.87085, -41.09053, -41.30251, 
    -41.50666, -41.70287, -41.89101, -42.07099, -42.24269, -42.40602, 
    -42.56086, -42.70713, -42.84472, -42.97356, -43.09357, -43.20465, 
    -43.30674, -43.39978, -43.48369, -43.55843, -43.62393, -43.68016, 
    -43.72708, -43.76466, -43.79286, -43.81168, -43.82109, -43.82109, 
    -43.81168, -43.79286, -43.76466, -43.72708, -43.68016, -43.62393, 
    -43.55843, -43.48369, -43.39978, -43.30674, -43.20465, -43.09357, 
    -42.97356, -42.84472, -42.70713, -42.56086, -42.40602, -42.24269, 
    -42.07099, -41.89101, -41.70287, -41.50666, -41.30251, -41.09053, 
    -40.87085, -40.64358, -40.40884, -40.16676, -39.91746, -39.66107, 
    -39.39772, -39.12755, -38.85067, -38.56721, -38.27731, -37.9811, 
    -37.67871, -37.37026, -37.05589, -36.73572, -36.40988, -36.0785, 
    -35.7417, -35.39962, -35.05236, -34.70005, -34.34282,
  -33.60628, -33.95987, -34.30869, -34.65261, -34.99154, -35.32531, 
    -35.65382, -35.97694, -36.29453, -36.60646, -36.91259, -37.21281, 
    -37.50697, -37.79493, -38.07658, -38.35176, -38.62035, -38.88222, 
    -39.13723, -39.38524, -39.62614, -39.85978, -40.08604, -40.30479, 
    -40.51591, -40.71927, -40.91476, -41.10225, -41.28164, -41.4528, 
    -41.61564, -41.77005, -41.91592, -42.05317, -42.18171, -42.30143, 
    -42.41228, -42.51416, -42.60701, -42.69076, -42.76536, -42.83075, 
    -42.88689, -42.93373, -42.97124, -42.9994, -43.01819, -43.02758, 
    -43.02758, -43.01819, -42.9994, -42.97124, -42.93373, -42.88689, 
    -42.83075, -42.76536, -42.69076, -42.60701, -42.51416, -42.41228, 
    -42.30143, -42.18171, -42.05317, -41.91592, -41.77005, -41.61564, 
    -41.4528, -41.28164, -41.10225, -40.91476, -40.71927, -40.51591, 
    -40.30479, -40.08604, -39.85978, -39.62614, -39.38524, -39.13723, 
    -38.88222, -38.62035, -38.35176, -38.07658, -37.79493, -37.50697, 
    -37.21281, -36.91259, -36.60646, -36.29453, -35.97694, -35.65382, 
    -35.32531, -34.99154, -34.65261, -34.30869, -33.95987, -33.60628,
  -32.86962, -33.21932, -33.56442, -33.90479, -34.2403, -34.57083, -34.89624, 
    -35.2164, -35.53117, -35.84042, -36.14403, -36.44184, -36.73372, 
    -37.01954, -37.29916, -37.57244, -37.83924, -38.09942, -38.35286, 
    -38.5994, -38.83891, -39.07127, -39.29634, -39.51399, -39.72409, 
    -39.9265, -40.12112, -40.30781, -40.48646, -40.65696, -40.81918, 
    -40.97303, -41.1184, -41.25519, -41.38331, -41.50267, -41.61318, 
    -41.71477, -41.80736, -41.89089, -41.96529, -42.03052, -42.08652, 
    -42.13324, -42.17067, -42.19876, -42.2175, -42.22688, -42.22688, 
    -42.2175, -42.19876, -42.17067, -42.13324, -42.08652, -42.03052, 
    -41.96529, -41.89089, -41.80736, -41.71477, -41.61318, -41.50267, 
    -41.38331, -41.25519, -41.1184, -40.97303, -40.81918, -40.65696, 
    -40.48646, -40.30781, -40.12112, -39.9265, -39.72409, -39.51399, 
    -39.29634, -39.07127, -38.83891, -38.5994, -38.35286, -38.09942, 
    -37.83924, -37.57244, -37.29916, -37.01954, -36.73372, -36.44184, 
    -36.14403, -35.84042, -35.53117, -35.2164, -34.89624, -34.57083, 
    -34.2403, -33.90479, -33.56442, -33.21932, -32.86962,
  -32.13284, -32.47842, -32.81957, -33.15614, -33.48802, -33.81506, 
    -34.13713, -34.4541, -34.76583, -35.07218, -35.37302, -35.66821, 
    -35.9576, -36.24105, -36.51843, -36.78959, -37.05439, -37.31269, 
    -37.56434, -37.80922, -38.04717, -38.27806, -38.50176, -38.71813, 
    -38.92703, -39.12834, -39.32193, -39.50767, -39.68544, -39.85512, 
    -40.0166, -40.16977, -40.31451, -40.45074, -40.57834, -40.69724, 
    -40.80733, -40.90854, -41.0008, -41.08404, -41.15818, -41.22319, -41.279, 
    -41.32558, -41.36288, -41.39089, -41.40957, -41.41891, -41.41891, 
    -41.40957, -41.39089, -41.36288, -41.32558, -41.279, -41.22319, 
    -41.15818, -41.08404, -41.0008, -40.90854, -40.80733, -40.69724, 
    -40.57834, -40.45074, -40.31451, -40.16977, -40.0166, -39.85512, 
    -39.68544, -39.50767, -39.32193, -39.12834, -38.92703, -38.71813, 
    -38.50176, -38.27806, -38.04717, -37.80922, -37.56434, -37.31269, 
    -37.05439, -36.78959, -36.51843, -36.24105, -35.9576, -35.66821, 
    -35.37302, -35.07218, -34.76583, -34.4541, -34.13713, -33.81506, 
    -33.48802, -33.15614, -32.81957, -32.47842, -32.13284,
  -31.39594, -31.73718, -32.07414, -32.40669, -32.73469, -33.05801, 
    -33.37651, -33.69006, -33.99852, -34.30174, -34.59959, -34.89193, 
    -35.1786, -35.45947, -35.73439, -36.00322, -36.26581, -36.52202, 
    -36.7717, -37.01471, -37.2509, -37.48015, -37.70229, -37.9172, -38.12474, 
    -38.32478, -38.51718, -38.70182, -38.87856, -39.04729, -39.20789, 
    -39.36025, -39.50425, -39.63979, -39.76678, -39.88511, -39.99469, 
    -40.09544, -40.18729, -40.27016, -40.34399, -40.40873, -40.46431, 
    -40.51069, -40.54784, -40.57574, -40.59435, -40.60365, -40.60365, 
    -40.59435, -40.57574, -40.54784, -40.51069, -40.46431, -40.40873, 
    -40.34399, -40.27016, -40.18729, -40.09544, -39.99469, -39.88511, 
    -39.76678, -39.63979, -39.50425, -39.36025, -39.20789, -39.04729, 
    -38.87856, -38.70182, -38.51718, -38.32478, -38.12474, -37.9172, 
    -37.70229, -37.48015, -37.2509, -37.01471, -36.7717, -36.52202, 
    -36.26581, -36.00322, -35.73439, -35.45947, -35.1786, -34.89193, 
    -34.59959, -34.30174, -33.99852, -33.69006, -33.37651, -33.05801, 
    -32.73469, -32.40669, -32.07414, -31.73718, -31.39594,
  -30.65893, -30.9956, -31.32814, -31.65643, -31.98032, -32.29969, -32.6144, 
    -32.9243, -33.22925, -33.52912, -33.82376, -34.11302, -34.39675, 
    -34.67482, -34.94707, -35.21335, -35.47353, -35.72744, -35.97494, 
    -36.21589, -36.45013, -36.67753, -36.89794, -37.11122, -37.31722, 
    -37.51582, -37.70687, -37.89024, -38.06581, -38.23346, -38.39304, 
    -38.54446, -38.6876, -38.82234, -38.94859, -39.06625, -39.17523, 
    -39.27544, -39.3668, -39.44924, -39.52269, -39.58709, -39.6424, 
    -39.68855, -39.72552, -39.75327, -39.77179, -39.78105, -39.78105, 
    -39.77179, -39.75327, -39.72552, -39.68855, -39.6424, -39.58709, 
    -39.52269, -39.44924, -39.3668, -39.27544, -39.17523, -39.06625, 
    -38.94859, -38.82234, -38.6876, -38.54446, -38.39304, -38.23346, 
    -38.06581, -37.89024, -37.70687, -37.51582, -37.31722, -37.11122, 
    -36.89794, -36.67753, -36.45013, -36.21589, -35.97494, -35.72744, 
    -35.47353, -35.21335, -34.94707, -34.67482, -34.39675, -34.11302, 
    -33.82376, -33.52912, -33.22925, -32.9243, -32.6144, -32.29969, 
    -31.98032, -31.65643, -31.32814, -30.9956, -30.65893,
  -29.92181, -30.25368, -30.58158, -30.90537, -31.22494, -31.54013, -31.8508, 
    -32.15683, -32.45805, -32.75434, -33.04553, -33.33149, -33.61207, 
    -33.88711, -34.15647, -34.42, -34.67754, -34.92895, -35.17407, -35.41275, 
    -35.64485, -35.87022, -36.08871, -36.30017, -36.50447, -36.70145, 
    -36.891, -37.07295, -37.2472, -37.4136, -37.57203, -37.72238, -37.86452, 
    -37.99836, -38.12377, -38.24066, -38.34894, -38.44851, -38.53931, 
    -38.62124, -38.69425, -38.75827, -38.81324, -38.85912, -38.89588, 
    -38.92347, -38.94188, -38.95109, -38.95109, -38.94188, -38.92347, 
    -38.89588, -38.85912, -38.81324, -38.75827, -38.69425, -38.62124, 
    -38.53931, -38.44851, -38.34894, -38.24066, -38.12377, -37.99836, 
    -37.86452, -37.72238, -37.57203, -37.4136, -37.2472, -37.07295, -36.891, 
    -36.70145, -36.50447, -36.30017, -36.08871, -35.87022, -35.64485, 
    -35.41275, -35.17407, -34.92895, -34.67754, -34.42, -34.15647, -33.88711, 
    -33.61207, -33.33149, -33.04553, -32.75434, -32.45805, -32.15683, 
    -31.8508, -31.54013, -31.22494, -30.90537, -30.58158, -30.25368, -29.92181,
  -29.18457, -29.51142, -29.83445, -30.15354, -30.46854, -30.77932, 
    -31.08575, -31.38766, -31.68493, -31.97741, -32.26494, -32.54737, 
    -32.82457, -33.09637, -33.36263, -33.62318, -33.87788, -34.12658, 
    -34.36911, -34.60533, -34.83509, -35.05824, -35.27462, -35.48409, 
    -35.68649, -35.8817, -36.06956, -36.24994, -36.42271, -36.58773, 
    -36.74487, -36.89401, -37.03504, -37.16784, -37.2923, -37.40832, 
    -37.5158, -37.61465, -37.7048, -37.78615, -37.85865, -37.92222, 
    -37.97682, -38.02239, -38.0589, -38.0863, -38.10459, -38.11374, 
    -38.11374, -38.10459, -38.0863, -38.0589, -38.02239, -37.97682, 
    -37.92222, -37.85865, -37.78615, -37.7048, -37.61465, -37.5158, 
    -37.40832, -37.2923, -37.16784, -37.03504, -36.89401, -36.74487, 
    -36.58773, -36.42271, -36.24994, -36.06956, -35.8817, -35.68649, 
    -35.48409, -35.27462, -35.05824, -34.83509, -34.60533, -34.36911, 
    -34.12658, -33.87788, -33.62318, -33.36263, -33.09637, -32.82457, 
    -32.54737, -32.26494, -31.97741, -31.68493, -31.38766, -31.08575, 
    -30.77932, -30.46854, -30.15354, -29.83445, -29.51142, -29.18457,
  -28.44723, -28.76883, -29.08677, -29.40093, -29.71115, -30.0173, -30.31924, 
    -30.61683, -30.90992, -31.19835, -31.482, -31.76069, -32.03428, 
    -32.30262, -32.56555, -32.82292, -33.07457, -33.32034, -33.56009, 
    -33.79364, -34.02087, -34.2416, -34.45568, -34.66297, -34.86331, 
    -35.05656, -35.24258, -35.42123, -35.59236, -35.75585, -35.91155, 
    -36.05936, -36.19914, -36.33079, -36.45418, -36.56922, -36.67581, 
    -36.77385, -36.86326, -36.94396, -37.01588, -37.07895, -37.13312, 
    -37.17834, -37.21456, -37.24176, -37.2599, -37.26898, -37.26898, 
    -37.2599, -37.24176, -37.21456, -37.17834, -37.13312, -37.07895, 
    -37.01588, -36.94396, -36.86326, -36.77385, -36.67581, -36.56922, 
    -36.45418, -36.33079, -36.19914, -36.05936, -35.91155, -35.75585, 
    -35.59236, -35.42123, -35.24258, -35.05656, -34.86331, -34.66297, 
    -34.45568, -34.2416, -34.02087, -33.79364, -33.56009, -33.32034, 
    -33.07457, -32.82292, -32.56555, -32.30262, -32.03428, -31.76069, 
    -31.482, -31.19835, -30.90992, -30.61683, -30.31924, -30.0173, -29.71115, 
    -29.40093, -29.08677, -28.76883, -28.44723,
  -27.70978, -28.02592, -28.33856, -28.64755, -28.95277, -29.25407, 
    -29.55131, -29.84434, -30.13302, -30.4172, -30.69673, -30.97146, 
    -31.24123, -31.50589, -31.76528, -32.01924, -32.26763, -32.51027, 
    -32.74702, -32.97771, -33.2022, -33.42032, -33.63192, -33.83684, 
    -34.03494, -34.22607, -34.41008, -34.58682, -34.75616, -34.91797, 
    -35.0721, -35.21843, -35.35684, -35.48721, -35.60942, -35.72337, 
    -35.82896, -35.9261, -36.01469, -36.09467, -36.16594, -36.22845, 
    -36.28214, -36.32696, -36.36287, -36.38982, -36.40781, -36.41681, 
    -36.41681, -36.40781, -36.38982, -36.36287, -36.32696, -36.28214, 
    -36.22845, -36.16594, -36.09467, -36.01469, -35.9261, -35.82896, 
    -35.72337, -35.60942, -35.48721, -35.35684, -35.21843, -35.0721, 
    -34.91797, -34.75616, -34.58682, -34.41008, -34.22607, -34.03494, 
    -33.83684, -33.63192, -33.42032, -33.2022, -32.97771, -32.74702, 
    -32.51027, -32.26763, -32.01924, -31.76528, -31.50589, -31.24123, 
    -30.97146, -30.69673, -30.4172, -30.13302, -29.84434, -29.55131, 
    -29.25407, -28.95277, -28.64755, -28.33856, -28.02592, -27.70978,
  -26.97222, -27.28269, -27.58981, -27.89343, -28.19342, -28.48965, 
    -28.78197, -29.07022, -29.35428, -29.63398, -29.90917, -30.17971, 
    -30.44544, -30.7062, -30.96183, -31.21218, -31.45709, -31.6964, 
    -31.92994, -32.15757, -32.37912, -32.59444, -32.80336, -33.00574, 
    -33.20141, -33.39024, -33.57207, -33.74675, -33.91414, -34.07411, 
    -34.22652, -34.37123, -34.50814, -34.6371, -34.75802, -34.87078, 
    -34.97528, -35.07141, -35.15911, -35.23827, -35.30883, -35.37072, 
    -35.42388, -35.46826, -35.50381, -35.53051, -35.54832, -35.55723, 
    -35.55723, -35.54832, -35.53051, -35.50381, -35.46826, -35.42388, 
    -35.37072, -35.30883, -35.23827, -35.15911, -35.07141, -34.97528, 
    -34.87078, -34.75802, -34.6371, -34.50814, -34.37123, -34.22652, 
    -34.07411, -33.91414, -33.74675, -33.57207, -33.39024, -33.20141, 
    -33.00574, -32.80336, -32.59444, -32.37912, -32.15757, -31.92994, 
    -31.6964, -31.45709, -31.21218, -30.96183, -30.7062, -30.44544, 
    -30.17971, -29.90917, -29.63398, -29.35428, -29.07022, -28.78197, 
    -28.48965, -28.19342, -27.89343, -27.58981, -27.28269, -26.97222,
  -26.23456, -26.53915, -26.84053, -27.13857, -27.43312, -27.72406, 
    -28.01123, -28.29449, -28.5737, -28.84871, -29.11935, -29.38548, 
    -29.64695, -29.90359, -30.15525, -30.40177, -30.643, -30.87876, 
    -31.10889, -31.33325, -31.55167, -31.76398, -31.97004, -32.16968, 
    -32.36275, -32.5491, -32.72858, -32.90103, -33.06631, -33.2243, 
    -33.37484, -33.5178, -33.65307, -33.78051, -33.90001, -34.01146, 
    -34.11476, -34.20981, -34.29651, -34.37479, -34.44456, -34.50577, 
    -34.55835, -34.60224, -34.63741, -34.66381, -34.68143, -34.69025, 
    -34.69025, -34.68143, -34.66381, -34.63741, -34.60224, -34.55835, 
    -34.50577, -34.44456, -34.37479, -34.29651, -34.20981, -34.11476, 
    -34.01146, -33.90001, -33.78051, -33.65307, -33.5178, -33.37484, 
    -33.2243, -33.06631, -32.90103, -32.72858, -32.5491, -32.36275, 
    -32.16968, -31.97004, -31.76398, -31.55167, -31.33325, -31.10889, 
    -30.87876, -30.643, -30.40177, -30.15525, -29.90359, -29.64695, 
    -29.38548, -29.11935, -28.84871, -28.5737, -28.29449, -28.01123, 
    -27.72406, -27.43312, -27.13857, -26.84053, -26.53915, -26.23456,
  -25.4968, -25.7953, -26.09074, -26.38298, -26.67189, -26.95732, -27.23913, 
    -27.51719, -27.79133, -28.06141, -28.32729, -28.5888, -28.84579, 
    -29.0981, -29.34557, -29.58805, -29.82537, -30.05738, -30.28391, 
    -30.50479, -30.71988, -30.929, -31.132, -31.32872, -31.519, -31.70269, 
    -31.87964, -32.0497, -32.21272, -32.36856, -32.51709, -32.65816, 
    -32.79165, -32.91744, -33.03541, -33.14545, -33.24744, -33.3413, 
    -33.42693, -33.50424, -33.57316, -33.63363, -33.68556, -33.72892, 
    -33.76367, -33.78976, -33.80717, -33.81588, -33.81588, -33.80717, 
    -33.78976, -33.76367, -33.72892, -33.68556, -33.63363, -33.57316, 
    -33.50424, -33.42693, -33.3413, -33.24744, -33.14545, -33.03541, 
    -32.91744, -32.79165, -32.65816, -32.51709, -32.36856, -32.21272, 
    -32.0497, -31.87964, -31.70269, -31.519, -31.32872, -31.132, -30.929, 
    -30.71988, -30.50479, -30.28391, -30.05738, -29.82537, -29.58805, 
    -29.34557, -29.0981, -28.84579, -28.5888, -28.32729, -28.06141, 
    -27.79133, -27.51719, -27.23913, -26.95732, -26.67189, -26.38298, 
    -26.09074, -25.7953, -25.4968,
  -24.75893, -25.05115, -25.34044, -25.62668, -25.90973, -26.18944, 
    -26.46569, -26.73832, -27.00718, -27.27213, -27.53302, -27.78969, 
    -28.04199, -28.28975, -28.53283, -28.77106, -29.00427, -29.23232, 
    -29.45502, -29.67224, -29.88379, -30.08952, -30.28927, -30.48288, 
    -30.6702, -30.85106, -31.02531, -31.19281, -31.3534, -31.50695, 
    -31.65331, -31.79235, -31.92393, -32.04794, -32.16426, -32.27277, 
    -32.37335, -32.46593, -32.55039, -32.62666, -32.69466, -32.75431, 
    -32.80555, -32.84834, -32.88263, -32.90837, -32.92555, -32.93415, 
    -32.93415, -32.92555, -32.90837, -32.88263, -32.84834, -32.80555, 
    -32.75431, -32.69466, -32.62666, -32.55039, -32.46593, -32.37335, 
    -32.27277, -32.16426, -32.04794, -31.92393, -31.79235, -31.65331, 
    -31.50695, -31.3534, -31.19281, -31.02531, -30.85106, -30.6702, 
    -30.48288, -30.28927, -30.08952, -29.88379, -29.67224, -29.45502, 
    -29.23232, -29.00427, -28.77106, -28.53283, -28.28975, -28.04199, 
    -27.78969, -27.53302, -27.27213, -27.00718, -26.73832, -26.46569, 
    -26.18944, -25.90973, -25.62668, -25.34044, -25.05115, -24.75893,
  -24.02097, -24.3067, -24.58965, -24.86968, -25.14667, -25.42046, -25.69092, 
    -25.95792, -26.22129, -26.4809, -26.73659, -26.98821, -27.2356, 
    -27.47861, -27.71707, -27.95084, -28.17974, -28.40361, -28.6223, 
    -28.83563, -29.04346, -29.2456, -29.44192, -29.63223, -29.81639, 
    -29.99424, -30.16563, -30.3304, -30.4884, -30.6395, -30.78355, -30.92041, 
    -31.04995, -31.17205, -31.28659, -31.39346, -31.49253, -31.58372, 
    -31.66694, -31.74208, -31.80908, -31.86786, -31.91836, -31.96053, 
    -31.99432, -32.01969, -32.03662, -32.04509, -32.04509, -32.03662, 
    -32.01969, -31.99432, -31.96053, -31.91836, -31.86786, -31.80908, 
    -31.74208, -31.66694, -31.58372, -31.49253, -31.39346, -31.28659, 
    -31.17205, -31.04995, -30.92041, -30.78355, -30.6395, -30.4884, -30.3304, 
    -30.16563, -29.99424, -29.81639, -29.63223, -29.44192, -29.2456, 
    -29.04346, -28.83563, -28.6223, -28.40361, -28.17974, -27.95084, 
    -27.71707, -27.47861, -27.2356, -26.98821, -26.73659, -26.4809, 
    -26.22129, -25.95792, -25.69092, -25.42046, -25.14667, -24.86968, 
    -24.58965, -24.3067, -24.02097,
  -23.28291, -23.56197, -23.83837, -24.112, -24.38272, -24.65038, -24.91487, 
    -25.17602, -25.43369, -25.68774, -25.93803, -26.18438, -26.42666, 
    -26.6647, -26.89834, -27.12744, -27.35181, -27.57131, -27.78577, 
    -27.99503, -28.19893, -28.3973, -28.58998, -28.77681, -28.95764, 
    -29.1323, -29.30065, -29.46252, -29.61777, -29.76627, -29.90785, 
    -30.04239, -30.16976, -30.28983, -30.40247, -30.50758, -30.60504, 
    -30.69475, -30.77662, -30.85055, -30.91648, -30.97433, -31.02403, 
    -31.06553, -31.09879, -31.12376, -31.14043, -31.14876, -31.14876, 
    -31.14043, -31.12376, -31.09879, -31.06553, -31.02403, -30.97433, 
    -30.91648, -30.85055, -30.77662, -30.69475, -30.60504, -30.50758, 
    -30.40247, -30.28983, -30.16976, -30.04239, -29.90785, -29.76627, 
    -29.61777, -29.46252, -29.30065, -29.1323, -28.95764, -28.77681, 
    -28.58998, -28.3973, -28.19893, -27.99503, -27.78577, -27.57131, 
    -27.35181, -27.12744, -26.89834, -26.6647, -26.42666, -26.18438, 
    -25.93803, -25.68774, -25.43369, -25.17602, -24.91487, -24.65038, 
    -24.38272, -24.112, -23.83837, -23.56197, -23.28291,
  -22.54476, -22.81695, -23.08662, -23.35365, -23.6179, -23.87924, -24.13754, 
    -24.39264, -24.64441, -24.89271, -25.13737, -25.37826, -25.61521, 
    -25.84807, -26.07669, -26.30091, -26.52055, -26.73548, -26.94551, 
    -27.1505, -27.35027, -27.54466, -27.73353, -27.91669, -28.094, -28.2653, 
    -28.43043, -28.58924, -28.74158, -28.88731, -29.02629, -29.15837, 
    -29.28342, -29.40132, -29.51195, -29.61518, -29.71092, -29.79905, 
    -29.87949, -29.95214, -30.01692, -30.07377, -30.12261, -30.1634, 
    -30.19609, -30.22064, -30.23702, -30.24521, -30.24521, -30.23702, 
    -30.22064, -30.19609, -30.1634, -30.12261, -30.07377, -30.01692, 
    -29.95214, -29.87949, -29.79905, -29.71092, -29.61518, -29.51195, 
    -29.40132, -29.28342, -29.15837, -29.02629, -28.88731, -28.74158, 
    -28.58924, -28.43043, -28.2653, -28.094, -27.91669, -27.73353, -27.54466, 
    -27.35027, -27.1505, -26.94551, -26.73548, -26.52055, -26.30091, 
    -26.07669, -25.84807, -25.61521, -25.37826, -25.13737, -24.89271, 
    -24.64441, -24.39264, -24.13754, -23.87924, -23.6179, -23.35365, 
    -23.08662, -22.81695, -22.54476,
  -21.80651, -22.07165, -22.33441, -22.59464, -22.85224, -23.10706, 
    -23.35897, -23.60783, -23.85349, -24.09582, -24.33467, -24.56988, 
    -24.8013, -25.02878, -25.25217, -25.4713, -25.68602, -25.89616, 
    -26.10157, -26.30208, -26.49753, -26.68777, -26.87262, -27.05193, 
    -27.22555, -27.3933, -27.55505, -27.71063, -27.8599, -28.00271, 
    -28.13892, -28.2684, -28.391, -28.50661, -28.6151, -28.71634, -28.81025, 
    -28.89671, -28.97562, -29.0469, -29.11047, -29.16625, -29.21418, 
    -29.25421, -29.28629, -29.31038, -29.32646, -29.33451, -29.33451, 
    -29.32646, -29.31038, -29.28629, -29.25421, -29.21418, -29.16625, 
    -29.11047, -29.0469, -28.97562, -28.89671, -28.81025, -28.71634, 
    -28.6151, -28.50661, -28.391, -28.2684, -28.13892, -28.00271, -27.8599, 
    -27.71063, -27.55505, -27.3933, -27.22555, -27.05193, -26.87262, 
    -26.68777, -26.49753, -26.30208, -26.10157, -25.89616, -25.68602, 
    -25.4713, -25.25217, -25.02878, -24.8013, -24.56988, -24.33467, 
    -24.09582, -23.85349, -23.60783, -23.35897, -23.10706, -22.85224, 
    -22.59464, -22.33441, -22.07165, -21.80651,
  -21.06818, -21.32609, -21.58174, -21.835, -22.08575, -22.33386, -22.57919, 
    -22.8216, -23.06096, -23.29713, -23.52995, -23.75929, -23.98498, 
    -24.20688, -24.42483, -24.63868, -24.84826, -25.05343, -25.25401, 
    -25.44986, -25.6408, -25.82668, -26.00734, -26.18261, -26.35234, 
    -26.51638, -26.67457, -26.82676, -26.9728, -27.11254, -27.24584, 
    -27.37256, -27.49258, -27.60576, -27.71199, -27.81114, -27.90311, 
    -27.98779, -28.06509, -28.13491, -28.19719, -28.25185, -28.29881, 
    -28.33804, -28.36947, -28.39308, -28.40884, -28.41672, -28.41672, 
    -28.40884, -28.39308, -28.36947, -28.33804, -28.29881, -28.25185, 
    -28.19719, -28.13491, -28.06509, -27.98779, -27.90311, -27.81114, 
    -27.71199, -27.60576, -27.49258, -27.37256, -27.24584, -27.11254, 
    -26.9728, -26.82676, -26.67457, -26.51638, -26.35234, -26.18261, 
    -26.00734, -25.82668, -25.6408, -25.44986, -25.25401, -25.05343, 
    -24.84826, -24.63868, -24.42483, -24.20688, -23.98498, -23.75929, 
    -23.52995, -23.29713, -23.06096, -22.8216, -22.57919, -22.33386, 
    -22.08575, -21.835, -21.58174, -21.32609, -21.06818,
  -20.32976, -20.58027, -20.82863, -21.07474, -21.31846, -21.55966, 
    -21.79822, -22.034, -22.26687, -22.49667, -22.72328, -22.94654, -23.1663, 
    -23.38242, -23.59474, -23.8031, -24.00736, -24.20735, -24.40292, 
    -24.5939, -24.78014, -24.96147, -25.13775, -25.3088, -25.47448, 
    -25.63463, -25.78909, -25.93772, -26.08036, -26.21687, -26.34712, 
    -26.47095, -26.58825, -26.69888, -26.80272, -26.89966, -26.98958, 
    -27.07239, -27.14798, -27.21628, -27.27719, -27.33065, -27.3766, 
    -27.41497, -27.44572, -27.46882, -27.48424, -27.49195, -27.49195, 
    -27.48424, -27.46882, -27.44572, -27.41497, -27.3766, -27.33065, 
    -27.27719, -27.21628, -27.14798, -27.07239, -26.98958, -26.89966, 
    -26.80272, -26.69888, -26.58825, -26.47095, -26.34712, -26.21687, 
    -26.08036, -25.93772, -25.78909, -25.63463, -25.47448, -25.3088, 
    -25.13775, -24.96147, -24.78014, -24.5939, -24.40292, -24.20735, 
    -24.00736, -23.8031, -23.59474, -23.38242, -23.1663, -22.94654, 
    -22.72328, -22.49667, -22.26687, -22.034, -21.79822, -21.55966, 
    -21.31846, -21.07474, -20.82863, -20.58027, -20.32976,
  -19.59126, -19.83419, -20.0751, -20.31387, -20.55038, -20.7845, -21.01611, 
    -21.24507, -21.47124, -21.6945, -21.91469, -22.13168, -22.34532, 
    -22.55546, -22.76195, -22.96464, -23.16337, -23.35799, -23.54835, 
    -23.73428, -23.91562, -24.09223, -24.26394, -24.43059, -24.59204, 
    -24.74813, -24.89869, -25.04359, -25.18268, -25.31582, -25.44285, 
    -25.56366, -25.6781, -25.78605, -25.88738, -25.98199, -26.06977, 
    -26.1506, -26.2244, -26.29108, -26.35056, -26.40276, -26.44763, -26.4851, 
    -26.51514, -26.5377, -26.55275, -26.56029, -26.56029, -26.55275, 
    -26.5377, -26.51514, -26.4851, -26.44763, -26.40276, -26.35056, 
    -26.29108, -26.2244, -26.1506, -26.06977, -25.98199, -25.88738, 
    -25.78605, -25.6781, -25.56366, -25.44285, -25.31582, -25.18268, 
    -25.04359, -24.89869, -24.74813, -24.59204, -24.43059, -24.26394, 
    -24.09223, -23.91562, -23.73428, -23.54835, -23.35799, -23.16337, 
    -22.96464, -22.76195, -22.55546, -22.34532, -22.13168, -21.91469, 
    -21.6945, -21.47124, -21.24507, -21.01611, -20.7845, -20.55038, 
    -20.31387, -20.0751, -19.83419, -19.59126,
  -18.85267, -19.08786, -19.32115, -19.55242, -19.78154, -20.0084, -20.23287, 
    -20.45482, -20.67413, -20.89065, -21.10424, -21.31477, -21.52209, 
    -21.72607, -21.92654, -22.12335, -22.31637, -22.50543, -22.69039, 
    -22.87107, -23.04734, -23.21904, -23.386, -23.54808, -23.70512, 
    -23.85697, -24.00347, -24.14449, -24.27987, -24.40947, -24.53315, 
    -24.65079, -24.76223, -24.86737, -24.96609, -25.05826, -25.14377, 
    -25.22254, -25.29446, -25.35944, -25.41741, -25.46829, -25.51202, 
    -25.54855, -25.57783, -25.59982, -25.6145, -25.62184, -25.62184, 
    -25.6145, -25.59982, -25.57783, -25.54855, -25.51202, -25.46829, 
    -25.41741, -25.35944, -25.29446, -25.22254, -25.14377, -25.05826, 
    -24.96609, -24.86737, -24.76223, -24.65079, -24.53315, -24.40947, 
    -24.27987, -24.14449, -24.00347, -23.85697, -23.70512, -23.54808, 
    -23.386, -23.21904, -23.04734, -22.87107, -22.69039, -22.50543, 
    -22.31637, -22.12335, -21.92654, -21.72607, -21.52209, -21.31477, 
    -21.10424, -20.89065, -20.67413, -20.45482, -20.23287, -20.0084, 
    -19.78154, -19.55242, -19.32115, -19.08786, -18.85267,
  -18.114, -18.3413, -18.5668, -18.79039, -19.01196, -19.23139, -19.44855, 
    -19.66332, -19.87557, -20.08517, -20.29198, -20.49586, -20.69669, 
    -20.8943, -21.08856, -21.27932, -21.46644, -21.64975, -21.82912, 
    -22.00438, -22.17539, -22.34199, -22.50403, -22.66135, -22.81381, 
    -22.96125, -23.10353, -23.2405, -23.37202, -23.49794, -23.61813, 
    -23.73245, -23.84077, -23.94298, -24.03895, -24.12856, -24.21172, 
    -24.28832, -24.35827, -24.42147, -24.47786, -24.52736, -24.5699, 
    -24.60544, -24.63392, -24.65532, -24.6696, -24.67674, -24.67674, 
    -24.6696, -24.65532, -24.63392, -24.60544, -24.5699, -24.52736, 
    -24.47786, -24.42147, -24.35827, -24.28832, -24.21172, -24.12856, 
    -24.03895, -23.94298, -23.84077, -23.73245, -23.61813, -23.49794, 
    -23.37202, -23.2405, -23.10353, -22.96125, -22.81381, -22.66135, 
    -22.50403, -22.34199, -22.17539, -22.00438, -21.82912, -21.64975, 
    -21.46644, -21.27932, -21.08856, -20.8943, -20.69669, -20.49586, 
    -20.29198, -20.08517, -19.87557, -19.66332, -19.44855, -19.23139, 
    -19.01196, -18.79039, -18.5668, -18.3413, -18.114,
  -17.37526, -17.59451, -17.81206, -18.02782, -18.24167, -18.45349, 
    -18.66317, -18.87058, -19.07561, -19.2781, -19.47795, -19.67501, 
    -19.86915, -20.06023, -20.2481, -20.43262, -20.61365, -20.79103, 
    -20.96463, -21.13428, -21.29985, -21.46118, -21.61812, -21.77052, 
    -21.91823, -22.0611, -22.19899, -22.33176, -22.45926, -22.58134, 
    -22.69789, -22.80877, -22.91384, -23.01299, -23.10609, -23.19304, 
    -23.27374, -23.34808, -23.41596, -23.47731, -23.53204, -23.58009, 
    -23.62139, -23.6559, -23.68355, -23.70432, -23.71819, -23.72513, 
    -23.72513, -23.71819, -23.70432, -23.68355, -23.6559, -23.62139, 
    -23.58009, -23.53204, -23.47731, -23.41596, -23.34808, -23.27374, 
    -23.19304, -23.10609, -23.01299, -22.91384, -22.80877, -22.69789, 
    -22.58134, -22.45926, -22.33176, -22.19899, -22.0611, -21.91823, 
    -21.77052, -21.61812, -21.46118, -21.29985, -21.13428, -20.96463, 
    -20.79103, -20.61365, -20.43262, -20.2481, -20.06023, -19.86915, 
    -19.67501, -19.47795, -19.2781, -19.07561, -18.87058, -18.66317, 
    -18.45349, -18.24167, -18.02782, -17.81206, -17.59451, -17.37526,
  -16.63645, -16.84749, -17.05695, -17.26471, -17.47068, -17.67474, 
    -17.87678, -18.07666, -18.27429, -18.46952, -18.66223, -18.85229, 
    -19.03956, -19.22392, -19.40522, -19.58332, -19.75808, -19.92936, 
    -20.09701, -20.26088, -20.42083, -20.57672, -20.72838, -20.87569, 
    -21.01848, -21.15662, -21.28997, -21.41838, -21.5417, -21.65982, 
    -21.77258, -21.87987, -21.98156, -22.07753, -22.16766, -22.25184, 
    -22.32997, -22.40195, -22.46768, -22.52709, -22.5801, -22.62664, 
    -22.66665, -22.70007, -22.72686, -22.74698, -22.76041, -22.76713, 
    -22.76713, -22.76041, -22.74698, -22.72686, -22.70007, -22.66665, 
    -22.62664, -22.5801, -22.52709, -22.46768, -22.40195, -22.32997, 
    -22.25184, -22.16766, -22.07753, -21.98156, -21.87987, -21.77258, 
    -21.65982, -21.5417, -21.41838, -21.28997, -21.15662, -21.01848, 
    -20.87569, -20.72838, -20.57672, -20.42083, -20.26088, -20.09701, 
    -19.92936, -19.75808, -19.58332, -19.40522, -19.22392, -19.03956, 
    -18.85229, -18.66223, -18.46952, -18.27429, -18.07666, -17.87678, 
    -17.67474, -17.47068, -17.26471, -17.05695, -16.84749, -16.63645,
  -15.89756, -16.10026, -16.30147, -16.50109, -16.69903, -16.89517, -17.0894, 
    -17.2816, -17.47165, -17.65945, -17.84485, -18.02774, -18.20799, 
    -18.38545, -18.56001, -18.73152, -18.89984, -19.06483, -19.22636, 
    -19.38427, -19.53844, -19.68871, -19.83493, -19.97698, -20.11469, 
    -20.24794, -20.37659, -20.50048, -20.61949, -20.73348, -20.84233, 
    -20.94591, -21.04409, -21.13675, -21.22379, -21.30509, -21.38055, 
    -21.45008, -21.51358, -21.57098, -21.6222, -21.66716, -21.70582, 
    -21.73811, -21.764, -21.78345, -21.79643, -21.80292, -21.80292, 
    -21.79643, -21.78345, -21.764, -21.73811, -21.70582, -21.66716, -21.6222, 
    -21.57098, -21.51358, -21.45008, -21.38055, -21.30509, -21.22379, 
    -21.13675, -21.04409, -20.94591, -20.84233, -20.73348, -20.61949, 
    -20.50048, -20.37659, -20.24794, -20.11469, -19.97698, -19.83493, 
    -19.68871, -19.53844, -19.38427, -19.22636, -19.06483, -18.89984, 
    -18.73152, -18.56001, -18.38545, -18.20799, -18.02774, -17.84485, 
    -17.65945, -17.47165, -17.2816, -17.0894, -16.89517, -16.69903, 
    -16.50109, -16.30147, -16.10026, -15.89756,
  -15.15861, -15.35282, -15.54564, -15.73699, -15.92674, -16.11481, 
    -16.30107, -16.48543, -16.66776, -16.84796, -17.02589, -17.20144, 
    -17.37449, -17.5449, -17.71254, -17.87728, -18.03899, -18.19754, 
    -18.35277, -18.50457, -18.65277, -18.79726, -18.93789, -19.07451, 
    -19.20699, -19.33519, -19.45897, -19.57821, -19.69276, -19.8025, 
    -19.90729, -20.00702, -20.10156, -20.19081, -20.27464, -20.35295, 
    -20.42565, -20.49264, -20.55383, -20.60913, -20.65849, -20.70182, 
    -20.73908, -20.7702, -20.79515, -20.81389, -20.8264, -20.83266, 
    -20.83266, -20.8264, -20.81389, -20.79515, -20.7702, -20.73908, 
    -20.70182, -20.65849, -20.60913, -20.55383, -20.49264, -20.42565, 
    -20.35295, -20.27464, -20.19081, -20.10156, -20.00702, -19.90729, 
    -19.8025, -19.69276, -19.57821, -19.45897, -19.33519, -19.20699, 
    -19.07451, -18.93789, -18.79726, -18.65277, -18.50457, -18.35277, 
    -18.19754, -18.03899, -17.87728, -17.71254, -17.5449, -17.37449, 
    -17.20144, -17.02589, -16.84796, -16.66776, -16.48543, -16.30107, 
    -16.11481, -15.92674, -15.73699, -15.54564, -15.35282, -15.15861,
  -14.41959, -14.60518, -14.78949, -14.9724, -15.15383, -15.33368, -15.51184, 
    -15.6882, -15.86266, -16.0351, -16.20541, -16.37346, -16.53915, 
    -16.70233, -16.8629, -17.02072, -17.17565, -17.32758, -17.47636, 
    -17.62187, -17.76396, -17.9025, -18.03736, -18.16841, -18.2955, -18.4185, 
    -18.53728, -18.65171, -18.76166, -18.867, -18.96761, -19.06337, 
    -19.15416, -19.23986, -19.32038, -19.39561, -19.46544, -19.5298, 
    -19.58859, -19.64173, -19.68916, -19.7308, -19.7666, -19.79651, 
    -19.82049, -19.8385, -19.85053, -19.85655, -19.85655, -19.85053, 
    -19.8385, -19.82049, -19.79651, -19.7666, -19.7308, -19.68916, -19.64173, 
    -19.58859, -19.5298, -19.46544, -19.39561, -19.32038, -19.23986, 
    -19.15416, -19.06337, -18.96761, -18.867, -18.76166, -18.65171, 
    -18.53728, -18.4185, -18.2955, -18.16841, -18.03736, -17.9025, -17.76396, 
    -17.62187, -17.47636, -17.32758, -17.17565, -17.02072, -16.8629, 
    -16.70233, -16.53915, -16.37346, -16.20541, -16.0351, -15.86266, 
    -15.6882, -15.51184, -15.33368, -15.15383, -14.9724, -14.78949, 
    -14.60518, -14.41959,
  -13.6805, -13.85736, -14.03301, -14.20737, -14.38034, -14.55183, -14.72173, 
    -14.88996, -15.05639, -15.22093, -15.38346, -15.54386, -15.70203, 
    -15.85784, -16.01117, -16.1619, -16.30991, -16.45506, -16.59723, 
    -16.73629, -16.87211, -17.00456, -17.1335, -17.25882, -17.38036, 
    -17.49802, -17.61165, -17.72114, -17.82635, -17.92716, -18.02345, 
    -18.11512, -18.20203, -18.28409, -18.36119, -18.43323, -18.50011, 
    -18.56174, -18.61805, -18.66896, -18.71439, -18.75428, -18.78858, 
    -18.81724, -18.84021, -18.85747, -18.86899, -18.87476, -18.87476, 
    -18.86899, -18.85747, -18.84021, -18.81724, -18.78858, -18.75428, 
    -18.71439, -18.66896, -18.61805, -18.56174, -18.50011, -18.43323, 
    -18.36119, -18.28409, -18.20203, -18.11512, -18.02345, -17.92716, 
    -17.82635, -17.72114, -17.61165, -17.49802, -17.38036, -17.25882, 
    -17.1335, -17.00456, -16.87211, -16.73629, -16.59723, -16.45506, 
    -16.30991, -16.1619, -16.01117, -15.85784, -15.70203, -15.54386, 
    -15.38346, -15.22093, -15.05639, -14.88996, -14.72173, -14.55183, 
    -14.38034, -14.20737, -14.03301, -13.85736, -13.6805,
  -12.94136, -13.10935, -13.27623, -13.4419, -13.60628, -13.76928, -13.9308, 
    -14.09074, -14.24901, -14.4055, -14.56011, -14.71272, -14.86322, 
    -15.0115, -15.15745, -15.30094, -15.44186, -15.58009, -15.71549, 
    -15.84795, -15.97735, -16.10355, -16.22643, -16.34587, -16.46173, 
    -16.57389, -16.68224, -16.78664, -16.88698, -16.98314, -17.075, 
    -17.16244, -17.24537, -17.32367, -17.39725, -17.466, -17.52983, 
    -17.58866, -17.64242, -17.69101, -17.73438, -17.77247, -17.80522, 
    -17.83258, -17.85452, -17.871, -17.882, -17.88751, -17.88751, -17.882, 
    -17.871, -17.85452, -17.83258, -17.80522, -17.77247, -17.73438, 
    -17.69101, -17.64242, -17.58866, -17.52983, -17.466, -17.39725, 
    -17.32367, -17.24537, -17.16244, -17.075, -16.98314, -16.88698, 
    -16.78664, -16.68224, -16.57389, -16.46173, -16.34587, -16.22643, 
    -16.10355, -15.97735, -15.84795, -15.71549, -15.58009, -15.44186, 
    -15.30094, -15.15745, -15.0115, -14.86322, -14.71272, -14.56011, 
    -14.4055, -14.24901, -14.09074, -13.9308, -13.76928, -13.60628, -13.4419, 
    -13.27623, -13.10935, -12.94136,
  -12.20216, -12.36118, -12.51916, -12.67602, -12.83169, -12.98607, 
    -13.13908, -13.29061, -13.44058, -13.58888, -13.73542, -13.88009, 
    -14.02279, -14.1634, -14.30182, -14.43793, -14.57162, -14.70277, 
    -14.83126, -14.95698, -15.07981, -15.19962, -15.31629, -15.42971, 
    -15.53974, -15.64629, -15.74921, -15.8484, -15.94374, -16.03511, 
    -16.12242, -16.20553, -16.28436, -16.3588, -16.42875, -16.49412, 
    -16.55482, -16.61077, -16.66188, -16.7081, -16.74936, -16.78558, 
    -16.81673, -16.84276, -16.86363, -16.87931, -16.88978, -16.89501, 
    -16.89501, -16.88978, -16.87931, -16.86363, -16.84276, -16.81673, 
    -16.78558, -16.74936, -16.7081, -16.66188, -16.61077, -16.55482, 
    -16.49412, -16.42875, -16.3588, -16.28436, -16.20553, -16.12242, 
    -16.03511, -15.94374, -15.8484, -15.74921, -15.64629, -15.53974, 
    -15.42971, -15.31629, -15.19962, -15.07981, -14.95698, -14.83126, 
    -14.70277, -14.57162, -14.43793, -14.30182, -14.1634, -14.02279, 
    -13.88009, -13.73542, -13.58888, -13.44058, -13.29061, -13.13908, 
    -12.98607, -12.83169, -12.67602, -12.51916, -12.36118, -12.20216,
  -11.46291, -11.61284, -11.76182, -11.90976, -12.05659, -12.20224, -12.3466, 
    -12.4896, -12.63114, -12.77113, -12.90947, -13.04607, -13.18083, 
    -13.31363, -13.44438, -13.57297, -13.69929, -13.82323, -13.94467, 
    -14.0635, -14.17962, -14.2929, -14.40323, -14.51049, -14.61457, 
    -14.71535, -14.81272, -14.90658, -14.99679, -15.08327, -15.1659, 
    -15.24457, -15.3192, -15.38967, -15.4559, -15.5178, -15.57528, -15.62826, 
    -15.67667, -15.72045, -15.75952, -15.79384, -15.82335, -15.84801, 
    -15.86777, -15.88263, -15.89254, -15.8975, -15.8975, -15.89254, 
    -15.88263, -15.86777, -15.84801, -15.82335, -15.79384, -15.75952, 
    -15.72045, -15.67667, -15.62826, -15.57528, -15.5178, -15.4559, 
    -15.38967, -15.3192, -15.24457, -15.1659, -15.08327, -14.99679, 
    -14.90658, -14.81272, -14.71535, -14.61457, -14.51049, -14.40323, 
    -14.2929, -14.17962, -14.0635, -13.94467, -13.82323, -13.69929, 
    -13.57297, -13.44438, -13.31363, -13.18083, -13.04607, -12.90947, 
    -12.77113, -12.63114, -12.4896, -12.3466, -12.20224, -12.05659, 
    -11.90976, -11.76182, -11.61284, -11.46291,
  -10.72361, -10.86435, -11.00421, -11.14313, -11.28102, -11.41781, 
    -11.55342, -11.68776, -11.82075, -11.9523, -12.08233, -12.21073, 
    -12.33741, -12.46228, -12.58523, -12.70616, -12.82498, -12.94157, 
    -13.05583, -13.16765, -13.27692, -13.38354, -13.48739, -13.58837, 
    -13.68636, -13.78126, -13.87296, -13.96135, -14.04633, -14.1278, 
    -14.20564, -14.27977, -14.35008, -14.4165, -14.47891, -14.53725, 
    -14.59143, -14.64138, -14.68701, -14.72828, -14.76512, -14.79747, 
    -14.8253, -14.84855, -14.86719, -14.88119, -14.89054, -14.89522, 
    -14.89522, -14.89054, -14.88119, -14.86719, -14.84855, -14.8253, 
    -14.79747, -14.76512, -14.72828, -14.68701, -14.64138, -14.59143, 
    -14.53725, -14.47891, -14.4165, -14.35008, -14.27977, -14.20564, 
    -14.1278, -14.04633, -13.96135, -13.87296, -13.78126, -13.68636, 
    -13.58837, -13.48739, -13.38354, -13.27692, -13.16765, -13.05583, 
    -12.94157, -12.82498, -12.70616, -12.58523, -12.46228, -12.33741, 
    -12.21073, -12.08233, -11.9523, -11.82075, -11.68776, -11.55342, 
    -11.41781, -11.28102, -11.14313, -11.00421, -10.86435, -10.72361,
  -9.984256, -10.11571, -10.24637, -10.37615, -10.505, -10.63283, -10.75957, 
    -10.88514, -11.00947, -11.13247, -11.25405, -11.37413, -11.49262, 
    -11.60943, -11.72446, -11.83762, -11.9488, -12.05792, -12.16487, 
    -12.26954, -12.37185, -12.47168, -12.56893, -12.66351, -12.75529, 
    -12.84419, -12.9301, -13.01292, -13.09255, -13.16889, -13.24185, 
    -13.31133, -13.37724, -13.43949, -13.49801, -13.55271, -13.60351, 
    -13.65034, -13.69314, -13.73184, -13.76639, -13.79673, -13.82283, 
    -13.84463, -13.86212, -13.87526, -13.88403, -13.88841, -13.88841, 
    -13.88403, -13.87526, -13.86212, -13.84463, -13.82283, -13.79673, 
    -13.76639, -13.73184, -13.69314, -13.65034, -13.60351, -13.55271, 
    -13.49801, -13.43949, -13.37724, -13.31133, -13.24185, -13.16889, 
    -13.09255, -13.01292, -12.9301, -12.84419, -12.75529, -12.66351, 
    -12.56893, -12.47168, -12.37185, -12.26954, -12.16487, -12.05792, 
    -11.9488, -11.83762, -11.72446, -11.60943, -11.49262, -11.37413, 
    -11.25405, -11.13247, -11.00947, -10.88514, -10.75957, -10.63283, 
    -10.505, -10.37615, -10.24637, -10.11571, -9.984256,
  -9.244861, -9.366945, -9.488298, -9.608856, -9.728554, -9.847324, 
    -9.965097, -10.0818, -10.19736, -10.31169, -10.42472, -10.53637, 
    -10.64656, -10.75519, -10.86218, -10.96744, -11.07087, -11.1724, 
    -11.27192, -11.36934, -11.46456, -11.55748, -11.64802, -11.73607, 
    -11.82154, -11.90432, -11.98433, -12.06147, -12.13564, -12.20676, 
    -12.27472, -12.33946, -12.40088, -12.45889, -12.51342, -12.5644, 
    -12.61175, -12.6554, -12.6953, -12.73137, -12.76358, -12.79187, -12.8162, 
    -12.83653, -12.85283, -12.86508, -12.87325, -12.87735, -12.87735, 
    -12.87325, -12.86508, -12.85283, -12.83653, -12.8162, -12.79187, 
    -12.76358, -12.73137, -12.6953, -12.6554, -12.61175, -12.5644, -12.51342, 
    -12.45889, -12.40088, -12.33946, -12.27472, -12.20676, -12.13564, 
    -12.06147, -11.98433, -11.90432, -11.82154, -11.73607, -11.64802, 
    -11.55748, -11.46456, -11.36934, -11.27192, -11.1724, -11.07087, 
    -10.96744, -10.86218, -10.75519, -10.64656, -10.53637, -10.42472, 
    -10.31169, -10.19736, -10.0818, -9.965097, -9.847324, -9.728554, 
    -9.608856, -9.488298, -9.366945, -9.244861,
  -8.505425, -8.618052, -8.730017, -8.84126, -8.951721, -9.061338, -9.170046, 
    -9.277779, -9.384465, -9.490034, -9.594414, -9.697527, -9.799295, 
    -9.899641, -9.998483, -10.09574, -10.19132, -10.28514, -10.37712, 
    -10.46716, -10.55519, -10.6411, -10.72481, -10.80623, -10.88527, 
    -10.96183, -11.03584, -11.10719, -11.17581, -11.2416, -11.30449, 
    -11.3644, -11.42123, -11.47492, -11.52539, -11.57257, -11.6164, 
    -11.65681, -11.69374, -11.72714, -11.75696, -11.78315, -11.80567, 
    -11.8245, -11.83959, -11.85093, -11.8585, -11.86229, -11.86229, -11.8585, 
    -11.85093, -11.83959, -11.8245, -11.80567, -11.78315, -11.75696, 
    -11.72714, -11.69374, -11.65681, -11.6164, -11.57257, -11.52539, 
    -11.47492, -11.42123, -11.3644, -11.30449, -11.2416, -11.17581, 
    -11.10719, -11.03584, -10.96183, -10.88527, -10.80623, -10.72481, 
    -10.6411, -10.55519, -10.46716, -10.37712, -10.28514, -10.19132, 
    -10.09574, -9.998483, -9.899641, -9.799295, -9.697527, -9.594414, 
    -9.490034, -9.384465, -9.277779, -9.170046, -9.061338, -8.951721, 
    -8.84126, -8.730017, -8.618052, -8.505425,
  -7.765951, -7.869044, -7.971541, -8.073387, -8.174527, -8.274905, -8.37446, 
    -8.473132, -8.570855, -8.667565, -8.763195, -8.857674, -8.95093, 
    -9.042892, -9.133484, -9.222629, -9.31025, -9.396269, -9.480604, 
    -9.563174, -9.643898, -9.722692, -9.799476, -9.874163, -9.946671, 
    -10.01692, -10.08482, -10.1503, -10.21327, -10.27365, -10.33138, 
    -10.38636, -10.43853, -10.48782, -10.53416, -10.57748, -10.61772, 
    -10.65482, -10.68873, -10.7194, -10.74679, -10.77084, -10.79152, 
    -10.80881, -10.82268, -10.83309, -10.84004, -10.84352, -10.84352, 
    -10.84004, -10.83309, -10.82268, -10.80881, -10.79152, -10.77084, 
    -10.74679, -10.7194, -10.68873, -10.65482, -10.61772, -10.57748, 
    -10.53416, -10.48782, -10.43853, -10.38636, -10.33138, -10.27365, 
    -10.21327, -10.1503, -10.08482, -10.01692, -9.946671, -9.874163, 
    -9.799476, -9.722692, -9.643898, -9.563174, -9.480604, -9.396269, 
    -9.31025, -9.222629, -9.133484, -9.042892, -8.95093, -8.857674, 
    -8.763195, -8.667565, -8.570855, -8.473132, -8.37446, -8.274905, 
    -8.174527, -8.073387, -7.971541, -7.869044, -7.765951,
  -7.026442, -7.119931, -7.212887, -7.305261, -7.397004, -7.488063, 
    -7.578384, -7.667912, -7.756588, -7.844352, -7.931143, -8.016898, 
    -8.101551, -8.185037, -8.267286, -8.34823, -8.427797, -8.505915, 
    -8.582511, -8.657512, -8.730841, -8.802423, -8.872184, -8.940046, 
    -9.005934, -9.069772, -9.131484, -9.190996, -9.248235, -9.303126, 
    -9.355601, -9.40559, -9.453025, -9.49784, -9.539974, -9.579368, 
    -9.615962, -9.649706, -9.680549, -9.708443, -9.733348, -9.755226, 
    -9.774042, -9.789767, -9.802377, -9.811852, -9.818177, -9.821342, 
    -9.821342, -9.818177, -9.811852, -9.802377, -9.789767, -9.774042, 
    -9.755226, -9.733348, -9.708443, -9.680549, -9.649706, -9.615962, 
    -9.579368, -9.539974, -9.49784, -9.453025, -9.40559, -9.355601, 
    -9.303126, -9.248235, -9.190996, -9.131484, -9.069772, -9.005934, 
    -8.940046, -8.872184, -8.802423, -8.730841, -8.657512, -8.582511, 
    -8.505915, -8.427797, -8.34823, -8.267286, -8.185037, -8.101551, 
    -8.016898, -7.931143, -7.844352, -7.756588, -7.667912, -7.578384, 
    -7.488063, -7.397004, -7.305261, -7.212887, -7.119931, -7.026442,
  -6.286901, -6.370722, -6.454072, -6.536906, -6.619181, -6.70085, -6.781863, 
    -6.862171, -6.941722, -7.020462, -7.098334, -7.175284, -7.251252, 
    -7.326178, -7.4, -7.472656, -7.544083, -7.614214, -7.682984, -7.750327, 
    -7.816175, -7.880459, -7.943112, -8.004064, -8.063247, -8.120593, 
    -8.176033, -8.229501, -8.280929, -8.330251, -8.377405, -8.422327, 
    -8.464956, -8.505234, -8.543103, -8.578511, -8.611405, -8.641738, 
    -8.669463, -8.69454, -8.716929, -8.736598, -8.753514, -8.767653, 
    -8.77899, -8.787509, -8.793196, -8.796041, -8.796041, -8.793196, 
    -8.787509, -8.77899, -8.767653, -8.753514, -8.736598, -8.716929, 
    -8.69454, -8.669463, -8.641738, -8.611405, -8.578511, -8.543103, 
    -8.505234, -8.464956, -8.422327, -8.377405, -8.330251, -8.280929, 
    -8.229501, -8.176033, -8.120593, -8.063247, -8.004064, -7.943112, 
    -7.880459, -7.816175, -7.750327, -7.682984, -7.614214, -7.544083, 
    -7.472656, -7.4, -7.326178, -7.251252, -7.175284, -7.098334, -7.020462, 
    -6.941722, -6.862171, -6.781863, -6.70085, -6.619181, -6.536906, 
    -6.454072, -6.370722, -6.286901,
  -5.547333, -5.621428, -5.695111, -5.768345, -5.84109, -5.913303, -5.984942, 
    -6.055964, -6.12632, -6.195964, -6.264847, -6.332918, -6.400125, 
    -6.466415, -6.531734, -6.596026, -6.659235, -6.721301, -6.782168, 
    -6.841775, -6.900063, -6.956971, -7.012438, -7.066403, -7.118805, 
    -7.169584, -7.218679, -7.266029, -7.311576, -7.355261, -7.397027, 
    -7.436818, -7.47458, -7.510261, -7.54381, -7.57518, -7.604323, -7.631198, 
    -7.655765, -7.677984, -7.697824, -7.715252, -7.730243, -7.742771, 
    -7.752818, -7.760367, -7.765407, -7.767929, -7.767929, -7.765407, 
    -7.760367, -7.752818, -7.742771, -7.730243, -7.715252, -7.697824, 
    -7.677984, -7.655765, -7.631198, -7.604323, -7.57518, -7.54381, 
    -7.510261, -7.47458, -7.436818, -7.397027, -7.355261, -7.311576, 
    -7.266029, -7.218679, -7.169584, -7.118805, -7.066403, -7.012438, 
    -6.956971, -6.900063, -6.841775, -6.782168, -6.721301, -6.659235, 
    -6.596026, -6.531734, -6.466415, -6.400125, -6.332918, -6.264847, 
    -6.195964, -6.12632, -6.055964, -5.984942, -5.913303, -5.84109, 
    -5.768345, -5.695111, -5.621428, -5.547333,
  -4.807739, -4.872057, -4.936023, -4.999602, -5.06276, -5.125462, -5.187668, 
    -5.249342, -5.310442, -5.370928, -5.430757, -5.489884, -5.548265, 
    -5.605854, -5.662601, -5.718461, -5.773382, -5.827315, -5.880208, 
    -5.93201, -5.982669, -6.032131, -6.080344, -6.127254, -6.172808, 
    -6.216953, -6.259636, -6.300805, -6.340407, -6.378393, -6.414712, 
    -6.449316, -6.482156, -6.513187, -6.542367, -6.56965, -6.594999, 
    -6.618376, -6.639744, -6.659072, -6.676331, -6.691492, -6.704533, 
    -6.715432, -6.724172, -6.73074, -6.735124, -6.737318, -6.737318, 
    -6.735124, -6.73074, -6.724172, -6.715432, -6.704533, -6.691492, 
    -6.676331, -6.659072, -6.639744, -6.618376, -6.594999, -6.56965, 
    -6.542367, -6.513187, -6.482156, -6.449316, -6.414712, -6.378393, 
    -6.340407, -6.300805, -6.259636, -6.216953, -6.172808, -6.127254, 
    -6.080344, -6.032131, -5.982669, -5.93201, -5.880208, -5.827315, 
    -5.773382, -5.718461, -5.662601, -5.605854, -5.548265, -5.489884, 
    -5.430757, -5.370928, -5.310442, -5.249342, -5.187668, -5.125462, 
    -5.06276, -4.999602, -4.936023, -4.872057, -4.807739,
  -4.068124, -4.122622, -4.176824, -4.230701, -4.284225, -4.337364, 
    -4.390087, -4.442361, -4.494153, -4.545426, -4.596145, -4.646272, 
    -4.695769, -4.744597, -4.792715, -4.840082, -4.886656, -4.932395, 
    -4.977254, -5.02119, -5.064158, -5.106114, -5.147013, -5.186808, 
    -5.225454, -5.262908, -5.299122, -5.334054, -5.367657, -5.399891, 
    -5.430711, -5.460076, -5.487947, -5.514283, -5.539048, -5.562205, 
    -5.58372, -5.603562, -5.6217, -5.638107, -5.652757, -5.665627, -5.676696, 
    -5.685948, -5.693368, -5.698944, -5.702665, -5.704528, -5.704528, 
    -5.702665, -5.698944, -5.693368, -5.685948, -5.676696, -5.665627, 
    -5.652757, -5.638107, -5.6217, -5.603562, -5.58372, -5.562205, -5.539048, 
    -5.514283, -5.487947, -5.460076, -5.430711, -5.399891, -5.367657, 
    -5.334054, -5.299122, -5.262908, -5.225454, -5.186808, -5.147013, 
    -5.106114, -5.064158, -5.02119, -4.977254, -4.932395, -4.886656, 
    -4.840082, -4.792715, -4.744597, -4.695769, -4.646272, -4.596145, 
    -4.545426, -4.494153, -4.442361, -4.390087, -4.337364, -4.284225, 
    -4.230701, -4.176824, -4.122622, -4.068124,
  -3.32849, -3.37313, -3.41753, -3.461666, -3.505514, -3.549049, -3.592245, 
    -3.635076, -3.677513, -3.719527, -3.761089, -3.802168, -3.842732, 
    -3.88275, -3.922188, -3.961012, -3.999188, -4.036681, -4.073455, 
    -4.109474, -4.144701, -4.179099, -4.212631, -4.245261, -4.27695, 
    -4.307662, -4.337358, -4.366004, -4.393563, -4.419998, -4.445276, 
    -4.46936, -4.49222, -4.513822, -4.534135, -4.55313, -4.570779, -4.587056, 
    -4.601935, -4.615394, -4.627412, -4.63797, -4.647052, -4.654643, 
    -4.660729, -4.665304, -4.668357, -4.669885, -4.669885, -4.668357, 
    -4.665304, -4.660729, -4.654643, -4.647052, -4.63797, -4.627412, 
    -4.615394, -4.601935, -4.587056, -4.570779, -4.55313, -4.534135, 
    -4.513822, -4.49222, -4.46936, -4.445276, -4.419998, -4.393563, 
    -4.366004, -4.337358, -4.307662, -4.27695, -4.245261, -4.212631, 
    -4.179099, -4.144701, -4.109474, -4.073455, -4.036681, -3.999188, 
    -3.961012, -3.922188, -3.88275, -3.842732, -3.802168, -3.761089, 
    -3.719527, -3.677513, -3.635076, -3.592245, -3.549049, -3.505514, 
    -3.461666, -3.41753, -3.37313, -3.32849,
  -2.588841, -2.623593, -2.658159, -2.692521, -2.72666, -2.760556, -2.79419, 
    -2.827541, -2.860586, -2.893303, -2.925669, -2.957661, -2.989253, 
    -3.02042, -3.051136, -3.081377, -3.111113, -3.140318, -3.168964, 
    -3.197022, -3.224465, -3.251263, -3.277388, -3.30281, -3.3275, -3.35143, 
    -3.374569, -3.39689, -3.418365, -3.438965, -3.458663, -3.477432, 
    -3.495247, -3.512082, -3.527913, -3.542717, -3.556473, -3.569159, 
    -3.580756, -3.591246, -3.600614, -3.608843, -3.615922, -3.621838, 
    -3.626583, -3.630148, -3.632529, -3.63372, -3.63372, -3.632529, 
    -3.630148, -3.626583, -3.621838, -3.615922, -3.608843, -3.600614, 
    -3.591246, -3.580756, -3.569159, -3.556473, -3.542717, -3.527913, 
    -3.512082, -3.495247, -3.477432, -3.458663, -3.438965, -3.418365, 
    -3.39689, -3.374569, -3.35143, -3.3275, -3.30281, -3.277388, -3.251263, 
    -3.224465, -3.197022, -3.168964, -3.140318, -3.111113, -3.081377, 
    -3.051136, -3.02042, -2.989253, -2.957661, -2.925669, -2.893303, 
    -2.860586, -2.827541, -2.79419, -2.760556, -2.72666, -2.692521, 
    -2.658159, -2.623593, -2.588841,
  -1.849181, -1.87402, -1.898728, -1.92329, -1.947694, -1.971925, -1.995969, 
    -2.019811, -2.043435, -2.066826, -2.089966, -2.112839, -2.135427, 
    -2.157712, -2.179676, -2.201299, -2.222563, -2.243447, -2.263932, 
    -2.283998, -2.303623, -2.322789, -2.341473, -2.359655, -2.377314, 
    -2.394429, -2.41098, -2.426945, -2.442306, -2.457041, -2.471131, 
    -2.484558, -2.497301, -2.509345, -2.52067, -2.53126, -2.541101, 
    -2.550177, -2.558473, -2.565979, -2.57268, -2.578568, -2.583632, 
    -2.587865, -2.59126, -2.593811, -2.595514, -2.596366, -2.596366, 
    -2.595514, -2.593811, -2.59126, -2.587865, -2.583632, -2.578568, 
    -2.57268, -2.565979, -2.558473, -2.550177, -2.541101, -2.53126, -2.52067, 
    -2.509345, -2.497301, -2.484558, -2.471131, -2.457041, -2.442306, 
    -2.426945, -2.41098, -2.394429, -2.377314, -2.359655, -2.341473, 
    -2.322789, -2.303623, -2.283998, -2.263932, -2.243447, -2.222563, 
    -2.201299, -2.179676, -2.157712, -2.135427, -2.112839, -2.089966, 
    -2.066826, -2.043435, -2.019811, -1.995969, -1.971925, -1.947694, 
    -1.92329, -1.898728, -1.87402, -1.849181,
  -1.109512, -1.124422, -1.139254, -1.153999, -1.168648, -1.183195, 
    -1.197629, -1.211942, -1.226125, -1.240168, -1.254061, -1.267794, 
    -1.281355, -1.294735, -1.307923, -1.320906, -1.333673, -1.346213, 
    -1.358514, -1.370563, -1.382348, -1.393856, -1.405076, -1.415995, 
    -1.4266, -1.436878, -1.446817, -1.456406, -1.46563, -1.47448, -1.482942, 
    -1.491006, -1.49866, -1.505893, -1.512695, -1.519056, -1.524966, 
    -1.530417, -1.535401, -1.539908, -1.543934, -1.54747, -1.550512, 
    -1.553055, -1.555094, -1.556626, -1.557649, -1.55816, -1.55816, 
    -1.557649, -1.556626, -1.555094, -1.553055, -1.550512, -1.54747, 
    -1.543934, -1.539908, -1.535401, -1.530417, -1.524966, -1.519056, 
    -1.512695, -1.505893, -1.49866, -1.491006, -1.482942, -1.47448, -1.46563, 
    -1.456406, -1.446817, -1.436878, -1.4266, -1.415995, -1.405076, 
    -1.393856, -1.382348, -1.370563, -1.358514, -1.346213, -1.333673, 
    -1.320906, -1.307923, -1.294735, -1.281355, -1.267794, -1.254061, 
    -1.240168, -1.226125, -1.211942, -1.197629, -1.183195, -1.168648, 
    -1.153999, -1.139254, -1.124422, -1.109512,
  -0.3698378, -0.3748092, -0.3797542, -0.3846703, -0.3895547, -0.3944048, 
    -0.3992176, -0.40399, -0.4087191, -0.4134014, -0.4180338, -0.4226128, 
    -0.4271349, -0.4315965, -0.4359938, -0.4403231, -0.4445804, -0.448762, 
    -0.4528638, -0.4568816, -0.4608116, -0.4646493, -0.4683909, -0.472032, 
    -0.4755684, -0.478996, -0.4823107, -0.4855082, -0.4885846, -0.4915359, 
    -0.494358, -0.4970472, -0.4995998, -0.502012, -0.5042805, -0.5064019, 
    -0.5083731, -0.510191, -0.511853, -0.5133564, -0.5146989, -0.5158784, 
    -0.5168929, -0.5177408, -0.5184209, -0.5189319, -0.519273, -0.5194437, 
    -0.5194437, -0.519273, -0.5189319, -0.5184209, -0.5177408, -0.5168929, 
    -0.5158784, -0.5146989, -0.5133564, -0.511853, -0.510191, -0.5083731, 
    -0.5064019, -0.5042805, -0.502012, -0.4995998, -0.4970472, -0.494358, 
    -0.4915359, -0.4885846, -0.4855082, -0.4823107, -0.478996, -0.4755684, 
    -0.472032, -0.4683909, -0.4646493, -0.4608116, -0.4568816, -0.4528638, 
    -0.448762, -0.4445804, -0.4403231, -0.4359938, -0.4315965, -0.4271349, 
    -0.4226128, -0.4180338, -0.4134014, -0.4087191, -0.40399, -0.3992176, 
    -0.3944048, -0.3895547, -0.3846703, -0.3797542, -0.3748092, -0.3698378,
  0.3698378, 0.3748092, 0.3797542, 0.3846703, 0.3895547, 0.3944048, 
    0.3992176, 0.40399, 0.4087191, 0.4134014, 0.4180338, 0.4226128, 
    0.4271349, 0.4315965, 0.4359938, 0.4403231, 0.4445804, 0.448762, 
    0.4528638, 0.4568816, 0.4608116, 0.4646493, 0.4683909, 0.472032, 
    0.4755684, 0.478996, 0.4823107, 0.4855082, 0.4885846, 0.4915359, 
    0.494358, 0.4970472, 0.4995998, 0.502012, 0.5042805, 0.5064019, 
    0.5083731, 0.510191, 0.511853, 0.5133564, 0.5146989, 0.5158784, 
    0.5168929, 0.5177408, 0.5184209, 0.5189319, 0.519273, 0.5194437, 
    0.5194437, 0.519273, 0.5189319, 0.5184209, 0.5177408, 0.5168929, 
    0.5158784, 0.5146989, 0.5133564, 0.511853, 0.510191, 0.5083731, 
    0.5064019, 0.5042805, 0.502012, 0.4995998, 0.4970472, 0.494358, 
    0.4915359, 0.4885846, 0.4855082, 0.4823107, 0.478996, 0.4755684, 
    0.472032, 0.4683909, 0.4646493, 0.4608116, 0.4568816, 0.4528638, 
    0.448762, 0.4445804, 0.4403231, 0.4359938, 0.4315965, 0.4271349, 
    0.4226128, 0.4180338, 0.4134014, 0.4087191, 0.40399, 0.3992176, 
    0.3944048, 0.3895547, 0.3846703, 0.3797542, 0.3748092, 0.3698378,
  1.109512, 1.124422, 1.139254, 1.153999, 1.168648, 1.183195, 1.197629, 
    1.211942, 1.226125, 1.240168, 1.254061, 1.267794, 1.281355, 1.294735, 
    1.307923, 1.320906, 1.333673, 1.346213, 1.358514, 1.370563, 1.382348, 
    1.393856, 1.405076, 1.415995, 1.4266, 1.436878, 1.446817, 1.456406, 
    1.46563, 1.47448, 1.482942, 1.491006, 1.49866, 1.505893, 1.512695, 
    1.519056, 1.524966, 1.530417, 1.535401, 1.539908, 1.543934, 1.54747, 
    1.550512, 1.553055, 1.555094, 1.556626, 1.557649, 1.55816, 1.55816, 
    1.557649, 1.556626, 1.555094, 1.553055, 1.550512, 1.54747, 1.543934, 
    1.539908, 1.535401, 1.530417, 1.524966, 1.519056, 1.512695, 1.505893, 
    1.49866, 1.491006, 1.482942, 1.47448, 1.46563, 1.456406, 1.446817, 
    1.436878, 1.4266, 1.415995, 1.405076, 1.393856, 1.382348, 1.370563, 
    1.358514, 1.346213, 1.333673, 1.320906, 1.307923, 1.294735, 1.281355, 
    1.267794, 1.254061, 1.240168, 1.226125, 1.211942, 1.197629, 1.183195, 
    1.168648, 1.153999, 1.139254, 1.124422, 1.109512,
  1.849181, 1.87402, 1.898728, 1.92329, 1.947694, 1.971925, 1.995969, 
    2.019811, 2.043435, 2.066826, 2.089966, 2.112839, 2.135427, 2.157712, 
    2.179676, 2.201299, 2.222563, 2.243447, 2.263932, 2.283998, 2.303623, 
    2.322789, 2.341473, 2.359655, 2.377314, 2.394429, 2.41098, 2.426945, 
    2.442306, 2.457041, 2.471131, 2.484558, 2.497301, 2.509345, 2.52067, 
    2.53126, 2.541101, 2.550177, 2.558473, 2.565979, 2.57268, 2.578568, 
    2.583632, 2.587865, 2.59126, 2.593811, 2.595514, 2.596366, 2.596366, 
    2.595514, 2.593811, 2.59126, 2.587865, 2.583632, 2.578568, 2.57268, 
    2.565979, 2.558473, 2.550177, 2.541101, 2.53126, 2.52067, 2.509345, 
    2.497301, 2.484558, 2.471131, 2.457041, 2.442306, 2.426945, 2.41098, 
    2.394429, 2.377314, 2.359655, 2.341473, 2.322789, 2.303623, 2.283998, 
    2.263932, 2.243447, 2.222563, 2.201299, 2.179676, 2.157712, 2.135427, 
    2.112839, 2.089966, 2.066826, 2.043435, 2.019811, 1.995969, 1.971925, 
    1.947694, 1.92329, 1.898728, 1.87402, 1.849181,
  2.588841, 2.623593, 2.658159, 2.692521, 2.72666, 2.760556, 2.79419, 
    2.827541, 2.860586, 2.893303, 2.925669, 2.957661, 2.989253, 3.02042, 
    3.051136, 3.081377, 3.111113, 3.140318, 3.168964, 3.197022, 3.224465, 
    3.251263, 3.277388, 3.30281, 3.3275, 3.35143, 3.374569, 3.39689, 
    3.418365, 3.438965, 3.458663, 3.477432, 3.495247, 3.512082, 3.527913, 
    3.542717, 3.556473, 3.569159, 3.580756, 3.591246, 3.600614, 3.608843, 
    3.615922, 3.621838, 3.626583, 3.630148, 3.632529, 3.63372, 3.63372, 
    3.632529, 3.630148, 3.626583, 3.621838, 3.615922, 3.608843, 3.600614, 
    3.591246, 3.580756, 3.569159, 3.556473, 3.542717, 3.527913, 3.512082, 
    3.495247, 3.477432, 3.458663, 3.438965, 3.418365, 3.39689, 3.374569, 
    3.35143, 3.3275, 3.30281, 3.277388, 3.251263, 3.224465, 3.197022, 
    3.168964, 3.140318, 3.111113, 3.081377, 3.051136, 3.02042, 2.989253, 
    2.957661, 2.925669, 2.893303, 2.860586, 2.827541, 2.79419, 2.760556, 
    2.72666, 2.692521, 2.658159, 2.623593, 2.588841,
  3.32849, 3.37313, 3.41753, 3.461666, 3.505514, 3.549049, 3.592245, 
    3.635076, 3.677513, 3.719527, 3.761089, 3.802168, 3.842732, 3.88275, 
    3.922188, 3.961012, 3.999188, 4.036681, 4.073455, 4.109474, 4.144701, 
    4.179099, 4.212631, 4.245261, 4.27695, 4.307662, 4.337358, 4.366004, 
    4.393563, 4.419998, 4.445276, 4.46936, 4.49222, 4.513822, 4.534135, 
    4.55313, 4.570779, 4.587056, 4.601935, 4.615394, 4.627412, 4.63797, 
    4.647052, 4.654643, 4.660729, 4.665304, 4.668357, 4.669885, 4.669885, 
    4.668357, 4.665304, 4.660729, 4.654643, 4.647052, 4.63797, 4.627412, 
    4.615394, 4.601935, 4.587056, 4.570779, 4.55313, 4.534135, 4.513822, 
    4.49222, 4.46936, 4.445276, 4.419998, 4.393563, 4.366004, 4.337358, 
    4.307662, 4.27695, 4.245261, 4.212631, 4.179099, 4.144701, 4.109474, 
    4.073455, 4.036681, 3.999188, 3.961012, 3.922188, 3.88275, 3.842732, 
    3.802168, 3.761089, 3.719527, 3.677513, 3.635076, 3.592245, 3.549049, 
    3.505514, 3.461666, 3.41753, 3.37313, 3.32849,
  4.068124, 4.122622, 4.176824, 4.230701, 4.284225, 4.337364, 4.390087, 
    4.442361, 4.494153, 4.545426, 4.596145, 4.646272, 4.695769, 4.744597, 
    4.792715, 4.840082, 4.886656, 4.932395, 4.977254, 5.02119, 5.064158, 
    5.106114, 5.147013, 5.186808, 5.225454, 5.262908, 5.299122, 5.334054, 
    5.367657, 5.399891, 5.430711, 5.460076, 5.487947, 5.514283, 5.539048, 
    5.562205, 5.58372, 5.603562, 5.6217, 5.638107, 5.652757, 5.665627, 
    5.676696, 5.685948, 5.693368, 5.698944, 5.702665, 5.704528, 5.704528, 
    5.702665, 5.698944, 5.693368, 5.685948, 5.676696, 5.665627, 5.652757, 
    5.638107, 5.6217, 5.603562, 5.58372, 5.562205, 5.539048, 5.514283, 
    5.487947, 5.460076, 5.430711, 5.399891, 5.367657, 5.334054, 5.299122, 
    5.262908, 5.225454, 5.186808, 5.147013, 5.106114, 5.064158, 5.02119, 
    4.977254, 4.932395, 4.886656, 4.840082, 4.792715, 4.744597, 4.695769, 
    4.646272, 4.596145, 4.545426, 4.494153, 4.442361, 4.390087, 4.337364, 
    4.284225, 4.230701, 4.176824, 4.122622, 4.068124,
  4.807739, 4.872057, 4.936023, 4.999602, 5.06276, 5.125462, 5.187668, 
    5.249342, 5.310442, 5.370928, 5.430757, 5.489884, 5.548265, 5.605854, 
    5.662601, 5.718461, 5.773382, 5.827315, 5.880208, 5.93201, 5.982669, 
    6.032131, 6.080344, 6.127254, 6.172808, 6.216953, 6.259636, 6.300805, 
    6.340407, 6.378393, 6.414712, 6.449316, 6.482156, 6.513187, 6.542367, 
    6.56965, 6.594999, 6.618376, 6.639744, 6.659072, 6.676331, 6.691492, 
    6.704533, 6.715432, 6.724172, 6.73074, 6.735124, 6.737318, 6.737318, 
    6.735124, 6.73074, 6.724172, 6.715432, 6.704533, 6.691492, 6.676331, 
    6.659072, 6.639744, 6.618376, 6.594999, 6.56965, 6.542367, 6.513187, 
    6.482156, 6.449316, 6.414712, 6.378393, 6.340407, 6.300805, 6.259636, 
    6.216953, 6.172808, 6.127254, 6.080344, 6.032131, 5.982669, 5.93201, 
    5.880208, 5.827315, 5.773382, 5.718461, 5.662601, 5.605854, 5.548265, 
    5.489884, 5.430757, 5.370928, 5.310442, 5.249342, 5.187668, 5.125462, 
    5.06276, 4.999602, 4.936023, 4.872057, 4.807739,
  5.547333, 5.621428, 5.695111, 5.768345, 5.84109, 5.913303, 5.984942, 
    6.055964, 6.12632, 6.195964, 6.264847, 6.332918, 6.400125, 6.466415, 
    6.531734, 6.596026, 6.659235, 6.721301, 6.782168, 6.841775, 6.900063, 
    6.956971, 7.012438, 7.066403, 7.118805, 7.169584, 7.218679, 7.266029, 
    7.311576, 7.355261, 7.397027, 7.436818, 7.47458, 7.510261, 7.54381, 
    7.57518, 7.604323, 7.631198, 7.655765, 7.677984, 7.697824, 7.715252, 
    7.730243, 7.742771, 7.752818, 7.760367, 7.765407, 7.767929, 7.767929, 
    7.765407, 7.760367, 7.752818, 7.742771, 7.730243, 7.715252, 7.697824, 
    7.677984, 7.655765, 7.631198, 7.604323, 7.57518, 7.54381, 7.510261, 
    7.47458, 7.436818, 7.397027, 7.355261, 7.311576, 7.266029, 7.218679, 
    7.169584, 7.118805, 7.066403, 7.012438, 6.956971, 6.900063, 6.841775, 
    6.782168, 6.721301, 6.659235, 6.596026, 6.531734, 6.466415, 6.400125, 
    6.332918, 6.264847, 6.195964, 6.12632, 6.055964, 5.984942, 5.913303, 
    5.84109, 5.768345, 5.695111, 5.621428, 5.547333,
  6.286901, 6.370722, 6.454072, 6.536906, 6.619181, 6.70085, 6.781863, 
    6.862171, 6.941722, 7.020462, 7.098334, 7.175284, 7.251252, 7.326178, 
    7.4, 7.472656, 7.544083, 7.614214, 7.682984, 7.750327, 7.816175, 
    7.880459, 7.943112, 8.004064, 8.063247, 8.120593, 8.176033, 8.229501, 
    8.280929, 8.330251, 8.377405, 8.422327, 8.464956, 8.505234, 8.543103, 
    8.578511, 8.611405, 8.641738, 8.669463, 8.69454, 8.716929, 8.736598, 
    8.753514, 8.767653, 8.77899, 8.787509, 8.793196, 8.796041, 8.796041, 
    8.793196, 8.787509, 8.77899, 8.767653, 8.753514, 8.736598, 8.716929, 
    8.69454, 8.669463, 8.641738, 8.611405, 8.578511, 8.543103, 8.505234, 
    8.464956, 8.422327, 8.377405, 8.330251, 8.280929, 8.229501, 8.176033, 
    8.120593, 8.063247, 8.004064, 7.943112, 7.880459, 7.816175, 7.750327, 
    7.682984, 7.614214, 7.544083, 7.472656, 7.4, 7.326178, 7.251252, 
    7.175284, 7.098334, 7.020462, 6.941722, 6.862171, 6.781863, 6.70085, 
    6.619181, 6.536906, 6.454072, 6.370722, 6.286901,
  7.026442, 7.119931, 7.212887, 7.305261, 7.397004, 7.488063, 7.578384, 
    7.667912, 7.756588, 7.844352, 7.931143, 8.016898, 8.101551, 8.185037, 
    8.267286, 8.34823, 8.427797, 8.505915, 8.582511, 8.657512, 8.730841, 
    8.802423, 8.872184, 8.940046, 9.005934, 9.069772, 9.131484, 9.190996, 
    9.248235, 9.303126, 9.355601, 9.40559, 9.453025, 9.49784, 9.539974, 
    9.579368, 9.615962, 9.649706, 9.680549, 9.708443, 9.733348, 9.755226, 
    9.774042, 9.789767, 9.802377, 9.811852, 9.818177, 9.821342, 9.821342, 
    9.818177, 9.811852, 9.802377, 9.789767, 9.774042, 9.755226, 9.733348, 
    9.708443, 9.680549, 9.649706, 9.615962, 9.579368, 9.539974, 9.49784, 
    9.453025, 9.40559, 9.355601, 9.303126, 9.248235, 9.190996, 9.131484, 
    9.069772, 9.005934, 8.940046, 8.872184, 8.802423, 8.730841, 8.657512, 
    8.582511, 8.505915, 8.427797, 8.34823, 8.267286, 8.185037, 8.101551, 
    8.016898, 7.931143, 7.844352, 7.756588, 7.667912, 7.578384, 7.488063, 
    7.397004, 7.305261, 7.212887, 7.119931, 7.026442,
  7.765951, 7.869044, 7.971541, 8.073387, 8.174527, 8.274905, 8.37446, 
    8.473132, 8.570855, 8.667565, 8.763195, 8.857674, 8.95093, 9.042892, 
    9.133484, 9.222629, 9.31025, 9.396269, 9.480604, 9.563174, 9.643898, 
    9.722692, 9.799476, 9.874163, 9.946671, 10.01692, 10.08482, 10.1503, 
    10.21327, 10.27365, 10.33138, 10.38636, 10.43853, 10.48782, 10.53416, 
    10.57748, 10.61772, 10.65482, 10.68873, 10.7194, 10.74679, 10.77084, 
    10.79152, 10.80881, 10.82268, 10.83309, 10.84004, 10.84352, 10.84352, 
    10.84004, 10.83309, 10.82268, 10.80881, 10.79152, 10.77084, 10.74679, 
    10.7194, 10.68873, 10.65482, 10.61772, 10.57748, 10.53416, 10.48782, 
    10.43853, 10.38636, 10.33138, 10.27365, 10.21327, 10.1503, 10.08482, 
    10.01692, 9.946671, 9.874163, 9.799476, 9.722692, 9.643898, 9.563174, 
    9.480604, 9.396269, 9.31025, 9.222629, 9.133484, 9.042892, 8.95093, 
    8.857674, 8.763195, 8.667565, 8.570855, 8.473132, 8.37446, 8.274905, 
    8.174527, 8.073387, 7.971541, 7.869044, 7.765951,
  8.505425, 8.618052, 8.730017, 8.84126, 8.951721, 9.061338, 9.170046, 
    9.277779, 9.384465, 9.490034, 9.594414, 9.697527, 9.799295, 9.899641, 
    9.998483, 10.09574, 10.19132, 10.28514, 10.37712, 10.46716, 10.55519, 
    10.6411, 10.72481, 10.80623, 10.88527, 10.96183, 11.03584, 11.10719, 
    11.17581, 11.2416, 11.30449, 11.3644, 11.42123, 11.47492, 11.52539, 
    11.57257, 11.6164, 11.65681, 11.69374, 11.72714, 11.75696, 11.78315, 
    11.80567, 11.8245, 11.83959, 11.85093, 11.8585, 11.86229, 11.86229, 
    11.8585, 11.85093, 11.83959, 11.8245, 11.80567, 11.78315, 11.75696, 
    11.72714, 11.69374, 11.65681, 11.6164, 11.57257, 11.52539, 11.47492, 
    11.42123, 11.3644, 11.30449, 11.2416, 11.17581, 11.10719, 11.03584, 
    10.96183, 10.88527, 10.80623, 10.72481, 10.6411, 10.55519, 10.46716, 
    10.37712, 10.28514, 10.19132, 10.09574, 9.998483, 9.899641, 9.799295, 
    9.697527, 9.594414, 9.490034, 9.384465, 9.277779, 9.170046, 9.061338, 
    8.951721, 8.84126, 8.730017, 8.618052, 8.505425,
  9.244861, 9.366945, 9.488298, 9.608856, 9.728554, 9.847324, 9.965097, 
    10.0818, 10.19736, 10.31169, 10.42472, 10.53637, 10.64656, 10.75519, 
    10.86218, 10.96744, 11.07087, 11.1724, 11.27192, 11.36934, 11.46456, 
    11.55748, 11.64802, 11.73607, 11.82154, 11.90432, 11.98433, 12.06147, 
    12.13564, 12.20676, 12.27472, 12.33946, 12.40088, 12.45889, 12.51342, 
    12.5644, 12.61175, 12.6554, 12.6953, 12.73137, 12.76358, 12.79187, 
    12.8162, 12.83653, 12.85283, 12.86508, 12.87325, 12.87735, 12.87735, 
    12.87325, 12.86508, 12.85283, 12.83653, 12.8162, 12.79187, 12.76358, 
    12.73137, 12.6953, 12.6554, 12.61175, 12.5644, 12.51342, 12.45889, 
    12.40088, 12.33946, 12.27472, 12.20676, 12.13564, 12.06147, 11.98433, 
    11.90432, 11.82154, 11.73607, 11.64802, 11.55748, 11.46456, 11.36934, 
    11.27192, 11.1724, 11.07087, 10.96744, 10.86218, 10.75519, 10.64656, 
    10.53637, 10.42472, 10.31169, 10.19736, 10.0818, 9.965097, 9.847324, 
    9.728554, 9.608856, 9.488298, 9.366945, 9.244861,
  9.984256, 10.11571, 10.24637, 10.37615, 10.505, 10.63283, 10.75957, 
    10.88514, 11.00947, 11.13247, 11.25405, 11.37413, 11.49262, 11.60943, 
    11.72446, 11.83762, 11.9488, 12.05792, 12.16487, 12.26954, 12.37185, 
    12.47168, 12.56893, 12.66351, 12.75529, 12.84419, 12.9301, 13.01292, 
    13.09255, 13.16889, 13.24185, 13.31133, 13.37724, 13.43949, 13.49801, 
    13.55271, 13.60351, 13.65034, 13.69314, 13.73184, 13.76639, 13.79673, 
    13.82283, 13.84463, 13.86212, 13.87526, 13.88403, 13.88841, 13.88841, 
    13.88403, 13.87526, 13.86212, 13.84463, 13.82283, 13.79673, 13.76639, 
    13.73184, 13.69314, 13.65034, 13.60351, 13.55271, 13.49801, 13.43949, 
    13.37724, 13.31133, 13.24185, 13.16889, 13.09255, 13.01292, 12.9301, 
    12.84419, 12.75529, 12.66351, 12.56893, 12.47168, 12.37185, 12.26954, 
    12.16487, 12.05792, 11.9488, 11.83762, 11.72446, 11.60943, 11.49262, 
    11.37413, 11.25405, 11.13247, 11.00947, 10.88514, 10.75957, 10.63283, 
    10.505, 10.37615, 10.24637, 10.11571, 9.984256,
  10.72361, 10.86435, 11.00421, 11.14313, 11.28102, 11.41781, 11.55342, 
    11.68776, 11.82075, 11.9523, 12.08233, 12.21073, 12.33741, 12.46228, 
    12.58523, 12.70616, 12.82498, 12.94157, 13.05583, 13.16765, 13.27692, 
    13.38354, 13.48739, 13.58837, 13.68636, 13.78126, 13.87296, 13.96135, 
    14.04633, 14.1278, 14.20564, 14.27977, 14.35008, 14.4165, 14.47891, 
    14.53725, 14.59143, 14.64138, 14.68701, 14.72828, 14.76512, 14.79747, 
    14.8253, 14.84855, 14.86719, 14.88119, 14.89054, 14.89522, 14.89522, 
    14.89054, 14.88119, 14.86719, 14.84855, 14.8253, 14.79747, 14.76512, 
    14.72828, 14.68701, 14.64138, 14.59143, 14.53725, 14.47891, 14.4165, 
    14.35008, 14.27977, 14.20564, 14.1278, 14.04633, 13.96135, 13.87296, 
    13.78126, 13.68636, 13.58837, 13.48739, 13.38354, 13.27692, 13.16765, 
    13.05583, 12.94157, 12.82498, 12.70616, 12.58523, 12.46228, 12.33741, 
    12.21073, 12.08233, 11.9523, 11.82075, 11.68776, 11.55342, 11.41781, 
    11.28102, 11.14313, 11.00421, 10.86435, 10.72361,
  11.46291, 11.61284, 11.76182, 11.90976, 12.05659, 12.20224, 12.3466, 
    12.4896, 12.63114, 12.77113, 12.90947, 13.04607, 13.18083, 13.31363, 
    13.44438, 13.57297, 13.69929, 13.82323, 13.94467, 14.0635, 14.17962, 
    14.2929, 14.40323, 14.51049, 14.61457, 14.71535, 14.81272, 14.90658, 
    14.99679, 15.08327, 15.1659, 15.24457, 15.3192, 15.38967, 15.4559, 
    15.5178, 15.57528, 15.62826, 15.67667, 15.72045, 15.75952, 15.79384, 
    15.82335, 15.84801, 15.86777, 15.88263, 15.89254, 15.8975, 15.8975, 
    15.89254, 15.88263, 15.86777, 15.84801, 15.82335, 15.79384, 15.75952, 
    15.72045, 15.67667, 15.62826, 15.57528, 15.5178, 15.4559, 15.38967, 
    15.3192, 15.24457, 15.1659, 15.08327, 14.99679, 14.90658, 14.81272, 
    14.71535, 14.61457, 14.51049, 14.40323, 14.2929, 14.17962, 14.0635, 
    13.94467, 13.82323, 13.69929, 13.57297, 13.44438, 13.31363, 13.18083, 
    13.04607, 12.90947, 12.77113, 12.63114, 12.4896, 12.3466, 12.20224, 
    12.05659, 11.90976, 11.76182, 11.61284, 11.46291,
  12.20216, 12.36118, 12.51916, 12.67602, 12.83169, 12.98607, 13.13908, 
    13.29061, 13.44058, 13.58888, 13.73542, 13.88009, 14.02279, 14.1634, 
    14.30182, 14.43793, 14.57162, 14.70277, 14.83126, 14.95698, 15.07981, 
    15.19962, 15.31629, 15.42971, 15.53974, 15.64629, 15.74921, 15.8484, 
    15.94374, 16.03511, 16.12242, 16.20553, 16.28436, 16.3588, 16.42875, 
    16.49412, 16.55482, 16.61077, 16.66188, 16.7081, 16.74936, 16.78558, 
    16.81673, 16.84276, 16.86363, 16.87931, 16.88978, 16.89501, 16.89501, 
    16.88978, 16.87931, 16.86363, 16.84276, 16.81673, 16.78558, 16.74936, 
    16.7081, 16.66188, 16.61077, 16.55482, 16.49412, 16.42875, 16.3588, 
    16.28436, 16.20553, 16.12242, 16.03511, 15.94374, 15.8484, 15.74921, 
    15.64629, 15.53974, 15.42971, 15.31629, 15.19962, 15.07981, 14.95698, 
    14.83126, 14.70277, 14.57162, 14.43793, 14.30182, 14.1634, 14.02279, 
    13.88009, 13.73542, 13.58888, 13.44058, 13.29061, 13.13908, 12.98607, 
    12.83169, 12.67602, 12.51916, 12.36118, 12.20216,
  12.94136, 13.10935, 13.27623, 13.4419, 13.60628, 13.76928, 13.9308, 
    14.09074, 14.24901, 14.4055, 14.56011, 14.71272, 14.86322, 15.0115, 
    15.15745, 15.30094, 15.44186, 15.58009, 15.71549, 15.84795, 15.97735, 
    16.10355, 16.22643, 16.34587, 16.46173, 16.57389, 16.68224, 16.78664, 
    16.88698, 16.98314, 17.075, 17.16244, 17.24537, 17.32367, 17.39725, 
    17.466, 17.52983, 17.58866, 17.64242, 17.69101, 17.73438, 17.77247, 
    17.80522, 17.83258, 17.85452, 17.871, 17.882, 17.88751, 17.88751, 17.882, 
    17.871, 17.85452, 17.83258, 17.80522, 17.77247, 17.73438, 17.69101, 
    17.64242, 17.58866, 17.52983, 17.466, 17.39725, 17.32367, 17.24537, 
    17.16244, 17.075, 16.98314, 16.88698, 16.78664, 16.68224, 16.57389, 
    16.46173, 16.34587, 16.22643, 16.10355, 15.97735, 15.84795, 15.71549, 
    15.58009, 15.44186, 15.30094, 15.15745, 15.0115, 14.86322, 14.71272, 
    14.56011, 14.4055, 14.24901, 14.09074, 13.9308, 13.76928, 13.60628, 
    13.4419, 13.27623, 13.10935, 12.94136,
  13.6805, 13.85736, 14.03301, 14.20737, 14.38034, 14.55183, 14.72173, 
    14.88996, 15.05639, 15.22093, 15.38346, 15.54386, 15.70203, 15.85784, 
    16.01117, 16.1619, 16.30991, 16.45506, 16.59723, 16.73629, 16.87211, 
    17.00456, 17.1335, 17.25882, 17.38036, 17.49802, 17.61165, 17.72114, 
    17.82635, 17.92716, 18.02345, 18.11512, 18.20203, 18.28409, 18.36119, 
    18.43323, 18.50011, 18.56174, 18.61805, 18.66896, 18.71439, 18.75428, 
    18.78858, 18.81724, 18.84021, 18.85747, 18.86899, 18.87476, 18.87476, 
    18.86899, 18.85747, 18.84021, 18.81724, 18.78858, 18.75428, 18.71439, 
    18.66896, 18.61805, 18.56174, 18.50011, 18.43323, 18.36119, 18.28409, 
    18.20203, 18.11512, 18.02345, 17.92716, 17.82635, 17.72114, 17.61165, 
    17.49802, 17.38036, 17.25882, 17.1335, 17.00456, 16.87211, 16.73629, 
    16.59723, 16.45506, 16.30991, 16.1619, 16.01117, 15.85784, 15.70203, 
    15.54386, 15.38346, 15.22093, 15.05639, 14.88996, 14.72173, 14.55183, 
    14.38034, 14.20737, 14.03301, 13.85736, 13.6805,
  14.41959, 14.60518, 14.78949, 14.9724, 15.15383, 15.33368, 15.51184, 
    15.6882, 15.86266, 16.0351, 16.20541, 16.37346, 16.53915, 16.70233, 
    16.8629, 17.02072, 17.17565, 17.32758, 17.47636, 17.62187, 17.76396, 
    17.9025, 18.03736, 18.16841, 18.2955, 18.4185, 18.53728, 18.65171, 
    18.76166, 18.867, 18.96761, 19.06337, 19.15416, 19.23986, 19.32038, 
    19.39561, 19.46544, 19.5298, 19.58859, 19.64173, 19.68916, 19.7308, 
    19.7666, 19.79651, 19.82049, 19.8385, 19.85053, 19.85655, 19.85655, 
    19.85053, 19.8385, 19.82049, 19.79651, 19.7666, 19.7308, 19.68916, 
    19.64173, 19.58859, 19.5298, 19.46544, 19.39561, 19.32038, 19.23986, 
    19.15416, 19.06337, 18.96761, 18.867, 18.76166, 18.65171, 18.53728, 
    18.4185, 18.2955, 18.16841, 18.03736, 17.9025, 17.76396, 17.62187, 
    17.47636, 17.32758, 17.17565, 17.02072, 16.8629, 16.70233, 16.53915, 
    16.37346, 16.20541, 16.0351, 15.86266, 15.6882, 15.51184, 15.33368, 
    15.15383, 14.9724, 14.78949, 14.60518, 14.41959,
  15.15861, 15.35282, 15.54564, 15.73699, 15.92674, 16.11481, 16.30107, 
    16.48543, 16.66776, 16.84796, 17.02589, 17.20144, 17.37449, 17.5449, 
    17.71254, 17.87728, 18.03899, 18.19754, 18.35277, 18.50457, 18.65277, 
    18.79726, 18.93789, 19.07451, 19.20699, 19.33519, 19.45897, 19.57821, 
    19.69276, 19.8025, 19.90729, 20.00702, 20.10156, 20.19081, 20.27464, 
    20.35295, 20.42565, 20.49264, 20.55383, 20.60913, 20.65849, 20.70182, 
    20.73908, 20.7702, 20.79515, 20.81389, 20.8264, 20.83266, 20.83266, 
    20.8264, 20.81389, 20.79515, 20.7702, 20.73908, 20.70182, 20.65849, 
    20.60913, 20.55383, 20.49264, 20.42565, 20.35295, 20.27464, 20.19081, 
    20.10156, 20.00702, 19.90729, 19.8025, 19.69276, 19.57821, 19.45897, 
    19.33519, 19.20699, 19.07451, 18.93789, 18.79726, 18.65277, 18.50457, 
    18.35277, 18.19754, 18.03899, 17.87728, 17.71254, 17.5449, 17.37449, 
    17.20144, 17.02589, 16.84796, 16.66776, 16.48543, 16.30107, 16.11481, 
    15.92674, 15.73699, 15.54564, 15.35282, 15.15861,
  15.89756, 16.10026, 16.30147, 16.50109, 16.69903, 16.89517, 17.0894, 
    17.2816, 17.47165, 17.65945, 17.84485, 18.02774, 18.20799, 18.38545, 
    18.56001, 18.73152, 18.89984, 19.06483, 19.22636, 19.38427, 19.53844, 
    19.68871, 19.83493, 19.97698, 20.11469, 20.24794, 20.37659, 20.50048, 
    20.61949, 20.73348, 20.84233, 20.94591, 21.04409, 21.13675, 21.22379, 
    21.30509, 21.38055, 21.45008, 21.51358, 21.57098, 21.6222, 21.66716, 
    21.70582, 21.73811, 21.764, 21.78345, 21.79643, 21.80292, 21.80292, 
    21.79643, 21.78345, 21.764, 21.73811, 21.70582, 21.66716, 21.6222, 
    21.57098, 21.51358, 21.45008, 21.38055, 21.30509, 21.22379, 21.13675, 
    21.04409, 20.94591, 20.84233, 20.73348, 20.61949, 20.50048, 20.37659, 
    20.24794, 20.11469, 19.97698, 19.83493, 19.68871, 19.53844, 19.38427, 
    19.22636, 19.06483, 18.89984, 18.73152, 18.56001, 18.38545, 18.20799, 
    18.02774, 17.84485, 17.65945, 17.47165, 17.2816, 17.0894, 16.89517, 
    16.69903, 16.50109, 16.30147, 16.10026, 15.89756,
  16.63645, 16.84749, 17.05695, 17.26471, 17.47068, 17.67474, 17.87678, 
    18.07666, 18.27429, 18.46952, 18.66223, 18.85229, 19.03956, 19.22392, 
    19.40522, 19.58332, 19.75808, 19.92936, 20.09701, 20.26088, 20.42083, 
    20.57672, 20.72838, 20.87569, 21.01848, 21.15662, 21.28997, 21.41838, 
    21.5417, 21.65982, 21.77258, 21.87987, 21.98156, 22.07753, 22.16766, 
    22.25184, 22.32997, 22.40195, 22.46768, 22.52709, 22.5801, 22.62664, 
    22.66665, 22.70007, 22.72686, 22.74698, 22.76041, 22.76713, 22.76713, 
    22.76041, 22.74698, 22.72686, 22.70007, 22.66665, 22.62664, 22.5801, 
    22.52709, 22.46768, 22.40195, 22.32997, 22.25184, 22.16766, 22.07753, 
    21.98156, 21.87987, 21.77258, 21.65982, 21.5417, 21.41838, 21.28997, 
    21.15662, 21.01848, 20.87569, 20.72838, 20.57672, 20.42083, 20.26088, 
    20.09701, 19.92936, 19.75808, 19.58332, 19.40522, 19.22392, 19.03956, 
    18.85229, 18.66223, 18.46952, 18.27429, 18.07666, 17.87678, 17.67474, 
    17.47068, 17.26471, 17.05695, 16.84749, 16.63645,
  17.37526, 17.59451, 17.81206, 18.02782, 18.24167, 18.45349, 18.66317, 
    18.87058, 19.07561, 19.2781, 19.47795, 19.67501, 19.86915, 20.06023, 
    20.2481, 20.43262, 20.61365, 20.79103, 20.96463, 21.13428, 21.29985, 
    21.46118, 21.61812, 21.77052, 21.91823, 22.0611, 22.19899, 22.33176, 
    22.45926, 22.58134, 22.69789, 22.80877, 22.91384, 23.01299, 23.10609, 
    23.19304, 23.27374, 23.34808, 23.41596, 23.47731, 23.53204, 23.58009, 
    23.62139, 23.6559, 23.68355, 23.70432, 23.71819, 23.72513, 23.72513, 
    23.71819, 23.70432, 23.68355, 23.6559, 23.62139, 23.58009, 23.53204, 
    23.47731, 23.41596, 23.34808, 23.27374, 23.19304, 23.10609, 23.01299, 
    22.91384, 22.80877, 22.69789, 22.58134, 22.45926, 22.33176, 22.19899, 
    22.0611, 21.91823, 21.77052, 21.61812, 21.46118, 21.29985, 21.13428, 
    20.96463, 20.79103, 20.61365, 20.43262, 20.2481, 20.06023, 19.86915, 
    19.67501, 19.47795, 19.2781, 19.07561, 18.87058, 18.66317, 18.45349, 
    18.24167, 18.02782, 17.81206, 17.59451, 17.37526,
  18.114, 18.3413, 18.5668, 18.79039, 19.01196, 19.23139, 19.44855, 19.66332, 
    19.87557, 20.08517, 20.29198, 20.49586, 20.69669, 20.8943, 21.08856, 
    21.27932, 21.46644, 21.64975, 21.82912, 22.00438, 22.17539, 22.34199, 
    22.50403, 22.66135, 22.81381, 22.96125, 23.10353, 23.2405, 23.37202, 
    23.49794, 23.61813, 23.73245, 23.84077, 23.94298, 24.03895, 24.12856, 
    24.21172, 24.28832, 24.35827, 24.42147, 24.47786, 24.52736, 24.5699, 
    24.60544, 24.63392, 24.65532, 24.6696, 24.67674, 24.67674, 24.6696, 
    24.65532, 24.63392, 24.60544, 24.5699, 24.52736, 24.47786, 24.42147, 
    24.35827, 24.28832, 24.21172, 24.12856, 24.03895, 23.94298, 23.84077, 
    23.73245, 23.61813, 23.49794, 23.37202, 23.2405, 23.10353, 22.96125, 
    22.81381, 22.66135, 22.50403, 22.34199, 22.17539, 22.00438, 21.82912, 
    21.64975, 21.46644, 21.27932, 21.08856, 20.8943, 20.69669, 20.49586, 
    20.29198, 20.08517, 19.87557, 19.66332, 19.44855, 19.23139, 19.01196, 
    18.79039, 18.5668, 18.3413, 18.114,
  18.85267, 19.08786, 19.32115, 19.55242, 19.78154, 20.0084, 20.23287, 
    20.45482, 20.67413, 20.89065, 21.10424, 21.31477, 21.52209, 21.72607, 
    21.92654, 22.12335, 22.31637, 22.50543, 22.69039, 22.87107, 23.04734, 
    23.21904, 23.386, 23.54808, 23.70512, 23.85697, 24.00347, 24.14449, 
    24.27987, 24.40947, 24.53315, 24.65079, 24.76223, 24.86737, 24.96609, 
    25.05826, 25.14377, 25.22254, 25.29446, 25.35944, 25.41741, 25.46829, 
    25.51202, 25.54855, 25.57783, 25.59982, 25.6145, 25.62184, 25.62184, 
    25.6145, 25.59982, 25.57783, 25.54855, 25.51202, 25.46829, 25.41741, 
    25.35944, 25.29446, 25.22254, 25.14377, 25.05826, 24.96609, 24.86737, 
    24.76223, 24.65079, 24.53315, 24.40947, 24.27987, 24.14449, 24.00347, 
    23.85697, 23.70512, 23.54808, 23.386, 23.21904, 23.04734, 22.87107, 
    22.69039, 22.50543, 22.31637, 22.12335, 21.92654, 21.72607, 21.52209, 
    21.31477, 21.10424, 20.89065, 20.67413, 20.45482, 20.23287, 20.0084, 
    19.78154, 19.55242, 19.32115, 19.08786, 18.85267,
  19.59126, 19.83419, 20.0751, 20.31387, 20.55038, 20.7845, 21.01611, 
    21.24507, 21.47124, 21.6945, 21.91469, 22.13168, 22.34532, 22.55546, 
    22.76195, 22.96464, 23.16337, 23.35799, 23.54835, 23.73428, 23.91562, 
    24.09223, 24.26394, 24.43059, 24.59204, 24.74813, 24.89869, 25.04359, 
    25.18268, 25.31582, 25.44285, 25.56366, 25.6781, 25.78605, 25.88738, 
    25.98199, 26.06977, 26.1506, 26.2244, 26.29108, 26.35056, 26.40276, 
    26.44763, 26.4851, 26.51514, 26.5377, 26.55275, 26.56029, 26.56029, 
    26.55275, 26.5377, 26.51514, 26.4851, 26.44763, 26.40276, 26.35056, 
    26.29108, 26.2244, 26.1506, 26.06977, 25.98199, 25.88738, 25.78605, 
    25.6781, 25.56366, 25.44285, 25.31582, 25.18268, 25.04359, 24.89869, 
    24.74813, 24.59204, 24.43059, 24.26394, 24.09223, 23.91562, 23.73428, 
    23.54835, 23.35799, 23.16337, 22.96464, 22.76195, 22.55546, 22.34532, 
    22.13168, 21.91469, 21.6945, 21.47124, 21.24507, 21.01611, 20.7845, 
    20.55038, 20.31387, 20.0751, 19.83419, 19.59126,
  20.32976, 20.58027, 20.82863, 21.07474, 21.31846, 21.55966, 21.79822, 
    22.034, 22.26687, 22.49667, 22.72328, 22.94654, 23.1663, 23.38242, 
    23.59474, 23.8031, 24.00736, 24.20735, 24.40292, 24.5939, 24.78014, 
    24.96147, 25.13775, 25.3088, 25.47448, 25.63463, 25.78909, 25.93772, 
    26.08036, 26.21687, 26.34712, 26.47095, 26.58825, 26.69888, 26.80272, 
    26.89966, 26.98958, 27.07239, 27.14798, 27.21628, 27.27719, 27.33065, 
    27.3766, 27.41497, 27.44572, 27.46882, 27.48424, 27.49195, 27.49195, 
    27.48424, 27.46882, 27.44572, 27.41497, 27.3766, 27.33065, 27.27719, 
    27.21628, 27.14798, 27.07239, 26.98958, 26.89966, 26.80272, 26.69888, 
    26.58825, 26.47095, 26.34712, 26.21687, 26.08036, 25.93772, 25.78909, 
    25.63463, 25.47448, 25.3088, 25.13775, 24.96147, 24.78014, 24.5939, 
    24.40292, 24.20735, 24.00736, 23.8031, 23.59474, 23.38242, 23.1663, 
    22.94654, 22.72328, 22.49667, 22.26687, 22.034, 21.79822, 21.55966, 
    21.31846, 21.07474, 20.82863, 20.58027, 20.32976,
  21.06818, 21.32609, 21.58174, 21.835, 22.08575, 22.33386, 22.57919, 
    22.8216, 23.06096, 23.29713, 23.52995, 23.75929, 23.98498, 24.20688, 
    24.42483, 24.63868, 24.84826, 25.05343, 25.25401, 25.44986, 25.6408, 
    25.82668, 26.00734, 26.18261, 26.35234, 26.51638, 26.67457, 26.82676, 
    26.9728, 27.11254, 27.24584, 27.37256, 27.49258, 27.60576, 27.71199, 
    27.81114, 27.90311, 27.98779, 28.06509, 28.13491, 28.19719, 28.25185, 
    28.29881, 28.33804, 28.36947, 28.39308, 28.40884, 28.41672, 28.41672, 
    28.40884, 28.39308, 28.36947, 28.33804, 28.29881, 28.25185, 28.19719, 
    28.13491, 28.06509, 27.98779, 27.90311, 27.81114, 27.71199, 27.60576, 
    27.49258, 27.37256, 27.24584, 27.11254, 26.9728, 26.82676, 26.67457, 
    26.51638, 26.35234, 26.18261, 26.00734, 25.82668, 25.6408, 25.44986, 
    25.25401, 25.05343, 24.84826, 24.63868, 24.42483, 24.20688, 23.98498, 
    23.75929, 23.52995, 23.29713, 23.06096, 22.8216, 22.57919, 22.33386, 
    22.08575, 21.835, 21.58174, 21.32609, 21.06818,
  21.80651, 22.07165, 22.33441, 22.59464, 22.85224, 23.10706, 23.35897, 
    23.60783, 23.85349, 24.09582, 24.33467, 24.56988, 24.8013, 25.02878, 
    25.25217, 25.4713, 25.68602, 25.89616, 26.10157, 26.30208, 26.49753, 
    26.68777, 26.87262, 27.05193, 27.22555, 27.3933, 27.55505, 27.71063, 
    27.8599, 28.00271, 28.13892, 28.2684, 28.391, 28.50661, 28.6151, 
    28.71634, 28.81025, 28.89671, 28.97562, 29.0469, 29.11047, 29.16625, 
    29.21418, 29.25421, 29.28629, 29.31038, 29.32646, 29.33451, 29.33451, 
    29.32646, 29.31038, 29.28629, 29.25421, 29.21418, 29.16625, 29.11047, 
    29.0469, 28.97562, 28.89671, 28.81025, 28.71634, 28.6151, 28.50661, 
    28.391, 28.2684, 28.13892, 28.00271, 27.8599, 27.71063, 27.55505, 
    27.3933, 27.22555, 27.05193, 26.87262, 26.68777, 26.49753, 26.30208, 
    26.10157, 25.89616, 25.68602, 25.4713, 25.25217, 25.02878, 24.8013, 
    24.56988, 24.33467, 24.09582, 23.85349, 23.60783, 23.35897, 23.10706, 
    22.85224, 22.59464, 22.33441, 22.07165, 21.80651,
  22.54476, 22.81695, 23.08662, 23.35365, 23.6179, 23.87924, 24.13754, 
    24.39264, 24.64441, 24.89271, 25.13737, 25.37826, 25.61521, 25.84807, 
    26.07669, 26.30091, 26.52055, 26.73548, 26.94551, 27.1505, 27.35027, 
    27.54466, 27.73353, 27.91669, 28.094, 28.2653, 28.43043, 28.58924, 
    28.74158, 28.88731, 29.02629, 29.15837, 29.28342, 29.40132, 29.51195, 
    29.61518, 29.71092, 29.79905, 29.87949, 29.95214, 30.01692, 30.07377, 
    30.12261, 30.1634, 30.19609, 30.22064, 30.23702, 30.24521, 30.24521, 
    30.23702, 30.22064, 30.19609, 30.1634, 30.12261, 30.07377, 30.01692, 
    29.95214, 29.87949, 29.79905, 29.71092, 29.61518, 29.51195, 29.40132, 
    29.28342, 29.15837, 29.02629, 28.88731, 28.74158, 28.58924, 28.43043, 
    28.2653, 28.094, 27.91669, 27.73353, 27.54466, 27.35027, 27.1505, 
    26.94551, 26.73548, 26.52055, 26.30091, 26.07669, 25.84807, 25.61521, 
    25.37826, 25.13737, 24.89271, 24.64441, 24.39264, 24.13754, 23.87924, 
    23.6179, 23.35365, 23.08662, 22.81695, 22.54476,
  23.28291, 23.56197, 23.83837, 24.112, 24.38272, 24.65038, 24.91487, 
    25.17602, 25.43369, 25.68774, 25.93803, 26.18438, 26.42666, 26.6647, 
    26.89834, 27.12744, 27.35181, 27.57131, 27.78577, 27.99503, 28.19893, 
    28.3973, 28.58998, 28.77681, 28.95764, 29.1323, 29.30065, 29.46252, 
    29.61777, 29.76627, 29.90785, 30.04239, 30.16976, 30.28983, 30.40247, 
    30.50758, 30.60504, 30.69475, 30.77662, 30.85055, 30.91648, 30.97433, 
    31.02403, 31.06553, 31.09879, 31.12376, 31.14043, 31.14876, 31.14876, 
    31.14043, 31.12376, 31.09879, 31.06553, 31.02403, 30.97433, 30.91648, 
    30.85055, 30.77662, 30.69475, 30.60504, 30.50758, 30.40247, 30.28983, 
    30.16976, 30.04239, 29.90785, 29.76627, 29.61777, 29.46252, 29.30065, 
    29.1323, 28.95764, 28.77681, 28.58998, 28.3973, 28.19893, 27.99503, 
    27.78577, 27.57131, 27.35181, 27.12744, 26.89834, 26.6647, 26.42666, 
    26.18438, 25.93803, 25.68774, 25.43369, 25.17602, 24.91487, 24.65038, 
    24.38272, 24.112, 23.83837, 23.56197, 23.28291,
  24.02097, 24.3067, 24.58965, 24.86968, 25.14667, 25.42046, 25.69092, 
    25.95792, 26.22129, 26.4809, 26.73659, 26.98821, 27.2356, 27.47861, 
    27.71707, 27.95084, 28.17974, 28.40361, 28.6223, 28.83563, 29.04346, 
    29.2456, 29.44192, 29.63223, 29.81639, 29.99424, 30.16563, 30.3304, 
    30.4884, 30.6395, 30.78355, 30.92041, 31.04995, 31.17205, 31.28659, 
    31.39346, 31.49253, 31.58372, 31.66694, 31.74208, 31.80908, 31.86786, 
    31.91836, 31.96053, 31.99432, 32.01969, 32.03662, 32.04509, 32.04509, 
    32.03662, 32.01969, 31.99432, 31.96053, 31.91836, 31.86786, 31.80908, 
    31.74208, 31.66694, 31.58372, 31.49253, 31.39346, 31.28659, 31.17205, 
    31.04995, 30.92041, 30.78355, 30.6395, 30.4884, 30.3304, 30.16563, 
    29.99424, 29.81639, 29.63223, 29.44192, 29.2456, 29.04346, 28.83563, 
    28.6223, 28.40361, 28.17974, 27.95084, 27.71707, 27.47861, 27.2356, 
    26.98821, 26.73659, 26.4809, 26.22129, 25.95792, 25.69092, 25.42046, 
    25.14667, 24.86968, 24.58965, 24.3067, 24.02097,
  24.75893, 25.05115, 25.34044, 25.62668, 25.90973, 26.18944, 26.46569, 
    26.73832, 27.00718, 27.27213, 27.53302, 27.78969, 28.04199, 28.28975, 
    28.53283, 28.77106, 29.00427, 29.23232, 29.45502, 29.67224, 29.88379, 
    30.08952, 30.28927, 30.48288, 30.6702, 30.85106, 31.02531, 31.19281, 
    31.3534, 31.50695, 31.65331, 31.79235, 31.92393, 32.04794, 32.16426, 
    32.27277, 32.37335, 32.46593, 32.55039, 32.62666, 32.69466, 32.75431, 
    32.80555, 32.84834, 32.88263, 32.90837, 32.92555, 32.93415, 32.93415, 
    32.92555, 32.90837, 32.88263, 32.84834, 32.80555, 32.75431, 32.69466, 
    32.62666, 32.55039, 32.46593, 32.37335, 32.27277, 32.16426, 32.04794, 
    31.92393, 31.79235, 31.65331, 31.50695, 31.3534, 31.19281, 31.02531, 
    30.85106, 30.6702, 30.48288, 30.28927, 30.08952, 29.88379, 29.67224, 
    29.45502, 29.23232, 29.00427, 28.77106, 28.53283, 28.28975, 28.04199, 
    27.78969, 27.53302, 27.27213, 27.00718, 26.73832, 26.46569, 26.18944, 
    25.90973, 25.62668, 25.34044, 25.05115, 24.75893,
  25.4968, 25.7953, 26.09074, 26.38298, 26.67189, 26.95732, 27.23913, 
    27.51719, 27.79133, 28.06141, 28.32729, 28.5888, 28.84579, 29.0981, 
    29.34557, 29.58805, 29.82537, 30.05738, 30.28391, 30.50479, 30.71988, 
    30.929, 31.132, 31.32872, 31.519, 31.70269, 31.87964, 32.0497, 32.21272, 
    32.36856, 32.51709, 32.65816, 32.79165, 32.91744, 33.03541, 33.14545, 
    33.24744, 33.3413, 33.42693, 33.50424, 33.57316, 33.63363, 33.68556, 
    33.72892, 33.76367, 33.78976, 33.80717, 33.81588, 33.81588, 33.80717, 
    33.78976, 33.76367, 33.72892, 33.68556, 33.63363, 33.57316, 33.50424, 
    33.42693, 33.3413, 33.24744, 33.14545, 33.03541, 32.91744, 32.79165, 
    32.65816, 32.51709, 32.36856, 32.21272, 32.0497, 31.87964, 31.70269, 
    31.519, 31.32872, 31.132, 30.929, 30.71988, 30.50479, 30.28391, 30.05738, 
    29.82537, 29.58805, 29.34557, 29.0981, 28.84579, 28.5888, 28.32729, 
    28.06141, 27.79133, 27.51719, 27.23913, 26.95732, 26.67189, 26.38298, 
    26.09074, 25.7953, 25.4968,
  26.23456, 26.53915, 26.84053, 27.13857, 27.43312, 27.72406, 28.01123, 
    28.29449, 28.5737, 28.84871, 29.11935, 29.38548, 29.64695, 29.90359, 
    30.15525, 30.40177, 30.643, 30.87876, 31.10889, 31.33325, 31.55167, 
    31.76398, 31.97004, 32.16968, 32.36275, 32.5491, 32.72858, 32.90103, 
    33.06631, 33.2243, 33.37484, 33.5178, 33.65307, 33.78051, 33.90001, 
    34.01146, 34.11476, 34.20981, 34.29651, 34.37479, 34.44456, 34.50577, 
    34.55835, 34.60224, 34.63741, 34.66381, 34.68143, 34.69025, 34.69025, 
    34.68143, 34.66381, 34.63741, 34.60224, 34.55835, 34.50577, 34.44456, 
    34.37479, 34.29651, 34.20981, 34.11476, 34.01146, 33.90001, 33.78051, 
    33.65307, 33.5178, 33.37484, 33.2243, 33.06631, 32.90103, 32.72858, 
    32.5491, 32.36275, 32.16968, 31.97004, 31.76398, 31.55167, 31.33325, 
    31.10889, 30.87876, 30.643, 30.40177, 30.15525, 29.90359, 29.64695, 
    29.38548, 29.11935, 28.84871, 28.5737, 28.29449, 28.01123, 27.72406, 
    27.43312, 27.13857, 26.84053, 26.53915, 26.23456,
  26.97222, 27.28269, 27.58981, 27.89343, 28.19342, 28.48965, 28.78197, 
    29.07022, 29.35428, 29.63398, 29.90917, 30.17971, 30.44544, 30.7062, 
    30.96183, 31.21218, 31.45709, 31.6964, 31.92994, 32.15757, 32.37912, 
    32.59444, 32.80336, 33.00574, 33.20141, 33.39024, 33.57207, 33.74675, 
    33.91414, 34.07411, 34.22652, 34.37123, 34.50814, 34.6371, 34.75802, 
    34.87078, 34.97528, 35.07141, 35.15911, 35.23827, 35.30883, 35.37072, 
    35.42388, 35.46826, 35.50381, 35.53051, 35.54832, 35.55723, 35.55723, 
    35.54832, 35.53051, 35.50381, 35.46826, 35.42388, 35.37072, 35.30883, 
    35.23827, 35.15911, 35.07141, 34.97528, 34.87078, 34.75802, 34.6371, 
    34.50814, 34.37123, 34.22652, 34.07411, 33.91414, 33.74675, 33.57207, 
    33.39024, 33.20141, 33.00574, 32.80336, 32.59444, 32.37912, 32.15757, 
    31.92994, 31.6964, 31.45709, 31.21218, 30.96183, 30.7062, 30.44544, 
    30.17971, 29.90917, 29.63398, 29.35428, 29.07022, 28.78197, 28.48965, 
    28.19342, 27.89343, 27.58981, 27.28269, 26.97222,
  27.70978, 28.02592, 28.33856, 28.64755, 28.95277, 29.25407, 29.55131, 
    29.84434, 30.13302, 30.4172, 30.69673, 30.97146, 31.24123, 31.50589, 
    31.76528, 32.01924, 32.26763, 32.51027, 32.74702, 32.97771, 33.2022, 
    33.42032, 33.63192, 33.83684, 34.03494, 34.22607, 34.41008, 34.58682, 
    34.75616, 34.91797, 35.0721, 35.21843, 35.35684, 35.48721, 35.60942, 
    35.72337, 35.82896, 35.9261, 36.01469, 36.09467, 36.16594, 36.22845, 
    36.28214, 36.32696, 36.36287, 36.38982, 36.40781, 36.41681, 36.41681, 
    36.40781, 36.38982, 36.36287, 36.32696, 36.28214, 36.22845, 36.16594, 
    36.09467, 36.01469, 35.9261, 35.82896, 35.72337, 35.60942, 35.48721, 
    35.35684, 35.21843, 35.0721, 34.91797, 34.75616, 34.58682, 34.41008, 
    34.22607, 34.03494, 33.83684, 33.63192, 33.42032, 33.2022, 32.97771, 
    32.74702, 32.51027, 32.26763, 32.01924, 31.76528, 31.50589, 31.24123, 
    30.97146, 30.69673, 30.4172, 30.13302, 29.84434, 29.55131, 29.25407, 
    28.95277, 28.64755, 28.33856, 28.02592, 27.70978,
  28.44723, 28.76883, 29.08677, 29.40093, 29.71115, 30.0173, 30.31924, 
    30.61683, 30.90992, 31.19835, 31.482, 31.76069, 32.03428, 32.30262, 
    32.56555, 32.82292, 33.07457, 33.32034, 33.56009, 33.79364, 34.02087, 
    34.2416, 34.45568, 34.66297, 34.86331, 35.05656, 35.24258, 35.42123, 
    35.59236, 35.75585, 35.91155, 36.05936, 36.19914, 36.33079, 36.45418, 
    36.56922, 36.67581, 36.77385, 36.86326, 36.94396, 37.01588, 37.07895, 
    37.13312, 37.17834, 37.21456, 37.24176, 37.2599, 37.26898, 37.26898, 
    37.2599, 37.24176, 37.21456, 37.17834, 37.13312, 37.07895, 37.01588, 
    36.94396, 36.86326, 36.77385, 36.67581, 36.56922, 36.45418, 36.33079, 
    36.19914, 36.05936, 35.91155, 35.75585, 35.59236, 35.42123, 35.24258, 
    35.05656, 34.86331, 34.66297, 34.45568, 34.2416, 34.02087, 33.79364, 
    33.56009, 33.32034, 33.07457, 32.82292, 32.56555, 32.30262, 32.03428, 
    31.76069, 31.482, 31.19835, 30.90992, 30.61683, 30.31924, 30.0173, 
    29.71115, 29.40093, 29.08677, 28.76883, 28.44723,
  29.18457, 29.51142, 29.83445, 30.15354, 30.46854, 30.77932, 31.08575, 
    31.38766, 31.68493, 31.97741, 32.26494, 32.54737, 32.82457, 33.09637, 
    33.36263, 33.62318, 33.87788, 34.12658, 34.36911, 34.60533, 34.83509, 
    35.05824, 35.27462, 35.48409, 35.68649, 35.8817, 36.06956, 36.24994, 
    36.42271, 36.58773, 36.74487, 36.89401, 37.03504, 37.16784, 37.2923, 
    37.40832, 37.5158, 37.61465, 37.7048, 37.78615, 37.85865, 37.92222, 
    37.97682, 38.02239, 38.0589, 38.0863, 38.10459, 38.11374, 38.11374, 
    38.10459, 38.0863, 38.0589, 38.02239, 37.97682, 37.92222, 37.85865, 
    37.78615, 37.7048, 37.61465, 37.5158, 37.40832, 37.2923, 37.16784, 
    37.03504, 36.89401, 36.74487, 36.58773, 36.42271, 36.24994, 36.06956, 
    35.8817, 35.68649, 35.48409, 35.27462, 35.05824, 34.83509, 34.60533, 
    34.36911, 34.12658, 33.87788, 33.62318, 33.36263, 33.09637, 32.82457, 
    32.54737, 32.26494, 31.97741, 31.68493, 31.38766, 31.08575, 30.77932, 
    30.46854, 30.15354, 29.83445, 29.51142, 29.18457,
  29.92181, 30.25368, 30.58158, 30.90537, 31.22494, 31.54013, 31.8508, 
    32.15683, 32.45805, 32.75434, 33.04553, 33.33149, 33.61207, 33.88711, 
    34.15647, 34.42, 34.67754, 34.92895, 35.17407, 35.41275, 35.64485, 
    35.87022, 36.08871, 36.30017, 36.50447, 36.70145, 36.891, 37.07295, 
    37.2472, 37.4136, 37.57203, 37.72238, 37.86452, 37.99836, 38.12377, 
    38.24066, 38.34894, 38.44851, 38.53931, 38.62124, 38.69425, 38.75827, 
    38.81324, 38.85912, 38.89588, 38.92347, 38.94188, 38.95109, 38.95109, 
    38.94188, 38.92347, 38.89588, 38.85912, 38.81324, 38.75827, 38.69425, 
    38.62124, 38.53931, 38.44851, 38.34894, 38.24066, 38.12377, 37.99836, 
    37.86452, 37.72238, 37.57203, 37.4136, 37.2472, 37.07295, 36.891, 
    36.70145, 36.50447, 36.30017, 36.08871, 35.87022, 35.64485, 35.41275, 
    35.17407, 34.92895, 34.67754, 34.42, 34.15647, 33.88711, 33.61207, 
    33.33149, 33.04553, 32.75434, 32.45805, 32.15683, 31.8508, 31.54013, 
    31.22494, 30.90537, 30.58158, 30.25368, 29.92181,
  30.65893, 30.9956, 31.32814, 31.65643, 31.98032, 32.29969, 32.6144, 
    32.9243, 33.22925, 33.52912, 33.82376, 34.11302, 34.39675, 34.67482, 
    34.94707, 35.21335, 35.47353, 35.72744, 35.97494, 36.21589, 36.45013, 
    36.67753, 36.89794, 37.11122, 37.31722, 37.51582, 37.70687, 37.89024, 
    38.06581, 38.23346, 38.39304, 38.54446, 38.6876, 38.82234, 38.94859, 
    39.06625, 39.17523, 39.27544, 39.3668, 39.44924, 39.52269, 39.58709, 
    39.6424, 39.68855, 39.72552, 39.75327, 39.77179, 39.78105, 39.78105, 
    39.77179, 39.75327, 39.72552, 39.68855, 39.6424, 39.58709, 39.52269, 
    39.44924, 39.3668, 39.27544, 39.17523, 39.06625, 38.94859, 38.82234, 
    38.6876, 38.54446, 38.39304, 38.23346, 38.06581, 37.89024, 37.70687, 
    37.51582, 37.31722, 37.11122, 36.89794, 36.67753, 36.45013, 36.21589, 
    35.97494, 35.72744, 35.47353, 35.21335, 34.94707, 34.67482, 34.39675, 
    34.11302, 33.82376, 33.52912, 33.22925, 32.9243, 32.6144, 32.29969, 
    31.98032, 31.65643, 31.32814, 30.9956, 30.65893,
  31.39594, 31.73718, 32.07414, 32.40669, 32.73469, 33.05801, 33.37651, 
    33.69006, 33.99852, 34.30174, 34.59959, 34.89193, 35.1786, 35.45947, 
    35.73439, 36.00322, 36.26581, 36.52202, 36.7717, 37.01471, 37.2509, 
    37.48015, 37.70229, 37.9172, 38.12474, 38.32478, 38.51718, 38.70182, 
    38.87856, 39.04729, 39.20789, 39.36025, 39.50425, 39.63979, 39.76678, 
    39.88511, 39.99469, 40.09544, 40.18729, 40.27016, 40.34399, 40.40873, 
    40.46431, 40.51069, 40.54784, 40.57574, 40.59435, 40.60365, 40.60365, 
    40.59435, 40.57574, 40.54784, 40.51069, 40.46431, 40.40873, 40.34399, 
    40.27016, 40.18729, 40.09544, 39.99469, 39.88511, 39.76678, 39.63979, 
    39.50425, 39.36025, 39.20789, 39.04729, 38.87856, 38.70182, 38.51718, 
    38.32478, 38.12474, 37.9172, 37.70229, 37.48015, 37.2509, 37.01471, 
    36.7717, 36.52202, 36.26581, 36.00322, 35.73439, 35.45947, 35.1786, 
    34.89193, 34.59959, 34.30174, 33.99852, 33.69006, 33.37651, 33.05801, 
    32.73469, 32.40669, 32.07414, 31.73718, 31.39594,
  32.13284, 32.47842, 32.81957, 33.15614, 33.48802, 33.81506, 34.13713, 
    34.4541, 34.76583, 35.07218, 35.37302, 35.66821, 35.9576, 36.24105, 
    36.51843, 36.78959, 37.05439, 37.31269, 37.56434, 37.80922, 38.04717, 
    38.27806, 38.50176, 38.71813, 38.92703, 39.12834, 39.32193, 39.50767, 
    39.68544, 39.85512, 40.0166, 40.16977, 40.31451, 40.45074, 40.57834, 
    40.69724, 40.80733, 40.90854, 41.0008, 41.08404, 41.15818, 41.22319, 
    41.279, 41.32558, 41.36288, 41.39089, 41.40957, 41.41891, 41.41891, 
    41.40957, 41.39089, 41.36288, 41.32558, 41.279, 41.22319, 41.15818, 
    41.08404, 41.0008, 40.90854, 40.80733, 40.69724, 40.57834, 40.45074, 
    40.31451, 40.16977, 40.0166, 39.85512, 39.68544, 39.50767, 39.32193, 
    39.12834, 38.92703, 38.71813, 38.50176, 38.27806, 38.04717, 37.80922, 
    37.56434, 37.31269, 37.05439, 36.78959, 36.51843, 36.24105, 35.9576, 
    35.66821, 35.37302, 35.07218, 34.76583, 34.4541, 34.13713, 33.81506, 
    33.48802, 33.15614, 32.81957, 32.47842, 32.13284,
  32.86962, 33.21932, 33.56442, 33.90479, 34.2403, 34.57083, 34.89624, 
    35.2164, 35.53117, 35.84042, 36.14403, 36.44184, 36.73372, 37.01954, 
    37.29916, 37.57244, 37.83924, 38.09942, 38.35286, 38.5994, 38.83891, 
    39.07127, 39.29634, 39.51399, 39.72409, 39.9265, 40.12112, 40.30781, 
    40.48646, 40.65696, 40.81918, 40.97303, 41.1184, 41.25519, 41.38331, 
    41.50267, 41.61318, 41.71477, 41.80736, 41.89089, 41.96529, 42.03052, 
    42.08652, 42.13324, 42.17067, 42.19876, 42.2175, 42.22688, 42.22688, 
    42.2175, 42.19876, 42.17067, 42.13324, 42.08652, 42.03052, 41.96529, 
    41.89089, 41.80736, 41.71477, 41.61318, 41.50267, 41.38331, 41.25519, 
    41.1184, 40.97303, 40.81918, 40.65696, 40.48646, 40.30781, 40.12112, 
    39.9265, 39.72409, 39.51399, 39.29634, 39.07127, 38.83891, 38.5994, 
    38.35286, 38.09942, 37.83924, 37.57244, 37.29916, 37.01954, 36.73372, 
    36.44184, 36.14403, 35.84042, 35.53117, 35.2164, 34.89624, 34.57083, 
    34.2403, 33.90479, 33.56442, 33.21932, 32.86962,
  33.60628, 33.95987, 34.30869, 34.65261, 34.99154, 35.32531, 35.65382, 
    35.97694, 36.29453, 36.60646, 36.91259, 37.21281, 37.50697, 37.79493, 
    38.07658, 38.35176, 38.62035, 38.88222, 39.13723, 39.38524, 39.62614, 
    39.85978, 40.08604, 40.30479, 40.51591, 40.71927, 40.91476, 41.10225, 
    41.28164, 41.4528, 41.61564, 41.77005, 41.91592, 42.05317, 42.18171, 
    42.30143, 42.41228, 42.51416, 42.60701, 42.69076, 42.76536, 42.83075, 
    42.88689, 42.93373, 42.97124, 42.9994, 43.01819, 43.02758, 43.02758, 
    43.01819, 42.9994, 42.97124, 42.93373, 42.88689, 42.83075, 42.76536, 
    42.69076, 42.60701, 42.51416, 42.41228, 42.30143, 42.18171, 42.05317, 
    41.91592, 41.77005, 41.61564, 41.4528, 41.28164, 41.10225, 40.91476, 
    40.71927, 40.51591, 40.30479, 40.08604, 39.85978, 39.62614, 39.38524, 
    39.13723, 38.88222, 38.62035, 38.35176, 38.07658, 37.79493, 37.50697, 
    37.21281, 36.91259, 36.60646, 36.29453, 35.97694, 35.65382, 35.32531, 
    34.99154, 34.65261, 34.30869, 33.95987, 33.60628,
  34.34282, 34.70005, 35.05236, 35.39962, 35.7417, 36.0785, 36.40988, 
    36.73572, 37.05589, 37.37026, 37.67871, 37.9811, 38.27731, 38.56721, 
    38.85067, 39.12755, 39.39772, 39.66107, 39.91746, 40.16676, 40.40884, 
    40.64358, 40.87085, 41.09053, 41.30251, 41.50666, 41.70287, 41.89101, 
    42.07099, 42.24269, 42.40602, 42.56086, 42.70713, 42.84472, 42.97356, 
    43.09357, 43.20465, 43.30674, 43.39978, 43.48369, 43.55843, 43.62393, 
    43.68016, 43.72708, 43.76466, 43.79286, 43.81168, 43.82109, 43.82109, 
    43.81168, 43.79286, 43.76466, 43.72708, 43.68016, 43.62393, 43.55843, 
    43.48369, 43.39978, 43.30674, 43.20465, 43.09357, 42.97356, 42.84472, 
    42.70713, 42.56086, 42.40602, 42.24269, 42.07099, 41.89101, 41.70287, 
    41.50666, 41.30251, 41.09053, 40.87085, 40.64358, 40.40884, 40.16676, 
    39.91746, 39.66107, 39.39772, 39.12755, 38.85067, 38.56721, 38.27731, 
    37.9811, 37.67871, 37.37026, 37.05589, 36.73572, 36.40988, 36.0785, 
    35.7417, 35.39962, 35.05236, 34.70005, 34.34282,
  35.07925, 35.43988, 35.79544, 36.14578, 36.4908, 36.83038, 37.1644, 
    37.49273, 37.81525, 38.13184, 38.44237, 38.74672, 39.04476, 39.33637, 
    39.62142, 39.89979, 40.17135, 40.43598, 40.69355, 40.94394, 41.18702, 
    41.42268, 41.65079, 41.87124, 42.08391, 42.28868, 42.48545, 42.67411, 
    42.85454, 43.02665, 43.19033, 43.34549, 43.49203, 43.62987, 43.75893, 
    43.87911, 43.99035, 44.09258, 44.18572, 44.26973, 44.34454, 44.41011, 
    44.46639, 44.51335, 44.55096, 44.57919, 44.59801, 44.60743, 44.60743, 
    44.59801, 44.57919, 44.55096, 44.51335, 44.46639, 44.41011, 44.34454, 
    44.26973, 44.18572, 44.09258, 43.99035, 43.87911, 43.75893, 43.62987, 
    43.49203, 43.34549, 43.19033, 43.02665, 42.85454, 42.67411, 42.48545, 
    42.28868, 42.08391, 41.87124, 41.65079, 41.42268, 41.18702, 40.94394, 
    40.69355, 40.43598, 40.17135, 39.89979, 39.62142, 39.33637, 39.04476, 
    38.74672, 38.44237, 38.13184, 37.81525, 37.49273, 37.1644, 36.83038, 
    36.4908, 36.14578, 35.79544, 35.43988, 35.07925 ;

 area =
  5.832426e+09, 5.885548e+09, 5.937712e+09, 5.988909e+09, 6.039129e+09, 
    6.088361e+09, 6.136596e+09, 6.183825e+09, 6.230037e+09, 6.275223e+09, 
    6.319373e+09, 6.362479e+09, 6.404531e+09, 6.445522e+09, 6.485442e+09, 
    6.524282e+09, 6.562035e+09, 6.598693e+09, 6.634248e+09, 6.668692e+09, 
    6.702019e+09, 6.734221e+09, 6.76529e+09, 6.795221e+09, 6.824007e+09, 
    6.851641e+09, 6.878117e+09, 6.903431e+09, 6.927576e+09, 6.950547e+09, 
    6.972339e+09, 6.992947e+09, 7.012366e+09, 7.030593e+09, 7.047623e+09, 
    7.063453e+09, 7.078078e+09, 7.091497e+09, 7.103705e+09, 7.1147e+09, 
    7.124479e+09, 7.133041e+09, 7.140384e+09, 7.146505e+09, 7.151404e+09, 
    7.155078e+09, 7.157529e+09, 7.158754e+09, 7.158754e+09, 7.157529e+09, 
    7.155078e+09, 7.151404e+09, 7.146505e+09, 7.140384e+09, 7.133041e+09, 
    7.124479e+09, 7.1147e+09, 7.103705e+09, 7.091497e+09, 7.078078e+09, 
    7.063453e+09, 7.047623e+09, 7.030593e+09, 7.012366e+09, 6.992947e+09, 
    6.972339e+09, 6.950547e+09, 6.927576e+09, 6.903431e+09, 6.878117e+09, 
    6.851641e+09, 6.824007e+09, 6.795221e+09, 6.76529e+09, 6.734221e+09, 
    6.702019e+09, 6.668692e+09, 6.634248e+09, 6.598693e+09, 6.562035e+09, 
    6.524282e+09, 6.485442e+09, 6.445522e+09, 6.404531e+09, 6.362479e+09, 
    6.319373e+09, 6.275223e+09, 6.230037e+09, 6.183825e+09, 6.136596e+09, 
    6.088361e+09, 6.039129e+09, 5.988909e+09, 5.937712e+09, 5.885548e+09, 
    5.832426e+09,
  5.885548e+09, 5.942029e+09, 5.99757e+09, 6.052155e+09, 6.105772e+09, 
    6.158404e+09, 6.210038e+09, 6.260659e+09, 6.310255e+09, 6.35881e+09, 
    6.406312e+09, 6.452746e+09, 6.4981e+09, 6.54236e+09, 6.585513e+09, 
    6.627547e+09, 6.668449e+09, 6.708208e+09, 6.74681e+09, 6.784244e+09, 
    6.8205e+09, 6.855565e+09, 6.889429e+09, 6.922081e+09, 6.953512e+09, 
    6.98371e+09, 7.012667e+09, 7.040374e+09, 7.066821e+09, 7.092e+09, 
    7.115902e+09, 7.138521e+09, 7.159848e+09, 7.179877e+09, 7.198601e+09, 
    7.216014e+09, 7.23211e+09, 7.246883e+09, 7.260329e+09, 7.272444e+09, 
    7.283223e+09, 7.292662e+09, 7.30076e+09, 7.307511e+09, 7.312915e+09, 
    7.316969e+09, 7.319673e+09, 7.321026e+09, 7.321026e+09, 7.319673e+09, 
    7.316969e+09, 7.312915e+09, 7.307511e+09, 7.30076e+09, 7.292662e+09, 
    7.283223e+09, 7.272444e+09, 7.260329e+09, 7.246883e+09, 7.23211e+09, 
    7.216014e+09, 7.198601e+09, 7.179877e+09, 7.159848e+09, 7.138521e+09, 
    7.115902e+09, 7.092e+09, 7.066821e+09, 7.040374e+09, 7.012667e+09, 
    6.98371e+09, 6.953512e+09, 6.922081e+09, 6.889429e+09, 6.855565e+09, 
    6.8205e+09, 6.784244e+09, 6.74681e+09, 6.708208e+09, 6.668449e+09, 
    6.627547e+09, 6.585513e+09, 6.54236e+09, 6.4981e+09, 6.452746e+09, 
    6.406312e+09, 6.35881e+09, 6.310255e+09, 6.260659e+09, 6.210038e+09, 
    6.158404e+09, 6.105772e+09, 6.052155e+09, 5.99757e+09, 5.942029e+09, 
    5.885548e+09,
  5.937712e+09, 5.99757e+09, 6.056508e+09, 6.114508e+09, 6.171552e+09, 
    6.227619e+09, 6.282692e+09, 6.336752e+09, 6.38978e+09, 6.441759e+09, 
    6.492669e+09, 6.542493e+09, 6.591213e+09, 6.638811e+09, 6.685269e+09, 
    6.730571e+09, 6.774699e+09, 6.817636e+09, 6.859367e+09, 6.899874e+09, 
    6.939143e+09, 6.977157e+09, 7.013901e+09, 7.049361e+09, 7.083523e+09, 
    7.116371e+09, 7.147894e+09, 7.178077e+09, 7.206909e+09, 7.234377e+09, 
    7.260469e+09, 7.285175e+09, 7.308484e+09, 7.330385e+09, 7.350871e+09, 
    7.36993e+09, 7.387556e+09, 7.403741e+09, 7.418477e+09, 7.431758e+09, 
    7.443579e+09, 7.453934e+09, 7.462817e+09, 7.470226e+09, 7.476158e+09, 
    7.480609e+09, 7.483577e+09, 7.485062e+09, 7.485062e+09, 7.483577e+09, 
    7.480609e+09, 7.476158e+09, 7.470226e+09, 7.462817e+09, 7.453934e+09, 
    7.443579e+09, 7.431758e+09, 7.418477e+09, 7.403741e+09, 7.387556e+09, 
    7.36993e+09, 7.350871e+09, 7.330385e+09, 7.308484e+09, 7.285175e+09, 
    7.260469e+09, 7.234377e+09, 7.206909e+09, 7.178077e+09, 7.147894e+09, 
    7.116371e+09, 7.083523e+09, 7.049361e+09, 7.013901e+09, 6.977157e+09, 
    6.939143e+09, 6.899874e+09, 6.859367e+09, 6.817636e+09, 6.774699e+09, 
    6.730571e+09, 6.685269e+09, 6.638811e+09, 6.591213e+09, 6.542493e+09, 
    6.492669e+09, 6.441759e+09, 6.38978e+09, 6.336752e+09, 6.282692e+09, 
    6.227619e+09, 6.171552e+09, 6.114508e+09, 6.056508e+09, 5.99757e+09, 
    5.937712e+09,
  5.988909e+09, 6.052155e+09, 6.114508e+09, 6.175945e+09, 6.236442e+09, 
    6.295976e+09, 6.354524e+09, 6.412062e+09, 6.468569e+09, 6.52402e+09, 
    6.578392e+09, 6.631664e+09, 6.683811e+09, 6.734811e+09, 6.784643e+09, 
    6.833284e+09, 6.880711e+09, 6.926904e+09, 6.971842e+09, 7.015503e+09, 
    7.057866e+09, 7.098912e+09, 7.13862e+09, 7.176973e+09, 7.21395e+09, 
    7.249533e+09, 7.283705e+09, 7.316448e+09, 7.347746e+09, 7.377583e+09, 
    7.405943e+09, 7.432813e+09, 7.458176e+09, 7.482021e+09, 7.504335e+09, 
    7.525106e+09, 7.544322e+09, 7.561974e+09, 7.578052e+09, 7.592547e+09, 
    7.605452e+09, 7.616759e+09, 7.626462e+09, 7.634556e+09, 7.641037e+09, 
    7.645901e+09, 7.649145e+09, 7.650767e+09, 7.650767e+09, 7.649145e+09, 
    7.645901e+09, 7.641037e+09, 7.634556e+09, 7.626462e+09, 7.616759e+09, 
    7.605452e+09, 7.592547e+09, 7.578052e+09, 7.561974e+09, 7.544322e+09, 
    7.525106e+09, 7.504335e+09, 7.482021e+09, 7.458176e+09, 7.432813e+09, 
    7.405943e+09, 7.377583e+09, 7.347746e+09, 7.316448e+09, 7.283705e+09, 
    7.249533e+09, 7.21395e+09, 7.176973e+09, 7.13862e+09, 7.098912e+09, 
    7.057866e+09, 7.015503e+09, 6.971842e+09, 6.926904e+09, 6.880711e+09, 
    6.833284e+09, 6.784643e+09, 6.734811e+09, 6.683811e+09, 6.631664e+09, 
    6.578392e+09, 6.52402e+09, 6.468569e+09, 6.412062e+09, 6.354524e+09, 
    6.295976e+09, 6.236442e+09, 6.175945e+09, 6.114508e+09, 6.052155e+09, 
    5.988909e+09,
  6.039129e+09, 6.105772e+09, 6.171552e+09, 6.236442e+09, 6.300414e+09, 
    6.363442e+09, 6.425497e+09, 6.486551e+09, 6.546576e+09, 6.605544e+09, 
    6.663429e+09, 6.720201e+09, 6.775833e+09, 6.830297e+09, 6.883567e+09, 
    6.935614e+09, 6.986412e+09, 7.035934e+09, 7.084154e+09, 7.131045e+09, 
    7.176583e+09, 7.220742e+09, 7.263496e+09, 7.304823e+09, 7.344698e+09, 
    7.383099e+09, 7.420003e+09, 7.455388e+09, 7.489233e+09, 7.521518e+09, 
    7.552224e+09, 7.581331e+09, 7.608822e+09, 7.634681e+09, 7.65889e+09, 
    7.681435e+09, 7.702302e+09, 7.721477e+09, 7.738948e+09, 7.754704e+09, 
    7.768736e+09, 7.781033e+09, 7.791588e+09, 7.800395e+09, 7.807448e+09, 
    7.812741e+09, 7.816271e+09, 7.818037e+09, 7.818037e+09, 7.816271e+09, 
    7.812741e+09, 7.807448e+09, 7.800395e+09, 7.791588e+09, 7.781033e+09, 
    7.768736e+09, 7.754704e+09, 7.738948e+09, 7.721477e+09, 7.702302e+09, 
    7.681435e+09, 7.65889e+09, 7.634681e+09, 7.608822e+09, 7.581331e+09, 
    7.552224e+09, 7.521518e+09, 7.489233e+09, 7.455388e+09, 7.420003e+09, 
    7.383099e+09, 7.344698e+09, 7.304823e+09, 7.263496e+09, 7.220742e+09, 
    7.176583e+09, 7.131045e+09, 7.084154e+09, 7.035934e+09, 6.986412e+09, 
    6.935614e+09, 6.883567e+09, 6.830297e+09, 6.775833e+09, 6.720201e+09, 
    6.663429e+09, 6.605544e+09, 6.546576e+09, 6.486551e+09, 6.425497e+09, 
    6.363442e+09, 6.300414e+09, 6.236442e+09, 6.171552e+09, 6.105772e+09, 
    6.039129e+09,
  6.088361e+09, 6.158404e+09, 6.227619e+09, 6.295976e+09, 6.363442e+09, 
    6.429985e+09, 6.495574e+09, 6.560175e+09, 6.623755e+09, 6.686283e+09, 
    6.747724e+09, 6.808046e+09, 6.867216e+09, 6.925201e+09, 6.981969e+09, 
    7.037487e+09, 7.091722e+09, 7.144643e+09, 7.196217e+09, 7.246414e+09, 
    7.295202e+09, 7.342552e+09, 7.388432e+09, 7.432814e+09, 7.475667e+09, 
    7.516966e+09, 7.556683e+09, 7.594789e+09, 7.631261e+09, 7.666072e+09, 
    7.699199e+09, 7.73062e+09, 7.760311e+09, 7.788252e+09, 7.814423e+09, 
    7.838806e+09, 7.861382e+09, 7.882135e+09, 7.901051e+09, 7.918115e+09, 
    7.933316e+09, 7.946641e+09, 7.958081e+09, 7.967627e+09, 7.975273e+09, 
    7.981012e+09, 7.984841e+09, 7.986756e+09, 7.986756e+09, 7.984841e+09, 
    7.981012e+09, 7.975273e+09, 7.967627e+09, 7.958081e+09, 7.946641e+09, 
    7.933316e+09, 7.918115e+09, 7.901051e+09, 7.882135e+09, 7.861382e+09, 
    7.838806e+09, 7.814423e+09, 7.788252e+09, 7.760311e+09, 7.73062e+09, 
    7.699199e+09, 7.666072e+09, 7.631261e+09, 7.594789e+09, 7.556683e+09, 
    7.516966e+09, 7.475667e+09, 7.432814e+09, 7.388432e+09, 7.342552e+09, 
    7.295202e+09, 7.246414e+09, 7.196217e+09, 7.144643e+09, 7.091722e+09, 
    7.037487e+09, 6.981969e+09, 6.925201e+09, 6.867216e+09, 6.808046e+09, 
    6.747724e+09, 6.686283e+09, 6.623755e+09, 6.560175e+09, 6.495574e+09, 
    6.429985e+09, 6.363442e+09, 6.295976e+09, 6.227619e+09, 6.158404e+09, 
    6.088361e+09,
  6.136596e+09, 6.210038e+09, 6.282692e+09, 6.354524e+09, 6.425497e+09, 
    6.495574e+09, 6.564719e+09, 6.632894e+09, 6.700061e+09, 6.766183e+09, 
    6.831222e+09, 6.895139e+09, 6.957896e+09, 7.019455e+09, 7.079777e+09, 
    7.138825e+09, 7.196561e+09, 7.252946e+09, 7.307944e+09, 7.361518e+09, 
    7.41363e+09, 7.464245e+09, 7.513327e+09, 7.56084e+09, 7.606751e+09, 
    7.651027e+09, 7.693634e+09, 7.734541e+09, 7.773715e+09, 7.811129e+09, 
    7.846753e+09, 7.880559e+09, 7.912521e+09, 7.942612e+09, 7.970811e+09, 
    7.997093e+09, 8.021437e+09, 8.043825e+09, 8.064236e+09, 8.082655e+09, 
    8.099066e+09, 8.113456e+09, 8.125813e+09, 8.136126e+09, 8.144387e+09, 
    8.150589e+09, 8.154726e+09, 8.156796e+09, 8.156796e+09, 8.154726e+09, 
    8.150589e+09, 8.144387e+09, 8.136126e+09, 8.125813e+09, 8.113456e+09, 
    8.099066e+09, 8.082655e+09, 8.064236e+09, 8.043825e+09, 8.021437e+09, 
    7.997093e+09, 7.970811e+09, 7.942612e+09, 7.912521e+09, 7.880559e+09, 
    7.846753e+09, 7.811129e+09, 7.773715e+09, 7.734541e+09, 7.693634e+09, 
    7.651027e+09, 7.606751e+09, 7.56084e+09, 7.513327e+09, 7.464245e+09, 
    7.41363e+09, 7.361518e+09, 7.307944e+09, 7.252946e+09, 7.196561e+09, 
    7.138825e+09, 7.079777e+09, 7.019455e+09, 6.957896e+09, 6.895139e+09, 
    6.831222e+09, 6.766183e+09, 6.700061e+09, 6.632894e+09, 6.564719e+09, 
    6.495574e+09, 6.425497e+09, 6.354524e+09, 6.282692e+09, 6.210038e+09, 
    6.136596e+09,
  6.183825e+09, 6.260659e+09, 6.336752e+09, 6.412062e+09, 6.486551e+09, 
    6.560175e+09, 6.632894e+09, 6.704666e+09, 6.775447e+09, 6.845195e+09, 
    6.913867e+09, 6.981418e+09, 7.047806e+09, 7.112987e+09, 7.176916e+09, 
    7.23955e+09, 7.300845e+09, 7.360757e+09, 7.419243e+09, 7.47626e+09, 
    7.531766e+09, 7.585717e+09, 7.638074e+09, 7.688794e+09, 7.737838e+09, 
    7.785166e+09, 7.830739e+09, 7.874522e+09, 7.916475e+09, 7.956566e+09, 
    7.994759e+09, 8.031022e+09, 8.065324e+09, 8.097633e+09, 8.127923e+09, 
    8.156166e+09, 8.182336e+09, 8.20641e+09, 8.228367e+09, 8.248187e+09, 
    8.26585e+09, 8.281342e+09, 8.294647e+09, 8.305754e+09, 8.314652e+09, 
    8.321333e+09, 8.32579e+09, 8.32802e+09, 8.32802e+09, 8.32579e+09, 
    8.321333e+09, 8.314652e+09, 8.305754e+09, 8.294647e+09, 8.281342e+09, 
    8.26585e+09, 8.248187e+09, 8.228367e+09, 8.20641e+09, 8.182336e+09, 
    8.156166e+09, 8.127923e+09, 8.097633e+09, 8.065324e+09, 8.031022e+09, 
    7.994759e+09, 7.956566e+09, 7.916475e+09, 7.874522e+09, 7.830739e+09, 
    7.785166e+09, 7.737838e+09, 7.688794e+09, 7.638074e+09, 7.585717e+09, 
    7.531766e+09, 7.47626e+09, 7.419243e+09, 7.360757e+09, 7.300845e+09, 
    7.23955e+09, 7.176916e+09, 7.112987e+09, 7.047806e+09, 6.981418e+09, 
    6.913867e+09, 6.845195e+09, 6.775447e+09, 6.704666e+09, 6.632894e+09, 
    6.560175e+09, 6.486551e+09, 6.412062e+09, 6.336752e+09, 6.260659e+09, 
    6.183825e+09,
  6.230037e+09, 6.310255e+09, 6.38978e+09, 6.468569e+09, 6.546576e+09, 
    6.623755e+09, 6.700061e+09, 6.775447e+09, 6.849864e+09, 6.923265e+09, 
    6.9956e+09, 7.066822e+09, 7.136881e+09, 7.205726e+09, 7.273309e+09, 
    7.339579e+09, 7.404488e+09, 7.467984e+09, 7.530018e+09, 7.590542e+09, 
    7.649507e+09, 7.706863e+09, 7.762563e+09, 7.816561e+09, 7.868808e+09, 
    7.919261e+09, 7.967875e+09, 8.014606e+09, 8.059411e+09, 8.10225e+09, 
    8.143084e+09, 8.181873e+09, 8.218582e+09, 8.253174e+09, 8.285618e+09, 
    8.31588e+09, 8.343933e+09, 8.369748e+09, 8.3933e+09, 8.414565e+09, 
    8.433522e+09, 8.450151e+09, 8.464436e+09, 8.476363e+09, 8.485919e+09, 
    8.493095e+09, 8.497883e+09, 8.500278e+09, 8.500278e+09, 8.497883e+09, 
    8.493095e+09, 8.485919e+09, 8.476363e+09, 8.464436e+09, 8.450151e+09, 
    8.433522e+09, 8.414565e+09, 8.3933e+09, 8.369748e+09, 8.343933e+09, 
    8.31588e+09, 8.285618e+09, 8.253174e+09, 8.218582e+09, 8.181873e+09, 
    8.143084e+09, 8.10225e+09, 8.059411e+09, 8.014606e+09, 7.967875e+09, 
    7.919261e+09, 7.868808e+09, 7.816561e+09, 7.762563e+09, 7.706863e+09, 
    7.649507e+09, 7.590542e+09, 7.530018e+09, 7.467984e+09, 7.404488e+09, 
    7.339579e+09, 7.273309e+09, 7.205726e+09, 7.136881e+09, 7.066822e+09, 
    6.9956e+09, 6.923265e+09, 6.849864e+09, 6.775447e+09, 6.700061e+09, 
    6.623755e+09, 6.546576e+09, 6.468569e+09, 6.38978e+09, 6.310255e+09, 
    6.230037e+09,
  6.275223e+09, 6.35881e+09, 6.441759e+09, 6.52402e+09, 6.605544e+09, 
    6.686283e+09, 6.766183e+09, 6.845195e+09, 6.923265e+09, 7.000339e+09, 
    7.076365e+09, 7.151286e+09, 7.225049e+09, 7.297597e+09, 7.368877e+09, 
    7.438829e+09, 7.5074e+09, 7.574533e+09, 7.640172e+09, 7.704261e+09, 
    7.766745e+09, 7.827569e+09, 7.886679e+09, 7.94402e+09, 7.99954e+09, 
    8.053188e+09, 8.10491e+09, 8.15466e+09, 8.202386e+09, 8.248043e+09, 
    8.291585e+09, 8.332967e+09, 8.372148e+09, 8.409087e+09, 8.443745e+09, 
    8.476086e+09, 8.506077e+09, 8.533684e+09, 8.558878e+09, 8.581632e+09, 
    8.601922e+09, 8.619724e+09, 8.63502e+09, 8.647793e+09, 8.658028e+09, 
    8.665715e+09, 8.670843e+09, 8.673409e+09, 8.673409e+09, 8.670843e+09, 
    8.665715e+09, 8.658028e+09, 8.647793e+09, 8.63502e+09, 8.619724e+09, 
    8.601922e+09, 8.581632e+09, 8.558878e+09, 8.533684e+09, 8.506077e+09, 
    8.476086e+09, 8.443745e+09, 8.409087e+09, 8.372148e+09, 8.332967e+09, 
    8.291585e+09, 8.248043e+09, 8.202386e+09, 8.15466e+09, 8.10491e+09, 
    8.053188e+09, 7.99954e+09, 7.94402e+09, 7.886679e+09, 7.827569e+09, 
    7.766745e+09, 7.704261e+09, 7.640172e+09, 7.574533e+09, 7.5074e+09, 
    7.438829e+09, 7.368877e+09, 7.297597e+09, 7.225049e+09, 7.151286e+09, 
    7.076365e+09, 7.000339e+09, 6.923265e+09, 6.845195e+09, 6.766183e+09, 
    6.686283e+09, 6.605544e+09, 6.52402e+09, 6.441759e+09, 6.35881e+09, 
    6.275223e+09,
  6.319373e+09, 6.406312e+09, 6.492669e+09, 6.578392e+09, 6.663429e+09, 
    6.747724e+09, 6.831222e+09, 6.913867e+09, 6.9956e+09, 7.076365e+09, 
    7.1561e+09, 7.234745e+09, 7.312241e+09, 7.388526e+09, 7.463537e+09, 
    7.537212e+09, 7.60949e+09, 7.680307e+09, 7.749601e+09, 7.817309e+09, 
    7.883369e+09, 7.94772e+09, 8.010299e+09, 8.071048e+09, 8.129904e+09, 
    8.186811e+09, 8.241709e+09, 8.294543e+09, 8.345257e+09, 8.393798e+09, 
    8.440113e+09, 8.484152e+09, 8.525868e+09, 8.565214e+09, 8.602145e+09, 
    8.636621e+09, 8.668601e+09, 8.698051e+09, 8.724934e+09, 8.749221e+09, 
    8.770882e+09, 8.789891e+09, 8.806228e+09, 8.819871e+09, 8.830806e+09, 
    8.839017e+09, 8.844498e+09, 8.84724e+09, 8.84724e+09, 8.844498e+09, 
    8.839017e+09, 8.830806e+09, 8.819871e+09, 8.806228e+09, 8.789891e+09, 
    8.770882e+09, 8.749221e+09, 8.724934e+09, 8.698051e+09, 8.668601e+09, 
    8.636621e+09, 8.602145e+09, 8.565214e+09, 8.525868e+09, 8.484152e+09, 
    8.440113e+09, 8.393798e+09, 8.345257e+09, 8.294543e+09, 8.241709e+09, 
    8.186811e+09, 8.129904e+09, 8.071048e+09, 8.010299e+09, 7.94772e+09, 
    7.883369e+09, 7.817309e+09, 7.749601e+09, 7.680307e+09, 7.60949e+09, 
    7.537212e+09, 7.463537e+09, 7.388526e+09, 7.312241e+09, 7.234745e+09, 
    7.1561e+09, 7.076365e+09, 6.9956e+09, 6.913867e+09, 6.831222e+09, 
    6.747724e+09, 6.663429e+09, 6.578392e+09, 6.492669e+09, 6.406312e+09, 
    6.319373e+09,
  6.362479e+09, 6.452746e+09, 6.542493e+09, 6.631664e+09, 6.720201e+09, 
    6.808046e+09, 6.895139e+09, 6.981418e+09, 7.066822e+09, 7.151286e+09, 
    7.234745e+09, 7.317134e+09, 7.398386e+09, 7.478433e+09, 7.557208e+09, 
    7.634641e+09, 7.710664e+09, 7.785207e+09, 7.858201e+09, 7.929576e+09, 
    7.999264e+09, 8.067195e+09, 8.133301e+09, 8.197513e+09, 8.259766e+09, 
    8.319992e+09, 8.378128e+09, 8.434108e+09, 8.487873e+09, 8.539359e+09, 
    8.58851e+09, 8.635267e+09, 8.679578e+09, 8.721389e+09, 8.760649e+09, 
    8.797313e+09, 8.831335e+09, 8.862674e+09, 8.891291e+09, 8.917151e+09, 
    8.940219e+09, 8.96047e+09, 8.977876e+09, 8.992415e+09, 9.004068e+09, 
    9.012821e+09, 9.018663e+09, 9.021585e+09, 9.021585e+09, 9.018663e+09, 
    9.012821e+09, 9.004068e+09, 8.992415e+09, 8.977876e+09, 8.96047e+09, 
    8.940219e+09, 8.917151e+09, 8.891291e+09, 8.862674e+09, 8.831335e+09, 
    8.797313e+09, 8.760649e+09, 8.721389e+09, 8.679578e+09, 8.635267e+09, 
    8.58851e+09, 8.539359e+09, 8.487873e+09, 8.434108e+09, 8.378128e+09, 
    8.319992e+09, 8.259766e+09, 8.197513e+09, 8.133301e+09, 8.067195e+09, 
    7.999264e+09, 7.929576e+09, 7.858201e+09, 7.785207e+09, 7.710664e+09, 
    7.634641e+09, 7.557208e+09, 7.478433e+09, 7.398386e+09, 7.317134e+09, 
    7.234745e+09, 7.151286e+09, 7.066822e+09, 6.981418e+09, 6.895139e+09, 
    6.808046e+09, 6.720201e+09, 6.631664e+09, 6.542493e+09, 6.452746e+09, 
    6.362479e+09,
  6.404531e+09, 6.4981e+09, 6.591213e+09, 6.683811e+09, 6.775833e+09, 
    6.867216e+09, 6.957896e+09, 7.047806e+09, 7.136881e+09, 7.225049e+09, 
    7.312241e+09, 7.398386e+09, 7.483411e+09, 7.567242e+09, 7.649805e+09, 
    7.731025e+09, 7.810825e+09, 7.889131e+09, 7.965864e+09, 8.04095e+09, 
    8.11431e+09, 8.18587e+09, 8.255552e+09, 8.323282e+09, 8.388985e+09, 
    8.452588e+09, 8.514017e+09, 8.573202e+09, 8.630074e+09, 8.684566e+09, 
    8.736609e+09, 8.786142e+09, 8.833104e+09, 8.877434e+09, 8.919077e+09, 
    8.95798e+09, 8.994092e+09, 9.027367e+09, 9.05776e+09, 9.085231e+09, 
    9.109745e+09, 9.131267e+09, 9.14977e+09, 9.165227e+09, 9.177618e+09, 
    9.186927e+09, 9.193139e+09, 9.196247e+09, 9.196247e+09, 9.193139e+09, 
    9.186927e+09, 9.177618e+09, 9.165227e+09, 9.14977e+09, 9.131267e+09, 
    9.109745e+09, 9.085231e+09, 9.05776e+09, 9.027367e+09, 8.994092e+09, 
    8.95798e+09, 8.919077e+09, 8.877434e+09, 8.833104e+09, 8.786142e+09, 
    8.736609e+09, 8.684566e+09, 8.630074e+09, 8.573202e+09, 8.514017e+09, 
    8.452588e+09, 8.388985e+09, 8.323282e+09, 8.255552e+09, 8.18587e+09, 
    8.11431e+09, 8.04095e+09, 7.965864e+09, 7.889131e+09, 7.810825e+09, 
    7.731025e+09, 7.649805e+09, 7.567242e+09, 7.483411e+09, 7.398386e+09, 
    7.312241e+09, 7.225049e+09, 7.136881e+09, 7.047806e+09, 6.957896e+09, 
    6.867216e+09, 6.775833e+09, 6.683811e+09, 6.591213e+09, 6.4981e+09, 
    6.404531e+09,
  6.445522e+09, 6.54236e+09, 6.638811e+09, 6.734811e+09, 6.830297e+09, 
    6.925201e+09, 7.019455e+09, 7.112987e+09, 7.205726e+09, 7.297597e+09, 
    7.388526e+09, 7.478433e+09, 7.567242e+09, 7.654872e+09, 7.741242e+09, 
    7.826271e+09, 7.909876e+09, 7.991974e+09, 8.072481e+09, 8.151313e+09, 
    8.228386e+09, 8.303616e+09, 8.37692e+09, 8.448214e+09, 8.517416e+09, 
    8.584445e+09, 8.649221e+09, 8.711665e+09, 8.771699e+09, 8.829247e+09, 
    8.884238e+09, 8.936601e+09, 8.986266e+09, 9.033167e+09, 9.077242e+09, 
    9.118431e+09, 9.156679e+09, 9.191932e+09, 9.224142e+09, 9.253263e+09, 
    9.279254e+09, 9.302078e+09, 9.321703e+09, 9.338102e+09, 9.351248e+09, 
    9.361125e+09, 9.367718e+09, 9.371016e+09, 9.371016e+09, 9.367718e+09, 
    9.361125e+09, 9.351248e+09, 9.338102e+09, 9.321703e+09, 9.302078e+09, 
    9.279254e+09, 9.253263e+09, 9.224142e+09, 9.191932e+09, 9.156679e+09, 
    9.118431e+09, 9.077242e+09, 9.033167e+09, 8.986266e+09, 8.936601e+09, 
    8.884238e+09, 8.829247e+09, 8.771699e+09, 8.711665e+09, 8.649221e+09, 
    8.584445e+09, 8.517416e+09, 8.448214e+09, 8.37692e+09, 8.303616e+09, 
    8.228386e+09, 8.151313e+09, 8.072481e+09, 7.991974e+09, 7.909876e+09, 
    7.826271e+09, 7.741242e+09, 7.654872e+09, 7.567242e+09, 7.478433e+09, 
    7.388526e+09, 7.297597e+09, 7.205726e+09, 7.112987e+09, 7.019455e+09, 
    6.925201e+09, 6.830297e+09, 6.734811e+09, 6.638811e+09, 6.54236e+09, 
    6.445522e+09,
  6.485442e+09, 6.585513e+09, 6.685269e+09, 6.784643e+09, 6.883567e+09, 
    6.981969e+09, 7.079777e+09, 7.176916e+09, 7.273309e+09, 7.368877e+09, 
    7.463537e+09, 7.557208e+09, 7.649805e+09, 7.741242e+09, 7.831433e+09, 
    7.920287e+09, 8.007716e+09, 8.093629e+09, 8.177936e+09, 8.260545e+09, 
    8.341364e+09, 8.420301e+09, 8.497266e+09, 8.572165e+09, 8.64491e+09, 
    8.715411e+09, 8.78358e+09, 8.849328e+09, 8.912572e+09, 8.973229e+09, 
    9.031216e+09, 9.086456e+09, 9.138871e+09, 9.188391e+09, 9.234944e+09, 
    9.278465e+09, 9.318892e+09, 9.356163e+09, 9.390226e+09, 9.421031e+09, 
    9.448532e+09, 9.472687e+09, 9.49346e+09, 9.510819e+09, 9.524738e+09, 
    9.535196e+09, 9.542177e+09, 9.54567e+09, 9.54567e+09, 9.542177e+09, 
    9.535196e+09, 9.524738e+09, 9.510819e+09, 9.49346e+09, 9.472687e+09, 
    9.448532e+09, 9.421031e+09, 9.390226e+09, 9.356163e+09, 9.318892e+09, 
    9.278465e+09, 9.234944e+09, 9.188391e+09, 9.138871e+09, 9.086456e+09, 
    9.031216e+09, 8.973229e+09, 8.912572e+09, 8.849328e+09, 8.78358e+09, 
    8.715411e+09, 8.64491e+09, 8.572165e+09, 8.497266e+09, 8.420301e+09, 
    8.341364e+09, 8.260545e+09, 8.177936e+09, 8.093629e+09, 8.007716e+09, 
    7.920287e+09, 7.831433e+09, 7.741242e+09, 7.649805e+09, 7.557208e+09, 
    7.463537e+09, 7.368877e+09, 7.273309e+09, 7.176916e+09, 7.079777e+09, 
    6.981969e+09, 6.883567e+09, 6.784643e+09, 6.685269e+09, 6.585513e+09, 
    6.485442e+09,
  6.524282e+09, 6.627547e+09, 6.730571e+09, 6.833284e+09, 6.935614e+09, 
    7.037487e+09, 7.138825e+09, 7.23955e+09, 7.339579e+09, 7.438829e+09, 
    7.537212e+09, 7.634641e+09, 7.731025e+09, 7.826271e+09, 7.920287e+09, 
    8.012976e+09, 8.104243e+09, 8.193989e+09, 8.282116e+09, 8.368525e+09, 
    8.453116e+09, 8.53579e+09, 8.616447e+09, 8.694987e+09, 8.771312e+09, 
    8.845323e+09, 8.916924e+09, 8.986021e+09, 9.052518e+09, 9.116325e+09, 
    9.177352e+09, 9.235513e+09, 9.290724e+09, 9.342905e+09, 9.391978e+09, 
    9.437871e+09, 9.480515e+09, 9.519842e+09, 9.555794e+09, 9.588315e+09, 
    9.617354e+09, 9.642865e+09, 9.664807e+09, 9.683147e+09, 9.697854e+09, 
    9.708905e+09, 9.716282e+09, 9.719975e+09, 9.719975e+09, 9.716282e+09, 
    9.708905e+09, 9.697854e+09, 9.683147e+09, 9.664807e+09, 9.642865e+09, 
    9.617354e+09, 9.588315e+09, 9.555794e+09, 9.519842e+09, 9.480515e+09, 
    9.437871e+09, 9.391978e+09, 9.342905e+09, 9.290724e+09, 9.235513e+09, 
    9.177352e+09, 9.116325e+09, 9.052518e+09, 8.986021e+09, 8.916924e+09, 
    8.845323e+09, 8.771312e+09, 8.694987e+09, 8.616447e+09, 8.53579e+09, 
    8.453116e+09, 8.368525e+09, 8.282116e+09, 8.193989e+09, 8.104243e+09, 
    8.012976e+09, 7.920287e+09, 7.826271e+09, 7.731025e+09, 7.634641e+09, 
    7.537212e+09, 7.438829e+09, 7.339579e+09, 7.23955e+09, 7.138825e+09, 
    7.037487e+09, 6.935614e+09, 6.833284e+09, 6.730571e+09, 6.627547e+09, 
    6.524282e+09,
  6.562035e+09, 6.668449e+09, 6.774699e+09, 6.880711e+09, 6.986412e+09, 
    7.091722e+09, 7.196561e+09, 7.300845e+09, 7.404488e+09, 7.5074e+09, 
    7.60949e+09, 7.710664e+09, 7.810825e+09, 7.909876e+09, 8.007716e+09, 
    8.104243e+09, 8.199353e+09, 8.292941e+09, 8.384902e+09, 8.475127e+09, 
    8.563511e+09, 8.649944e+09, 8.734319e+09, 8.816526e+09, 8.896461e+09, 
    8.974015e+09, 9.049084e+09, 9.121564e+09, 9.191351e+09, 9.258346e+09, 
    9.322452e+09, 9.383574e+09, 9.441618e+09, 9.496498e+09, 9.548129e+09, 
    9.596429e+09, 9.641325e+09, 9.68274e+09, 9.720613e+09, 9.754878e+09, 
    9.785482e+09, 9.812372e+09, 9.835507e+09, 9.854844e+09, 9.870353e+09, 
    9.882009e+09, 9.88979e+09, 9.893683e+09, 9.893683e+09, 9.88979e+09, 
    9.882009e+09, 9.870353e+09, 9.854844e+09, 9.835507e+09, 9.812372e+09, 
    9.785482e+09, 9.754878e+09, 9.720613e+09, 9.68274e+09, 9.641325e+09, 
    9.596429e+09, 9.548129e+09, 9.496498e+09, 9.441618e+09, 9.383574e+09, 
    9.322452e+09, 9.258346e+09, 9.191351e+09, 9.121564e+09, 9.049084e+09, 
    8.974015e+09, 8.896461e+09, 8.816526e+09, 8.734319e+09, 8.649944e+09, 
    8.563511e+09, 8.475127e+09, 8.384902e+09, 8.292941e+09, 8.199353e+09, 
    8.104243e+09, 8.007716e+09, 7.909876e+09, 7.810825e+09, 7.710664e+09, 
    7.60949e+09, 7.5074e+09, 7.404488e+09, 7.300845e+09, 7.196561e+09, 
    7.091722e+09, 6.986412e+09, 6.880711e+09, 6.774699e+09, 6.668449e+09, 
    6.562035e+09,
  6.598693e+09, 6.708208e+09, 6.817636e+09, 6.926904e+09, 7.035934e+09, 
    7.144643e+09, 7.252946e+09, 7.360757e+09, 7.467984e+09, 7.574533e+09, 
    7.680307e+09, 7.785207e+09, 7.889131e+09, 7.991974e+09, 8.093629e+09, 
    8.193989e+09, 8.292941e+09, 8.390374e+09, 8.486173e+09, 8.580225e+09, 
    8.672412e+09, 8.762619e+09, 8.85073e+09, 8.936627e+09, 9.020195e+09, 
    9.101317e+09, 9.17988e+09, 9.255772e+09, 9.32888e+09, 9.399095e+09, 
    9.466312e+09, 9.530426e+09, 9.591338e+09, 9.64895e+09, 9.703171e+09, 
    9.753911e+09, 9.801088e+09, 9.844622e+09, 9.884442e+09, 9.920478e+09, 
    9.95267e+09, 9.980962e+09, 1.00053e+10, 1.002566e+10, 1.004198e+10, 
    1.005425e+10, 1.006244e+10, 1.006654e+10, 1.006654e+10, 1.006244e+10, 
    1.005425e+10, 1.004198e+10, 1.002566e+10, 1.00053e+10, 9.980962e+09, 
    9.95267e+09, 9.920478e+09, 9.884442e+09, 9.844622e+09, 9.801088e+09, 
    9.753911e+09, 9.703171e+09, 9.64895e+09, 9.591338e+09, 9.530426e+09, 
    9.466312e+09, 9.399095e+09, 9.32888e+09, 9.255772e+09, 9.17988e+09, 
    9.101317e+09, 9.020195e+09, 8.936627e+09, 8.85073e+09, 8.762619e+09, 
    8.672412e+09, 8.580225e+09, 8.486173e+09, 8.390374e+09, 8.292941e+09, 
    8.193989e+09, 8.093629e+09, 7.991974e+09, 7.889131e+09, 7.785207e+09, 
    7.680307e+09, 7.574533e+09, 7.467984e+09, 7.360757e+09, 7.252946e+09, 
    7.144643e+09, 7.035934e+09, 6.926904e+09, 6.817636e+09, 6.708208e+09, 
    6.598693e+09,
  6.634248e+09, 6.74681e+09, 6.859367e+09, 6.971842e+09, 7.084154e+09, 
    7.196217e+09, 7.307944e+09, 7.419243e+09, 7.530018e+09, 7.640172e+09, 
    7.749601e+09, 7.858201e+09, 7.965864e+09, 8.072481e+09, 8.177936e+09, 
    8.282116e+09, 8.384902e+09, 8.486173e+09, 8.585809e+09, 8.683688e+09, 
    8.779684e+09, 8.873673e+09, 8.96553e+09, 9.055129e+09, 9.142345e+09, 
    9.227054e+09, 9.309132e+09, 9.388457e+09, 9.464909e+09, 9.53837e+09, 
    9.608722e+09, 9.675857e+09, 9.739662e+09, 9.800034e+09, 9.856871e+09, 
    9.910078e+09, 9.959563e+09, 1.000524e+10, 1.004703e+10, 1.008486e+10, 
    1.011866e+10, 1.014837e+10, 1.017394e+10, 1.019532e+10, 1.021247e+10, 
    1.022536e+10, 1.023397e+10, 1.023827e+10, 1.023827e+10, 1.023397e+10, 
    1.022536e+10, 1.021247e+10, 1.019532e+10, 1.017394e+10, 1.014837e+10, 
    1.011866e+10, 1.008486e+10, 1.004703e+10, 1.000524e+10, 9.959563e+09, 
    9.910078e+09, 9.856871e+09, 9.800034e+09, 9.739662e+09, 9.675857e+09, 
    9.608722e+09, 9.53837e+09, 9.464909e+09, 9.388457e+09, 9.309132e+09, 
    9.227054e+09, 9.142345e+09, 9.055129e+09, 8.96553e+09, 8.873673e+09, 
    8.779684e+09, 8.683688e+09, 8.585809e+09, 8.486173e+09, 8.384902e+09, 
    8.282116e+09, 8.177936e+09, 8.072481e+09, 7.965864e+09, 7.858201e+09, 
    7.749601e+09, 7.640172e+09, 7.530018e+09, 7.419243e+09, 7.307944e+09, 
    7.196217e+09, 7.084154e+09, 6.971842e+09, 6.859367e+09, 6.74681e+09, 
    6.634248e+09,
  6.668692e+09, 6.784244e+09, 6.899874e+09, 7.015503e+09, 7.131045e+09, 
    7.246414e+09, 7.361518e+09, 7.47626e+09, 7.590542e+09, 7.704261e+09, 
    7.817309e+09, 7.929576e+09, 8.04095e+09, 8.151313e+09, 8.260545e+09, 
    8.368525e+09, 8.475127e+09, 8.580225e+09, 8.683688e+09, 8.785385e+09, 
    8.885187e+09, 8.982957e+09, 9.078562e+09, 9.171869e+09, 9.262742e+09, 
    9.351046e+09, 9.436652e+09, 9.519426e+09, 9.599237e+09, 9.67596e+09, 
    9.749469e+09, 9.819643e+09, 9.886363e+09, 9.949515e+09, 1.000899e+10, 
    1.006469e+10, 1.01165e+10, 1.016434e+10, 1.020812e+10, 1.024776e+10, 
    1.028319e+10, 1.031433e+10, 1.034114e+10, 1.036355e+10, 1.038154e+10, 
    1.039506e+10, 1.040409e+10, 1.040861e+10, 1.040861e+10, 1.040409e+10, 
    1.039506e+10, 1.038154e+10, 1.036355e+10, 1.034114e+10, 1.031433e+10, 
    1.028319e+10, 1.024776e+10, 1.020812e+10, 1.016434e+10, 1.01165e+10, 
    1.006469e+10, 1.000899e+10, 9.949515e+09, 9.886363e+09, 9.819643e+09, 
    9.749469e+09, 9.67596e+09, 9.599237e+09, 9.519426e+09, 9.436652e+09, 
    9.351046e+09, 9.262742e+09, 9.171869e+09, 9.078562e+09, 8.982957e+09, 
    8.885187e+09, 8.785385e+09, 8.683688e+09, 8.580225e+09, 8.475127e+09, 
    8.368525e+09, 8.260545e+09, 8.151313e+09, 8.04095e+09, 7.929576e+09, 
    7.817309e+09, 7.704261e+09, 7.590542e+09, 7.47626e+09, 7.361518e+09, 
    7.246414e+09, 7.131045e+09, 7.015503e+09, 6.899874e+09, 6.784244e+09, 
    6.668692e+09,
  6.702019e+09, 6.8205e+09, 6.939143e+09, 7.057866e+09, 7.176583e+09, 
    7.295202e+09, 7.41363e+09, 7.531766e+09, 7.649507e+09, 7.766745e+09, 
    7.883369e+09, 7.999264e+09, 8.11431e+09, 8.228386e+09, 8.341364e+09, 
    8.453116e+09, 8.563511e+09, 8.672412e+09, 8.779684e+09, 8.885187e+09, 
    8.988781e+09, 9.090322e+09, 9.18967e+09, 9.286681e+09, 9.381209e+09, 
    9.473112e+09, 9.562249e+09, 9.648477e+09, 9.731658e+09, 9.811654e+09, 
    9.88833e+09, 9.961556e+09, 1.00312e+10, 1.009715e+10, 1.015928e+10, 
    1.021748e+10, 1.027164e+10, 1.032166e+10, 1.036744e+10, 1.040891e+10, 
    1.044597e+10, 1.047856e+10, 1.050662e+10, 1.053008e+10, 1.054891e+10, 
    1.056306e+10, 1.057252e+10, 1.057725e+10, 1.057725e+10, 1.057252e+10, 
    1.056306e+10, 1.054891e+10, 1.053008e+10, 1.050662e+10, 1.047856e+10, 
    1.044597e+10, 1.040891e+10, 1.036744e+10, 1.032166e+10, 1.027164e+10, 
    1.021748e+10, 1.015928e+10, 1.009715e+10, 1.00312e+10, 9.961556e+09, 
    9.88833e+09, 9.811654e+09, 9.731658e+09, 9.648477e+09, 9.562249e+09, 
    9.473112e+09, 9.381209e+09, 9.286681e+09, 9.18967e+09, 9.090322e+09, 
    8.988781e+09, 8.885187e+09, 8.779684e+09, 8.672412e+09, 8.563511e+09, 
    8.453116e+09, 8.341364e+09, 8.228386e+09, 8.11431e+09, 7.999264e+09, 
    7.883369e+09, 7.766745e+09, 7.649507e+09, 7.531766e+09, 7.41363e+09, 
    7.295202e+09, 7.176583e+09, 7.057866e+09, 6.939143e+09, 6.8205e+09, 
    6.702019e+09,
  6.734221e+09, 6.855565e+09, 6.977157e+09, 7.098912e+09, 7.220742e+09, 
    7.342552e+09, 7.464245e+09, 7.585717e+09, 7.706863e+09, 7.827569e+09, 
    7.94772e+09, 8.067195e+09, 8.18587e+09, 8.303616e+09, 8.420301e+09, 
    8.53579e+09, 8.649944e+09, 8.762619e+09, 8.873673e+09, 8.982957e+09, 
    9.090322e+09, 9.195619e+09, 9.298694e+09, 9.399396e+09, 9.497571e+09, 
    9.593066e+09, 9.68573e+09, 9.775411e+09, 9.861961e+09, 9.945231e+09, 
    1.002508e+10, 1.010136e+10, 1.017395e+10, 1.02427e+10, 1.030749e+10, 
    1.03682e+10, 1.042471e+10, 1.047692e+10, 1.052472e+10, 1.056802e+10, 
    1.060673e+10, 1.064077e+10, 1.067009e+10, 1.06946e+10, 1.071428e+10, 
    1.072907e+10, 1.073895e+10, 1.07439e+10, 1.07439e+10, 1.073895e+10, 
    1.072907e+10, 1.071428e+10, 1.06946e+10, 1.067009e+10, 1.064077e+10, 
    1.060673e+10, 1.056802e+10, 1.052472e+10, 1.047692e+10, 1.042471e+10, 
    1.03682e+10, 1.030749e+10, 1.02427e+10, 1.017395e+10, 1.010136e+10, 
    1.002508e+10, 9.945231e+09, 9.861961e+09, 9.775411e+09, 9.68573e+09, 
    9.593066e+09, 9.497571e+09, 9.399396e+09, 9.298694e+09, 9.195619e+09, 
    9.090322e+09, 8.982957e+09, 8.873673e+09, 8.762619e+09, 8.649944e+09, 
    8.53579e+09, 8.420301e+09, 8.303616e+09, 8.18587e+09, 8.067195e+09, 
    7.94772e+09, 7.827569e+09, 7.706863e+09, 7.585717e+09, 7.464245e+09, 
    7.342552e+09, 7.220742e+09, 7.098912e+09, 6.977157e+09, 6.855565e+09, 
    6.734221e+09,
  6.76529e+09, 6.889429e+09, 7.013901e+09, 7.13862e+09, 7.263496e+09, 
    7.388432e+09, 7.513327e+09, 7.638074e+09, 7.762563e+09, 7.886679e+09, 
    8.010299e+09, 8.133301e+09, 8.255552e+09, 8.37692e+09, 8.497266e+09, 
    8.616447e+09, 8.734319e+09, 8.85073e+09, 8.96553e+09, 9.078562e+09, 
    9.18967e+09, 9.298694e+09, 9.405474e+09, 9.509846e+09, 9.61165e+09, 
    9.710721e+09, 9.806899e+09, 9.900023e+09, 9.989933e+09, 1.007647e+10, 
    1.015949e+10, 1.023883e+10, 1.031435e+10, 1.03859e+10, 1.045336e+10, 
    1.051658e+10, 1.057545e+10, 1.062985e+10, 1.067967e+10, 1.07248e+10, 
    1.076517e+10, 1.080067e+10, 1.083124e+10, 1.085682e+10, 1.087735e+10, 
    1.089278e+10, 1.090309e+10, 1.090825e+10, 1.090825e+10, 1.090309e+10, 
    1.089278e+10, 1.087735e+10, 1.085682e+10, 1.083124e+10, 1.080067e+10, 
    1.076517e+10, 1.07248e+10, 1.067967e+10, 1.062985e+10, 1.057545e+10, 
    1.051658e+10, 1.045336e+10, 1.03859e+10, 1.031435e+10, 1.023883e+10, 
    1.015949e+10, 1.007647e+10, 9.989933e+09, 9.900023e+09, 9.806899e+09, 
    9.710721e+09, 9.61165e+09, 9.509846e+09, 9.405474e+09, 9.298694e+09, 
    9.18967e+09, 9.078562e+09, 8.96553e+09, 8.85073e+09, 8.734319e+09, 
    8.616447e+09, 8.497266e+09, 8.37692e+09, 8.255552e+09, 8.133301e+09, 
    8.010299e+09, 7.886679e+09, 7.762563e+09, 7.638074e+09, 7.513327e+09, 
    7.388432e+09, 7.263496e+09, 7.13862e+09, 7.013901e+09, 6.889429e+09, 
    6.76529e+09,
  6.795221e+09, 6.922081e+09, 7.049361e+09, 7.176973e+09, 7.304823e+09, 
    7.432814e+09, 7.56084e+09, 7.688794e+09, 7.816561e+09, 7.94402e+09, 
    8.071048e+09, 8.197513e+09, 8.323282e+09, 8.448214e+09, 8.572165e+09, 
    8.694987e+09, 8.816526e+09, 8.936627e+09, 9.055129e+09, 9.171869e+09, 
    9.286681e+09, 9.399396e+09, 9.509846e+09, 9.61786e+09, 9.723264e+09, 
    9.825887e+09, 9.925557e+09, 1.00221e+10, 1.011536e+10, 1.020515e+10, 
    1.029132e+10, 1.037371e+10, 1.045215e+10, 1.05265e+10, 1.059662e+10, 
    1.066235e+10, 1.072358e+10, 1.078017e+10, 1.0832e+10, 1.087898e+10, 
    1.092099e+10, 1.095795e+10, 1.098979e+10, 1.101642e+10, 1.10378e+10, 
    1.105388e+10, 1.106461e+10, 1.106999e+10, 1.106999e+10, 1.106461e+10, 
    1.105388e+10, 1.10378e+10, 1.101642e+10, 1.098979e+10, 1.095795e+10, 
    1.092099e+10, 1.087898e+10, 1.0832e+10, 1.078017e+10, 1.072358e+10, 
    1.066235e+10, 1.059662e+10, 1.05265e+10, 1.045215e+10, 1.037371e+10, 
    1.029132e+10, 1.020515e+10, 1.011536e+10, 1.00221e+10, 9.925557e+09, 
    9.825887e+09, 9.723264e+09, 9.61786e+09, 9.509846e+09, 9.399396e+09, 
    9.286681e+09, 9.171869e+09, 9.055129e+09, 8.936627e+09, 8.816526e+09, 
    8.694987e+09, 8.572165e+09, 8.448214e+09, 8.323282e+09, 8.197513e+09, 
    8.071048e+09, 7.94402e+09, 7.816561e+09, 7.688794e+09, 7.56084e+09, 
    7.432814e+09, 7.304823e+09, 7.176973e+09, 7.049361e+09, 6.922081e+09, 
    6.795221e+09,
  6.824007e+09, 6.953512e+09, 7.083523e+09, 7.21395e+09, 7.344698e+09, 
    7.475667e+09, 7.606751e+09, 7.737838e+09, 7.868808e+09, 7.99954e+09, 
    8.129904e+09, 8.259766e+09, 8.388985e+09, 8.517416e+09, 8.64491e+09, 
    8.771312e+09, 8.896461e+09, 9.020195e+09, 9.142345e+09, 9.262742e+09, 
    9.381209e+09, 9.497571e+09, 9.61165e+09, 9.723264e+09, 9.832232e+09, 
    9.938373e+09, 1.00415e+10, 1.014144e+10, 1.023802e+10, 1.033104e+10, 
    1.042034e+10, 1.050575e+10, 1.058711e+10, 1.066424e+10, 1.0737e+10, 
    1.080523e+10, 1.08688e+10, 1.092757e+10, 1.098142e+10, 1.103023e+10, 
    1.107389e+10, 1.111231e+10, 1.11454e+10, 1.117309e+10, 1.119532e+10, 
    1.121203e+10, 1.12232e+10, 1.122879e+10, 1.122879e+10, 1.12232e+10, 
    1.121203e+10, 1.119532e+10, 1.117309e+10, 1.11454e+10, 1.111231e+10, 
    1.107389e+10, 1.103023e+10, 1.098142e+10, 1.092757e+10, 1.08688e+10, 
    1.080523e+10, 1.0737e+10, 1.066424e+10, 1.058711e+10, 1.050575e+10, 
    1.042034e+10, 1.033104e+10, 1.023802e+10, 1.014144e+10, 1.00415e+10, 
    9.938373e+09, 9.832232e+09, 9.723264e+09, 9.61165e+09, 9.497571e+09, 
    9.381209e+09, 9.26274e+09, 9.142345e+09, 9.020195e+09, 8.896461e+09, 
    8.771312e+09, 8.64491e+09, 8.517416e+09, 8.388985e+09, 8.259766e+09, 
    8.129904e+09, 7.99954e+09, 7.868808e+09, 7.737838e+09, 7.606751e+09, 
    7.475667e+09, 7.344698e+09, 7.21395e+09, 7.083523e+09, 6.953512e+09, 
    6.824007e+09,
  6.851641e+09, 6.98371e+09, 7.116371e+09, 7.249533e+09, 7.383099e+09, 
    7.516966e+09, 7.651027e+09, 7.785166e+09, 7.919261e+09, 8.053188e+09, 
    8.186811e+09, 8.319992e+09, 8.452588e+09, 8.584445e+09, 8.715411e+09, 
    8.845323e+09, 8.974015e+09, 9.101317e+09, 9.227054e+09, 9.351046e+09, 
    9.473112e+09, 9.593066e+09, 9.710721e+09, 9.825887e+09, 9.938373e+09, 
    1.004799e+10, 1.015454e+10, 1.025783e+10, 1.035769e+10, 1.045391e+10, 
    1.054631e+10, 1.063472e+10, 1.071896e+10, 1.079885e+10, 1.087423e+10, 
    1.094495e+10, 1.101085e+10, 1.107179e+10, 1.112763e+10, 1.117826e+10, 
    1.122356e+10, 1.126342e+10, 1.129776e+10, 1.13265e+10, 1.134958e+10, 
    1.136693e+10, 1.137852e+10, 1.138432e+10, 1.138432e+10, 1.137852e+10, 
    1.136693e+10, 1.134958e+10, 1.13265e+10, 1.129776e+10, 1.126342e+10, 
    1.122356e+10, 1.117826e+10, 1.112763e+10, 1.107179e+10, 1.101085e+10, 
    1.094495e+10, 1.087423e+10, 1.079885e+10, 1.071896e+10, 1.063472e+10, 
    1.054631e+10, 1.045391e+10, 1.035769e+10, 1.025783e+10, 1.015454e+10, 
    1.004799e+10, 9.938373e+09, 9.825887e+09, 9.710721e+09, 9.593066e+09, 
    9.473112e+09, 9.351046e+09, 9.227054e+09, 9.101317e+09, 8.974015e+09, 
    8.845323e+09, 8.715411e+09, 8.584445e+09, 8.452588e+09, 8.319992e+09, 
    8.186811e+09, 8.053188e+09, 7.919261e+09, 7.785166e+09, 7.651027e+09, 
    7.516966e+09, 7.383099e+09, 7.249533e+09, 7.116371e+09, 6.98371e+09, 
    6.851641e+09,
  6.878117e+09, 7.012667e+09, 7.147894e+09, 7.283705e+09, 7.420003e+09, 
    7.556683e+09, 7.693634e+09, 7.830739e+09, 7.967875e+09, 8.10491e+09, 
    8.241709e+09, 8.378128e+09, 8.514017e+09, 8.649221e+09, 8.78358e+09, 
    8.916924e+09, 9.049084e+09, 9.17988e+09, 9.309132e+09, 9.436652e+09, 
    9.562249e+09, 9.68573e+09, 9.806899e+09, 9.925557e+09, 1.00415e+10, 
    1.015454e+10, 1.026446e+10, 1.037106e+10, 1.047415e+10, 1.057352e+10, 
    1.066899e+10, 1.076036e+10, 1.084745e+10, 1.093007e+10, 1.100805e+10, 
    1.108122e+10, 1.114942e+10, 1.12125e+10, 1.127033e+10, 1.132276e+10, 
    1.136968e+10, 1.141097e+10, 1.144656e+10, 1.147634e+10, 1.150025e+10, 
    1.151823e+10, 1.153025e+10, 1.153626e+10, 1.153626e+10, 1.153025e+10, 
    1.151823e+10, 1.150025e+10, 1.147634e+10, 1.144656e+10, 1.141097e+10, 
    1.136968e+10, 1.132276e+10, 1.127033e+10, 1.12125e+10, 1.114942e+10, 
    1.108122e+10, 1.100805e+10, 1.093007e+10, 1.084745e+10, 1.076036e+10, 
    1.066899e+10, 1.057352e+10, 1.047415e+10, 1.037106e+10, 1.026446e+10, 
    1.015454e+10, 1.00415e+10, 9.925557e+09, 9.806899e+09, 9.68573e+09, 
    9.562249e+09, 9.436652e+09, 9.309132e+09, 9.17988e+09, 9.049084e+09, 
    8.916924e+09, 8.78358e+09, 8.649221e+09, 8.514017e+09, 8.378128e+09, 
    8.241709e+09, 8.10491e+09, 7.967875e+09, 7.830739e+09, 7.693634e+09, 
    7.556683e+09, 7.420003e+09, 7.283705e+09, 7.147894e+09, 7.012667e+09, 
    6.878117e+09,
  6.903431e+09, 7.040374e+09, 7.178077e+09, 7.316448e+09, 7.455388e+09, 
    7.594789e+09, 7.734541e+09, 7.874522e+09, 8.014606e+09, 8.15466e+09, 
    8.294543e+09, 8.434108e+09, 8.573202e+09, 8.711665e+09, 8.849328e+09, 
    8.986021e+09, 9.121564e+09, 9.255772e+09, 9.388457e+09, 9.519426e+09, 
    9.648477e+09, 9.775411e+09, 9.900023e+09, 1.00221e+10, 1.014144e+10, 
    1.025783e+10, 1.037106e+10, 1.048091e+10, 1.058718e+10, 1.068966e+10, 
    1.078814e+10, 1.088243e+10, 1.097232e+10, 1.105763e+10, 1.113816e+10, 
    1.121375e+10, 1.128423e+10, 1.134943e+10, 1.14092e+10, 1.146341e+10, 
    1.151193e+10, 1.155465e+10, 1.159146e+10, 1.162227e+10, 1.164701e+10, 
    1.166561e+10, 1.167804e+10, 1.168427e+10, 1.168427e+10, 1.167804e+10, 
    1.166561e+10, 1.164701e+10, 1.162227e+10, 1.159146e+10, 1.155465e+10, 
    1.151193e+10, 1.146341e+10, 1.14092e+10, 1.134943e+10, 1.128423e+10, 
    1.121375e+10, 1.113816e+10, 1.105763e+10, 1.097232e+10, 1.088243e+10, 
    1.078814e+10, 1.068966e+10, 1.058718e+10, 1.048091e+10, 1.037106e+10, 
    1.025783e+10, 1.014144e+10, 1.00221e+10, 9.900023e+09, 9.775411e+09, 
    9.648477e+09, 9.519426e+09, 9.388457e+09, 9.255772e+09, 9.121564e+09, 
    8.986021e+09, 8.849328e+09, 8.711665e+09, 8.573202e+09, 8.434108e+09, 
    8.294543e+09, 8.15466e+09, 8.014606e+09, 7.874522e+09, 7.734541e+09, 
    7.594789e+09, 7.455388e+09, 7.316448e+09, 7.178077e+09, 7.040374e+09, 
    6.903431e+09,
  6.927576e+09, 7.066821e+09, 7.206909e+09, 7.347746e+09, 7.489233e+09, 
    7.631261e+09, 7.773715e+09, 7.916475e+09, 8.059411e+09, 8.202386e+09, 
    8.345257e+09, 8.487873e+09, 8.630074e+09, 8.771699e+09, 8.912572e+09, 
    9.052518e+09, 9.191351e+09, 9.32888e+09, 9.464909e+09, 9.599237e+09, 
    9.731658e+09, 9.861961e+09, 9.989933e+09, 1.011536e+10, 1.023802e+10, 
    1.035769e+10, 1.047415e+10, 1.058718e+10, 1.069657e+10, 1.080209e+10, 
    1.090352e+10, 1.100067e+10, 1.109331e+10, 1.118125e+10, 1.12643e+10, 
    1.134227e+10, 1.141498e+10, 1.148226e+10, 1.154395e+10, 1.159992e+10, 
    1.165001e+10, 1.169412e+10, 1.173213e+10, 1.176396e+10, 1.178951e+10, 
    1.180873e+10, 1.182158e+10, 1.1828e+10, 1.1828e+10, 1.182158e+10, 
    1.180873e+10, 1.178951e+10, 1.176396e+10, 1.173213e+10, 1.169412e+10, 
    1.165001e+10, 1.159992e+10, 1.154395e+10, 1.148226e+10, 1.141498e+10, 
    1.134227e+10, 1.12643e+10, 1.118125e+10, 1.109331e+10, 1.100067e+10, 
    1.090352e+10, 1.080209e+10, 1.069657e+10, 1.058718e+10, 1.047415e+10, 
    1.035769e+10, 1.023802e+10, 1.011536e+10, 9.989933e+09, 9.861961e+09, 
    9.731658e+09, 9.599237e+09, 9.464909e+09, 9.32888e+09, 9.191351e+09, 
    9.052518e+09, 8.912572e+09, 8.771699e+09, 8.630074e+09, 8.487873e+09, 
    8.345257e+09, 8.202386e+09, 8.059411e+09, 7.916475e+09, 7.773715e+09, 
    7.631261e+09, 7.489233e+09, 7.347746e+09, 7.206909e+09, 7.066821e+09, 
    6.927576e+09,
  6.950547e+09, 7.092e+09, 7.234377e+09, 7.377583e+09, 7.521518e+09, 
    7.666072e+09, 7.811129e+09, 7.956566e+09, 8.10225e+09, 8.248043e+09, 
    8.393798e+09, 8.539359e+09, 8.684566e+09, 8.829247e+09, 8.973229e+09, 
    9.116325e+09, 9.258346e+09, 9.399095e+09, 9.53837e+09, 9.67596e+09, 
    9.811654e+09, 9.945231e+09, 1.007647e+10, 1.020515e+10, 1.033104e+10, 
    1.045391e+10, 1.057352e+10, 1.068966e+10, 1.080209e+10, 1.091057e+10, 
    1.10149e+10, 1.111483e+10, 1.121017e+10, 1.130069e+10, 1.13862e+10, 
    1.146649e+10, 1.154138e+10, 1.16107e+10, 1.167428e+10, 1.173195e+10, 
    1.17836e+10, 1.182907e+10, 1.186826e+10, 1.190108e+10, 1.192743e+10, 
    1.194726e+10, 1.19605e+10, 1.196713e+10, 1.196713e+10, 1.19605e+10, 
    1.194726e+10, 1.192743e+10, 1.190108e+10, 1.186826e+10, 1.182907e+10, 
    1.17836e+10, 1.173195e+10, 1.167428e+10, 1.16107e+10, 1.154138e+10, 
    1.146649e+10, 1.13862e+10, 1.130069e+10, 1.121017e+10, 1.111483e+10, 
    1.10149e+10, 1.091057e+10, 1.080209e+10, 1.068966e+10, 1.057352e+10, 
    1.045391e+10, 1.033104e+10, 1.020515e+10, 1.007647e+10, 9.945231e+09, 
    9.811654e+09, 9.67596e+09, 9.53837e+09, 9.399095e+09, 9.258346e+09, 
    9.116325e+09, 8.973229e+09, 8.829247e+09, 8.684566e+09, 8.539359e+09, 
    8.393798e+09, 8.248043e+09, 8.10225e+09, 7.956566e+09, 7.811129e+09, 
    7.666072e+09, 7.521518e+09, 7.377583e+09, 7.234377e+09, 7.092e+09, 
    6.950547e+09,
  6.972339e+09, 7.115902e+09, 7.260469e+09, 7.405943e+09, 7.552224e+09, 
    7.699199e+09, 7.846753e+09, 7.994759e+09, 8.143084e+09, 8.291585e+09, 
    8.440113e+09, 8.58851e+09, 8.736609e+09, 8.884238e+09, 9.031216e+09, 
    9.177352e+09, 9.322452e+09, 9.466312e+09, 9.608722e+09, 9.749469e+09, 
    9.88833e+09, 1.002508e+10, 1.015949e+10, 1.029132e+10, 1.042034e+10, 
    1.054631e+10, 1.066899e+10, 1.078814e+10, 1.090352e+10, 1.10149e+10, 
    1.112203e+10, 1.122468e+10, 1.132264e+10, 1.141567e+10, 1.150357e+10, 
    1.158613e+10, 1.166315e+10, 1.173446e+10, 1.179987e+10, 1.185922e+10, 
    1.191237e+10, 1.195917e+10, 1.199952e+10, 1.203331e+10, 1.206044e+10, 
    1.208085e+10, 1.209449e+10, 1.210132e+10, 1.210132e+10, 1.209449e+10, 
    1.208085e+10, 1.206044e+10, 1.203331e+10, 1.199952e+10, 1.195917e+10, 
    1.191237e+10, 1.185922e+10, 1.179987e+10, 1.173446e+10, 1.166315e+10, 
    1.158613e+10, 1.150357e+10, 1.141567e+10, 1.132264e+10, 1.122468e+10, 
    1.112203e+10, 1.10149e+10, 1.090352e+10, 1.078814e+10, 1.066899e+10, 
    1.054631e+10, 1.042034e+10, 1.029132e+10, 1.015949e+10, 1.002508e+10, 
    9.88833e+09, 9.749469e+09, 9.608722e+09, 9.466312e+09, 9.322452e+09, 
    9.177352e+09, 9.031216e+09, 8.884238e+09, 8.736609e+09, 8.58851e+09, 
    8.440113e+09, 8.291585e+09, 8.143084e+09, 7.994759e+09, 7.846753e+09, 
    7.699199e+09, 7.552224e+09, 7.405943e+09, 7.260469e+09, 7.115902e+09, 
    6.972339e+09,
  6.992947e+09, 7.138521e+09, 7.285175e+09, 7.432813e+09, 7.581331e+09, 
    7.73062e+09, 7.880559e+09, 8.031022e+09, 8.181873e+09, 8.332967e+09, 
    8.484152e+09, 8.635267e+09, 8.786142e+09, 8.936601e+09, 9.086456e+09, 
    9.235513e+09, 9.383574e+09, 9.530426e+09, 9.675857e+09, 9.819643e+09, 
    9.961556e+09, 1.010136e+10, 1.023883e+10, 1.037371e+10, 1.050575e+10, 
    1.063472e+10, 1.076036e+10, 1.088243e+10, 1.100067e+10, 1.111483e+10, 
    1.122468e+10, 1.132997e+10, 1.143046e+10, 1.152593e+10, 1.161615e+10, 
    1.170091e+10, 1.178001e+10, 1.185324e+10, 1.192043e+10, 1.198141e+10, 
    1.203602e+10, 1.208412e+10, 1.212559e+10, 1.216031e+10, 1.218821e+10, 
    1.220919e+10, 1.222321e+10, 1.223023e+10, 1.223023e+10, 1.222321e+10, 
    1.220919e+10, 1.218821e+10, 1.216031e+10, 1.212559e+10, 1.208412e+10, 
    1.203602e+10, 1.198141e+10, 1.192043e+10, 1.185324e+10, 1.178001e+10, 
    1.170091e+10, 1.161615e+10, 1.152593e+10, 1.143046e+10, 1.132997e+10, 
    1.122468e+10, 1.111483e+10, 1.100067e+10, 1.088243e+10, 1.076036e+10, 
    1.063472e+10, 1.050575e+10, 1.037371e+10, 1.023883e+10, 1.010136e+10, 
    9.961556e+09, 9.819643e+09, 9.675857e+09, 9.530426e+09, 9.383574e+09, 
    9.235513e+09, 9.086456e+09, 8.936601e+09, 8.786142e+09, 8.635267e+09, 
    8.484152e+09, 8.332967e+09, 8.181873e+09, 8.031022e+09, 7.880559e+09, 
    7.73062e+09, 7.581331e+09, 7.432813e+09, 7.285175e+09, 7.138521e+09, 
    6.992947e+09,
  7.012366e+09, 7.159848e+09, 7.308484e+09, 7.458176e+09, 7.608822e+09, 
    7.760311e+09, 7.912521e+09, 8.065324e+09, 8.218582e+09, 8.372148e+09, 
    8.525868e+09, 8.679578e+09, 8.833104e+09, 8.986266e+09, 9.138871e+09, 
    9.290724e+09, 9.441618e+09, 9.591338e+09, 9.739662e+09, 9.886363e+09, 
    1.00312e+10, 1.017395e+10, 1.031435e+10, 1.045215e+10, 1.058711e+10, 
    1.071896e+10, 1.084745e+10, 1.097232e+10, 1.109331e+10, 1.121017e+10, 
    1.132264e+10, 1.143046e+10, 1.153341e+10, 1.163122e+10, 1.172369e+10, 
    1.181057e+10, 1.189166e+10, 1.196675e+10, 1.203567e+10, 1.209821e+10, 
    1.215424e+10, 1.220359e+10, 1.224615e+10, 1.228178e+10, 1.231041e+10, 
    1.233195e+10, 1.234634e+10, 1.235355e+10, 1.235355e+10, 1.234634e+10, 
    1.233195e+10, 1.231041e+10, 1.228178e+10, 1.224615e+10, 1.220359e+10, 
    1.215424e+10, 1.209821e+10, 1.203567e+10, 1.196675e+10, 1.189166e+10, 
    1.181057e+10, 1.172369e+10, 1.163122e+10, 1.153341e+10, 1.143046e+10, 
    1.132264e+10, 1.121017e+10, 1.109331e+10, 1.097232e+10, 1.084745e+10, 
    1.071896e+10, 1.058711e+10, 1.045215e+10, 1.031435e+10, 1.017395e+10, 
    1.00312e+10, 9.886363e+09, 9.739662e+09, 9.591338e+09, 9.441618e+09, 
    9.290724e+09, 9.138871e+09, 8.986266e+09, 8.833104e+09, 8.679578e+09, 
    8.525868e+09, 8.372148e+09, 8.218582e+09, 8.065324e+09, 7.912521e+09, 
    7.760311e+09, 7.608822e+09, 7.458176e+09, 7.308484e+09, 7.159848e+09, 
    7.012366e+09,
  7.030593e+09, 7.179877e+09, 7.330385e+09, 7.482021e+09, 7.634681e+09, 
    7.788252e+09, 7.942612e+09, 8.097633e+09, 8.253174e+09, 8.409087e+09, 
    8.565214e+09, 8.721389e+09, 8.877434e+09, 9.033167e+09, 9.188391e+09, 
    9.342905e+09, 9.496498e+09, 9.64895e+09, 9.800034e+09, 9.949515e+09, 
    1.009715e+10, 1.02427e+10, 1.03859e+10, 1.05265e+10, 1.066424e+10, 
    1.079885e+10, 1.093007e+10, 1.105763e+10, 1.118125e+10, 1.130069e+10, 
    1.141567e+10, 1.152593e+10, 1.163122e+10, 1.17313e+10, 1.182591e+10, 
    1.191483e+10, 1.199784e+10, 1.207473e+10, 1.214529e+10, 1.220935e+10, 
    1.226673e+10, 1.231729e+10, 1.236089e+10, 1.23974e+10, 1.242673e+10, 
    1.24488e+10, 1.246355e+10, 1.247093e+10, 1.247093e+10, 1.246355e+10, 
    1.24488e+10, 1.242673e+10, 1.23974e+10, 1.236089e+10, 1.231729e+10, 
    1.226673e+10, 1.220935e+10, 1.214529e+10, 1.207473e+10, 1.199784e+10, 
    1.191483e+10, 1.182591e+10, 1.17313e+10, 1.163122e+10, 1.152593e+10, 
    1.141567e+10, 1.130069e+10, 1.118125e+10, 1.105763e+10, 1.093007e+10, 
    1.079885e+10, 1.066424e+10, 1.05265e+10, 1.03859e+10, 1.02427e+10, 
    1.009715e+10, 9.949515e+09, 9.800034e+09, 9.64895e+09, 9.496498e+09, 
    9.342905e+09, 9.188391e+09, 9.033167e+09, 8.877434e+09, 8.721389e+09, 
    8.565214e+09, 8.409087e+09, 8.253174e+09, 8.097633e+09, 7.942612e+09, 
    7.788252e+09, 7.634681e+09, 7.482021e+09, 7.330385e+09, 7.179877e+09, 
    7.030593e+09,
  7.047623e+09, 7.198601e+09, 7.350871e+09, 7.504335e+09, 7.65889e+09, 
    7.814423e+09, 7.970811e+09, 8.127923e+09, 8.285618e+09, 8.443745e+09, 
    8.602145e+09, 8.760649e+09, 8.919077e+09, 9.077242e+09, 9.234944e+09, 
    9.391978e+09, 9.548129e+09, 9.703171e+09, 9.856871e+09, 1.000899e+10, 
    1.015928e+10, 1.030749e+10, 1.045336e+10, 1.059662e+10, 1.0737e+10, 
    1.087423e+10, 1.100805e+10, 1.113816e+10, 1.12643e+10, 1.13862e+10, 
    1.150357e+10, 1.161615e+10, 1.172369e+10, 1.182591e+10, 1.192258e+10, 
    1.201345e+10, 1.209829e+10, 1.217688e+10, 1.224902e+10, 1.231452e+10, 
    1.237321e+10, 1.242492e+10, 1.246951e+10, 1.250686e+10, 1.253687e+10, 
    1.255944e+10, 1.257453e+10, 1.258209e+10, 1.258209e+10, 1.257453e+10, 
    1.255944e+10, 1.253687e+10, 1.250686e+10, 1.246951e+10, 1.242492e+10, 
    1.237321e+10, 1.231452e+10, 1.224902e+10, 1.217688e+10, 1.209829e+10, 
    1.201345e+10, 1.192258e+10, 1.182591e+10, 1.172369e+10, 1.161615e+10, 
    1.150357e+10, 1.13862e+10, 1.12643e+10, 1.113816e+10, 1.100805e+10, 
    1.087423e+10, 1.0737e+10, 1.059662e+10, 1.045336e+10, 1.030749e+10, 
    1.015928e+10, 1.000899e+10, 9.856871e+09, 9.703171e+09, 9.548129e+09, 
    9.391978e+09, 9.234944e+09, 9.077242e+09, 8.919077e+09, 8.760649e+09, 
    8.602145e+09, 8.443745e+09, 8.285618e+09, 8.127923e+09, 7.970811e+09, 
    7.814423e+09, 7.65889e+09, 7.504335e+09, 7.350871e+09, 7.198601e+09, 
    7.047623e+09,
  7.063453e+09, 7.216014e+09, 7.36993e+09, 7.525106e+09, 7.681435e+09, 
    7.838806e+09, 7.997093e+09, 8.156166e+09, 8.31588e+09, 8.476086e+09, 
    8.636621e+09, 8.797313e+09, 8.95798e+09, 9.118431e+09, 9.278465e+09, 
    9.437871e+09, 9.596429e+09, 9.753911e+09, 9.910078e+09, 1.006469e+10, 
    1.021748e+10, 1.03682e+10, 1.051658e+10, 1.066235e+10, 1.080523e+10, 
    1.094495e+10, 1.108122e+10, 1.121375e+10, 1.134227e+10, 1.146649e+10, 
    1.158613e+10, 1.170091e+10, 1.181057e+10, 1.191483e+10, 1.201345e+10, 
    1.210616e+10, 1.219274e+10, 1.227295e+10, 1.234659e+10, 1.241347e+10, 
    1.247338e+10, 1.252618e+10, 1.257172e+10, 1.260987e+10, 1.264052e+10, 
    1.266358e+10, 1.267899e+10, 1.268671e+10, 1.268671e+10, 1.267899e+10, 
    1.266358e+10, 1.264052e+10, 1.260987e+10, 1.257172e+10, 1.252618e+10, 
    1.247338e+10, 1.241347e+10, 1.234659e+10, 1.227295e+10, 1.219274e+10, 
    1.210616e+10, 1.201345e+10, 1.191483e+10, 1.181057e+10, 1.170091e+10, 
    1.158613e+10, 1.146649e+10, 1.134227e+10, 1.121375e+10, 1.108122e+10, 
    1.094495e+10, 1.080523e+10, 1.066235e+10, 1.051658e+10, 1.03682e+10, 
    1.021748e+10, 1.006469e+10, 9.910078e+09, 9.753911e+09, 9.596429e+09, 
    9.437871e+09, 9.278465e+09, 9.118431e+09, 8.95798e+09, 8.797313e+09, 
    8.636621e+09, 8.476086e+09, 8.31588e+09, 8.156166e+09, 7.997093e+09, 
    7.838806e+09, 7.681435e+09, 7.525106e+09, 7.36993e+09, 7.216014e+09, 
    7.063453e+09,
  7.078078e+09, 7.23211e+09, 7.387556e+09, 7.544322e+09, 7.702302e+09, 
    7.861382e+09, 8.021437e+09, 8.182336e+09, 8.343933e+09, 8.506077e+09, 
    8.668601e+09, 8.831335e+09, 8.994092e+09, 9.156679e+09, 9.318892e+09, 
    9.480515e+09, 9.641325e+09, 9.801088e+09, 9.959563e+09, 1.01165e+10, 
    1.027164e+10, 1.042471e+10, 1.057545e+10, 1.072358e+10, 1.08688e+10, 
    1.101085e+10, 1.114942e+10, 1.128423e+10, 1.141498e+10, 1.154138e+10, 
    1.166315e+10, 1.178001e+10, 1.189166e+10, 1.199784e+10, 1.209829e+10, 
    1.219274e+10, 1.228095e+10, 1.236269e+10, 1.243775e+10, 1.250591e+10, 
    1.256699e+10, 1.262082e+10, 1.266725e+10, 1.270614e+10, 1.273739e+10, 
    1.276091e+10, 1.277663e+10, 1.27845e+10, 1.27845e+10, 1.277663e+10, 
    1.276091e+10, 1.273739e+10, 1.270614e+10, 1.266725e+10, 1.262082e+10, 
    1.256699e+10, 1.250591e+10, 1.243775e+10, 1.236269e+10, 1.228095e+10, 
    1.219274e+10, 1.209829e+10, 1.199784e+10, 1.189166e+10, 1.178001e+10, 
    1.166315e+10, 1.154138e+10, 1.141498e+10, 1.128423e+10, 1.114942e+10, 
    1.101085e+10, 1.08688e+10, 1.072358e+10, 1.057545e+10, 1.042471e+10, 
    1.027164e+10, 1.01165e+10, 9.959563e+09, 9.801088e+09, 9.641325e+09, 
    9.480515e+09, 9.318892e+09, 9.156679e+09, 8.994092e+09, 8.831335e+09, 
    8.668601e+09, 8.506077e+09, 8.343933e+09, 8.182336e+09, 8.021437e+09, 
    7.861382e+09, 7.702302e+09, 7.544322e+09, 7.387556e+09, 7.23211e+09, 
    7.078078e+09,
  7.091497e+09, 7.246883e+09, 7.403741e+09, 7.561974e+09, 7.721477e+09, 
    7.882135e+09, 8.043825e+09, 8.20641e+09, 8.369748e+09, 8.533684e+09, 
    8.698051e+09, 8.862674e+09, 9.027367e+09, 9.191932e+09, 9.356163e+09, 
    9.519842e+09, 9.68274e+09, 9.844622e+09, 1.000524e+10, 1.016434e+10, 
    1.032166e+10, 1.047692e+10, 1.062985e+10, 1.078017e+10, 1.092757e+10, 
    1.107179e+10, 1.12125e+10, 1.134943e+10, 1.148226e+10, 1.16107e+10, 
    1.173446e+10, 1.185324e+10, 1.196675e+10, 1.207473e+10, 1.217688e+10, 
    1.227295e+10, 1.236269e+10, 1.244586e+10, 1.252223e+10, 1.25916e+10, 
    1.265377e+10, 1.270856e+10, 1.275582e+10, 1.279542e+10, 1.282723e+10, 
    1.285118e+10, 1.286718e+10, 1.287519e+10, 1.287519e+10, 1.286718e+10, 
    1.285118e+10, 1.282723e+10, 1.279542e+10, 1.275582e+10, 1.270856e+10, 
    1.265377e+10, 1.25916e+10, 1.252223e+10, 1.244586e+10, 1.236269e+10, 
    1.227295e+10, 1.217688e+10, 1.207473e+10, 1.196675e+10, 1.185324e+10, 
    1.173446e+10, 1.16107e+10, 1.148226e+10, 1.134943e+10, 1.12125e+10, 
    1.107179e+10, 1.092757e+10, 1.078017e+10, 1.062985e+10, 1.047692e+10, 
    1.032166e+10, 1.016434e+10, 1.000524e+10, 9.844622e+09, 9.68274e+09, 
    9.519842e+09, 9.356163e+09, 9.191932e+09, 9.027367e+09, 8.862674e+09, 
    8.698051e+09, 8.533684e+09, 8.369748e+09, 8.20641e+09, 8.043825e+09, 
    7.882135e+09, 7.721477e+09, 7.561974e+09, 7.403741e+09, 7.246883e+09, 
    7.091497e+09,
  7.103705e+09, 7.260329e+09, 7.418477e+09, 7.578052e+09, 7.738948e+09, 
    7.901051e+09, 8.064236e+09, 8.228367e+09, 8.3933e+09, 8.558878e+09, 
    8.724934e+09, 8.891291e+09, 9.05776e+09, 9.224142e+09, 9.390226e+09, 
    9.555794e+09, 9.720613e+09, 9.884442e+09, 1.004703e+10, 1.020812e+10, 
    1.036744e+10, 1.052472e+10, 1.067967e+10, 1.0832e+10, 1.098142e+10, 
    1.112763e+10, 1.127033e+10, 1.14092e+10, 1.154395e+10, 1.167428e+10, 
    1.179987e+10, 1.192043e+10, 1.203567e+10, 1.214529e+10, 1.224902e+10, 
    1.234659e+10, 1.243775e+10, 1.252223e+10, 1.259983e+10, 1.267031e+10, 
    1.273348e+10, 1.278916e+10, 1.283719e+10, 1.287743e+10, 1.290977e+10, 
    1.293411e+10, 1.295038e+10, 1.295852e+10, 1.295852e+10, 1.295038e+10, 
    1.293411e+10, 1.290977e+10, 1.287743e+10, 1.283719e+10, 1.278916e+10, 
    1.273348e+10, 1.267031e+10, 1.259983e+10, 1.252223e+10, 1.243775e+10, 
    1.234659e+10, 1.224902e+10, 1.214529e+10, 1.203567e+10, 1.192043e+10, 
    1.179987e+10, 1.167428e+10, 1.154395e+10, 1.14092e+10, 1.127033e+10, 
    1.112763e+10, 1.098142e+10, 1.0832e+10, 1.067967e+10, 1.052472e+10, 
    1.036744e+10, 1.020812e+10, 1.004703e+10, 9.884442e+09, 9.720613e+09, 
    9.555794e+09, 9.390226e+09, 9.224142e+09, 9.05776e+09, 8.891291e+09, 
    8.724934e+09, 8.558878e+09, 8.3933e+09, 8.228367e+09, 8.064236e+09, 
    7.901051e+09, 7.738948e+09, 7.578052e+09, 7.418477e+09, 7.260329e+09, 
    7.103705e+09,
  7.1147e+09, 7.272444e+09, 7.431758e+09, 7.592547e+09, 7.754704e+09, 
    7.918115e+09, 8.082655e+09, 8.248187e+09, 8.414565e+09, 8.581632e+09, 
    8.749221e+09, 8.917151e+09, 9.085231e+09, 9.253263e+09, 9.421031e+09, 
    9.588315e+09, 9.754878e+09, 9.920478e+09, 1.008486e+10, 1.024776e+10, 
    1.040891e+10, 1.056802e+10, 1.07248e+10, 1.087898e+10, 1.103023e+10, 
    1.117826e+10, 1.132276e+10, 1.146341e+10, 1.159992e+10, 1.173195e+10, 
    1.185922e+10, 1.198141e+10, 1.209821e+10, 1.220935e+10, 1.231452e+10, 
    1.241347e+10, 1.250591e+10, 1.25916e+10, 1.267031e+10, 1.27418e+10, 
    1.280589e+10, 1.286239e+10, 1.291113e+10, 1.295196e+10, 1.298478e+10, 
    1.300948e+10, 1.302599e+10, 1.303425e+10, 1.303425e+10, 1.302599e+10, 
    1.300948e+10, 1.298478e+10, 1.295196e+10, 1.291113e+10, 1.286239e+10, 
    1.280589e+10, 1.27418e+10, 1.267031e+10, 1.25916e+10, 1.250591e+10, 
    1.241347e+10, 1.231452e+10, 1.220935e+10, 1.209821e+10, 1.198141e+10, 
    1.185922e+10, 1.173195e+10, 1.159992e+10, 1.146341e+10, 1.132276e+10, 
    1.117826e+10, 1.103023e+10, 1.087898e+10, 1.07248e+10, 1.056802e+10, 
    1.040891e+10, 1.024776e+10, 1.008486e+10, 9.920478e+09, 9.754878e+09, 
    9.588315e+09, 9.421031e+09, 9.253263e+09, 9.085231e+09, 8.917151e+09, 
    8.749221e+09, 8.581632e+09, 8.414565e+09, 8.248187e+09, 8.082655e+09, 
    7.918115e+09, 7.754704e+09, 7.592547e+09, 7.431758e+09, 7.272444e+09, 
    7.1147e+09,
  7.124479e+09, 7.283223e+09, 7.443579e+09, 7.605452e+09, 7.768736e+09, 
    7.933316e+09, 8.099066e+09, 8.26585e+09, 8.433522e+09, 8.601922e+09, 
    8.770882e+09, 8.940219e+09, 9.109745e+09, 9.279254e+09, 9.448532e+09, 
    9.617354e+09, 9.785482e+09, 9.95267e+09, 1.011866e+10, 1.028319e+10, 
    1.044597e+10, 1.060673e+10, 1.076517e+10, 1.092099e+10, 1.107389e+10, 
    1.122356e+10, 1.136968e+10, 1.151193e+10, 1.165001e+10, 1.17836e+10, 
    1.191237e+10, 1.203602e+10, 1.215424e+10, 1.226673e+10, 1.237321e+10, 
    1.247338e+10, 1.256699e+10, 1.265377e+10, 1.273348e+10, 1.280589e+10, 
    1.287081e+10, 1.292804e+10, 1.297741e+10, 1.301878e+10, 1.305203e+10, 
    1.307706e+10, 1.309378e+10, 1.310215e+10, 1.310215e+10, 1.309378e+10, 
    1.307706e+10, 1.305203e+10, 1.301878e+10, 1.297741e+10, 1.292804e+10, 
    1.287081e+10, 1.280589e+10, 1.273348e+10, 1.265377e+10, 1.256699e+10, 
    1.247338e+10, 1.237321e+10, 1.226673e+10, 1.215424e+10, 1.203602e+10, 
    1.191237e+10, 1.17836e+10, 1.165001e+10, 1.151193e+10, 1.136968e+10, 
    1.122356e+10, 1.107389e+10, 1.092099e+10, 1.076517e+10, 1.060673e+10, 
    1.044597e+10, 1.028319e+10, 1.011866e+10, 9.95267e+09, 9.785482e+09, 
    9.617354e+09, 9.448532e+09, 9.279254e+09, 9.109745e+09, 8.940219e+09, 
    8.770882e+09, 8.601922e+09, 8.433522e+09, 8.26585e+09, 8.099066e+09, 
    7.933316e+09, 7.768736e+09, 7.605452e+09, 7.443579e+09, 7.283223e+09, 
    7.124479e+09,
  7.133041e+09, 7.292662e+09, 7.453934e+09, 7.616759e+09, 7.781033e+09, 
    7.946641e+09, 8.113456e+09, 8.281342e+09, 8.450151e+09, 8.619724e+09, 
    8.789891e+09, 8.96047e+09, 9.131267e+09, 9.302078e+09, 9.472687e+09, 
    9.642865e+09, 9.812372e+09, 9.980962e+09, 1.014837e+10, 1.031433e+10, 
    1.047856e+10, 1.064077e+10, 1.080067e+10, 1.095795e+10, 1.111231e+10, 
    1.126342e+10, 1.141097e+10, 1.155465e+10, 1.169412e+10, 1.182907e+10, 
    1.195917e+10, 1.208412e+10, 1.220359e+10, 1.231729e+10, 1.242492e+10, 
    1.252618e+10, 1.262082e+10, 1.270856e+10, 1.278916e+10, 1.286239e+10, 
    1.292804e+10, 1.298592e+10, 1.303585e+10, 1.30777e+10, 1.311133e+10, 
    1.313664e+10, 1.315356e+10, 1.316203e+10, 1.316203e+10, 1.315356e+10, 
    1.313664e+10, 1.311133e+10, 1.30777e+10, 1.303585e+10, 1.298592e+10, 
    1.292804e+10, 1.286239e+10, 1.278916e+10, 1.270856e+10, 1.262082e+10, 
    1.252618e+10, 1.242492e+10, 1.231729e+10, 1.220359e+10, 1.208412e+10, 
    1.195917e+10, 1.182907e+10, 1.169412e+10, 1.155465e+10, 1.141097e+10, 
    1.126342e+10, 1.111231e+10, 1.095795e+10, 1.080067e+10, 1.064077e+10, 
    1.047856e+10, 1.031433e+10, 1.014837e+10, 9.980962e+09, 9.812372e+09, 
    9.642865e+09, 9.472687e+09, 9.302078e+09, 9.131267e+09, 8.96047e+09, 
    8.789891e+09, 8.619724e+09, 8.450151e+09, 8.281342e+09, 8.113456e+09, 
    7.946641e+09, 7.781033e+09, 7.616759e+09, 7.453934e+09, 7.292662e+09, 
    7.133041e+09,
  7.140384e+09, 7.30076e+09, 7.462817e+09, 7.626462e+09, 7.791588e+09, 
    7.958081e+09, 8.125813e+09, 8.294647e+09, 8.464436e+09, 8.63502e+09, 
    8.806228e+09, 8.977876e+09, 9.14977e+09, 9.321703e+09, 9.49346e+09, 
    9.664807e+09, 9.835507e+09, 1.00053e+10, 1.017394e+10, 1.034114e+10, 
    1.050662e+10, 1.067009e+10, 1.083124e+10, 1.098979e+10, 1.11454e+10, 
    1.129776e+10, 1.144656e+10, 1.159146e+10, 1.173213e+10, 1.186826e+10, 
    1.199952e+10, 1.212559e+10, 1.224615e+10, 1.236089e+10, 1.246951e+10, 
    1.257172e+10, 1.266725e+10, 1.275582e+10, 1.283719e+10, 1.291113e+10, 
    1.297741e+10, 1.303585e+10, 1.308628e+10, 1.312854e+10, 1.316249e+10, 
    1.318806e+10, 1.320514e+10, 1.32137e+10, 1.32137e+10, 1.320514e+10, 
    1.318806e+10, 1.316249e+10, 1.312854e+10, 1.308628e+10, 1.303585e+10, 
    1.297741e+10, 1.291113e+10, 1.283719e+10, 1.275582e+10, 1.266725e+10, 
    1.257172e+10, 1.246951e+10, 1.236089e+10, 1.224615e+10, 1.212559e+10, 
    1.199952e+10, 1.186826e+10, 1.173213e+10, 1.159146e+10, 1.144656e+10, 
    1.129776e+10, 1.11454e+10, 1.098979e+10, 1.083124e+10, 1.067009e+10, 
    1.050662e+10, 1.034114e+10, 1.017394e+10, 1.00053e+10, 9.835507e+09, 
    9.664807e+09, 9.49346e+09, 9.321703e+09, 9.14977e+09, 8.977876e+09, 
    8.806228e+09, 8.63502e+09, 8.464436e+09, 8.294647e+09, 8.125813e+09, 
    7.958081e+09, 7.791588e+09, 7.626462e+09, 7.462817e+09, 7.30076e+09, 
    7.140384e+09,
  7.146505e+09, 7.307511e+09, 7.470226e+09, 7.634556e+09, 7.800395e+09, 
    7.967627e+09, 8.136126e+09, 8.305754e+09, 8.476363e+09, 8.647793e+09, 
    8.819871e+09, 8.992415e+09, 9.165227e+09, 9.338102e+09, 9.510819e+09, 
    9.683147e+09, 9.854844e+09, 1.002566e+10, 1.019532e+10, 1.036355e+10, 
    1.053008e+10, 1.06946e+10, 1.085682e+10, 1.101642e+10, 1.117309e+10, 
    1.13265e+10, 1.147634e+10, 1.162227e+10, 1.176396e+10, 1.190108e+10, 
    1.203331e+10, 1.216031e+10, 1.228178e+10, 1.23974e+10, 1.250686e+10, 
    1.260987e+10, 1.270614e+10, 1.279542e+10, 1.287743e+10, 1.295196e+10, 
    1.301878e+10, 1.30777e+10, 1.312854e+10, 1.317114e+10, 1.320537e+10, 
    1.323115e+10, 1.324837e+10, 1.3257e+10, 1.3257e+10, 1.324837e+10, 
    1.323115e+10, 1.320537e+10, 1.317114e+10, 1.312854e+10, 1.30777e+10, 
    1.301878e+10, 1.295196e+10, 1.287743e+10, 1.279542e+10, 1.270614e+10, 
    1.260987e+10, 1.250686e+10, 1.23974e+10, 1.228178e+10, 1.216031e+10, 
    1.203331e+10, 1.190108e+10, 1.176396e+10, 1.162227e+10, 1.147634e+10, 
    1.13265e+10, 1.117309e+10, 1.101642e+10, 1.085682e+10, 1.06946e+10, 
    1.053008e+10, 1.036355e+10, 1.019532e+10, 1.002566e+10, 9.854844e+09, 
    9.683147e+09, 9.510819e+09, 9.338102e+09, 9.165227e+09, 8.992415e+09, 
    8.819871e+09, 8.647793e+09, 8.476363e+09, 8.305754e+09, 8.136126e+09, 
    7.967627e+09, 7.800395e+09, 7.634556e+09, 7.470226e+09, 7.307511e+09, 
    7.146505e+09,
  7.151404e+09, 7.312915e+09, 7.476158e+09, 7.641037e+09, 7.807448e+09, 
    7.975273e+09, 8.144387e+09, 8.314652e+09, 8.485919e+09, 8.658028e+09, 
    8.830806e+09, 9.004068e+09, 9.177618e+09, 9.351248e+09, 9.524738e+09, 
    9.697854e+09, 9.870353e+09, 1.004198e+10, 1.021247e+10, 1.038154e+10, 
    1.054891e+10, 1.071428e+10, 1.087735e+10, 1.10378e+10, 1.119532e+10, 
    1.134958e+10, 1.150025e+10, 1.164701e+10, 1.178951e+10, 1.192743e+10, 
    1.206044e+10, 1.218821e+10, 1.231041e+10, 1.242673e+10, 1.253687e+10, 
    1.264052e+10, 1.273739e+10, 1.282723e+10, 1.290977e+10, 1.298478e+10, 
    1.305203e+10, 1.311133e+10, 1.316249e+10, 1.320537e+10, 1.323984e+10, 
    1.326578e+10, 1.328312e+10, 1.32918e+10, 1.32918e+10, 1.328312e+10, 
    1.326578e+10, 1.323984e+10, 1.320537e+10, 1.316249e+10, 1.311133e+10, 
    1.305203e+10, 1.298478e+10, 1.290977e+10, 1.282723e+10, 1.273739e+10, 
    1.264052e+10, 1.253687e+10, 1.242673e+10, 1.231041e+10, 1.218821e+10, 
    1.206044e+10, 1.192743e+10, 1.178951e+10, 1.164701e+10, 1.150025e+10, 
    1.134958e+10, 1.119532e+10, 1.10378e+10, 1.087735e+10, 1.071428e+10, 
    1.054891e+10, 1.038154e+10, 1.021247e+10, 1.004198e+10, 9.870353e+09, 
    9.697854e+09, 9.524738e+09, 9.351248e+09, 9.177618e+09, 9.004068e+09, 
    8.830806e+09, 8.658028e+09, 8.485919e+09, 8.314652e+09, 8.144387e+09, 
    7.975273e+09, 7.807448e+09, 7.641037e+09, 7.476158e+09, 7.312915e+09, 
    7.151404e+09,
  7.155078e+09, 7.316969e+09, 7.480609e+09, 7.645901e+09, 7.812741e+09, 
    7.981012e+09, 8.150589e+09, 8.321333e+09, 8.493095e+09, 8.665715e+09, 
    8.839017e+09, 9.012821e+09, 9.186927e+09, 9.361125e+09, 9.535196e+09, 
    9.708905e+09, 9.882009e+09, 1.005425e+10, 1.022536e+10, 1.039506e+10, 
    1.056306e+10, 1.072907e+10, 1.089278e+10, 1.105388e+10, 1.121203e+10, 
    1.136693e+10, 1.151823e+10, 1.166561e+10, 1.180873e+10, 1.194726e+10, 
    1.208085e+10, 1.220919e+10, 1.233195e+10, 1.24488e+10, 1.255944e+10, 
    1.266358e+10, 1.276091e+10, 1.285118e+10, 1.293411e+10, 1.300948e+10, 
    1.307706e+10, 1.313664e+10, 1.318806e+10, 1.323115e+10, 1.326578e+10, 
    1.329185e+10, 1.330927e+10, 1.3318e+10, 1.3318e+10, 1.330927e+10, 
    1.329185e+10, 1.326578e+10, 1.323115e+10, 1.318806e+10, 1.313664e+10, 
    1.307706e+10, 1.300948e+10, 1.293411e+10, 1.285118e+10, 1.276091e+10, 
    1.266358e+10, 1.255944e+10, 1.24488e+10, 1.233195e+10, 1.220919e+10, 
    1.208085e+10, 1.194726e+10, 1.180873e+10, 1.166561e+10, 1.151823e+10, 
    1.136693e+10, 1.121203e+10, 1.105388e+10, 1.089278e+10, 1.072907e+10, 
    1.056306e+10, 1.039506e+10, 1.022536e+10, 1.005425e+10, 9.882009e+09, 
    9.708905e+09, 9.535196e+09, 9.361125e+09, 9.186927e+09, 9.012821e+09, 
    8.839017e+09, 8.665715e+09, 8.493095e+09, 8.321333e+09, 8.150589e+09, 
    7.981012e+09, 7.812741e+09, 7.645901e+09, 7.480609e+09, 7.316969e+09, 
    7.155078e+09,
  7.157529e+09, 7.319673e+09, 7.483577e+09, 7.649145e+09, 7.816271e+09, 
    7.984841e+09, 8.154726e+09, 8.32579e+09, 8.497883e+09, 8.670843e+09, 
    8.844498e+09, 9.018663e+09, 9.193139e+09, 9.367718e+09, 9.542177e+09, 
    9.716282e+09, 9.88979e+09, 1.006244e+10, 1.023397e+10, 1.040409e+10, 
    1.057252e+10, 1.073895e+10, 1.090309e+10, 1.106461e+10, 1.12232e+10, 
    1.137852e+10, 1.153025e+10, 1.167804e+10, 1.182158e+10, 1.19605e+10, 
    1.209449e+10, 1.222321e+10, 1.234634e+10, 1.246355e+10, 1.257453e+10, 
    1.267899e+10, 1.277663e+10, 1.286718e+10, 1.295038e+10, 1.302599e+10, 
    1.309378e+10, 1.315356e+10, 1.320514e+10, 1.324837e+10, 1.328312e+10, 
    1.330927e+10, 1.332675e+10, 1.333551e+10, 1.333551e+10, 1.332675e+10, 
    1.330927e+10, 1.328312e+10, 1.324837e+10, 1.320514e+10, 1.315356e+10, 
    1.309378e+10, 1.302599e+10, 1.295038e+10, 1.286718e+10, 1.277663e+10, 
    1.267899e+10, 1.257453e+10, 1.246355e+10, 1.234634e+10, 1.222321e+10, 
    1.209449e+10, 1.19605e+10, 1.182158e+10, 1.167804e+10, 1.153025e+10, 
    1.137852e+10, 1.12232e+10, 1.106461e+10, 1.090309e+10, 1.073895e+10, 
    1.057252e+10, 1.040409e+10, 1.023397e+10, 1.006244e+10, 9.88979e+09, 
    9.716282e+09, 9.542177e+09, 9.367718e+09, 9.193139e+09, 9.018663e+09, 
    8.844498e+09, 8.670843e+09, 8.497883e+09, 8.32579e+09, 8.154726e+09, 
    7.984841e+09, 7.816271e+09, 7.649145e+09, 7.483577e+09, 7.319673e+09, 
    7.157529e+09,
  7.158754e+09, 7.321026e+09, 7.485062e+09, 7.650767e+09, 7.818037e+09, 
    7.986756e+09, 8.156796e+09, 8.32802e+09, 8.500278e+09, 8.673409e+09, 
    8.84724e+09, 9.021585e+09, 9.196247e+09, 9.371016e+09, 9.54567e+09, 
    9.719975e+09, 9.893683e+09, 1.006654e+10, 1.023827e+10, 1.040861e+10, 
    1.057725e+10, 1.07439e+10, 1.090825e+10, 1.106999e+10, 1.122879e+10, 
    1.138432e+10, 1.153626e+10, 1.168427e+10, 1.1828e+10, 1.196713e+10, 
    1.210132e+10, 1.223023e+10, 1.235355e+10, 1.247093e+10, 1.258209e+10, 
    1.268671e+10, 1.27845e+10, 1.287519e+10, 1.295852e+10, 1.303425e+10, 
    1.310215e+10, 1.316203e+10, 1.32137e+10, 1.3257e+10, 1.32918e+10, 
    1.3318e+10, 1.333551e+10, 1.334428e+10, 1.334428e+10, 1.333551e+10, 
    1.3318e+10, 1.32918e+10, 1.3257e+10, 1.32137e+10, 1.316203e+10, 
    1.310215e+10, 1.303425e+10, 1.295852e+10, 1.287519e+10, 1.27845e+10, 
    1.268671e+10, 1.258209e+10, 1.247093e+10, 1.235355e+10, 1.223023e+10, 
    1.210132e+10, 1.196713e+10, 1.1828e+10, 1.168427e+10, 1.153626e+10, 
    1.138432e+10, 1.122879e+10, 1.106999e+10, 1.090825e+10, 1.07439e+10, 
    1.057725e+10, 1.040861e+10, 1.023827e+10, 1.006654e+10, 9.893683e+09, 
    9.719975e+09, 9.54567e+09, 9.371016e+09, 9.196247e+09, 9.021585e+09, 
    8.84724e+09, 8.673409e+09, 8.500278e+09, 8.32802e+09, 8.156796e+09, 
    7.986756e+09, 7.818037e+09, 7.650767e+09, 7.485062e+09, 7.321026e+09, 
    7.158754e+09,
  7.158754e+09, 7.321026e+09, 7.485062e+09, 7.650767e+09, 7.818037e+09, 
    7.986756e+09, 8.156796e+09, 8.32802e+09, 8.500278e+09, 8.673409e+09, 
    8.84724e+09, 9.021585e+09, 9.196247e+09, 9.371016e+09, 9.54567e+09, 
    9.719975e+09, 9.893683e+09, 1.006654e+10, 1.023827e+10, 1.040861e+10, 
    1.057725e+10, 1.07439e+10, 1.090825e+10, 1.106999e+10, 1.122879e+10, 
    1.138432e+10, 1.153626e+10, 1.168427e+10, 1.1828e+10, 1.196713e+10, 
    1.210132e+10, 1.223023e+10, 1.235355e+10, 1.247093e+10, 1.258209e+10, 
    1.268671e+10, 1.27845e+10, 1.287519e+10, 1.295852e+10, 1.303425e+10, 
    1.310215e+10, 1.316203e+10, 1.32137e+10, 1.3257e+10, 1.32918e+10, 
    1.3318e+10, 1.333551e+10, 1.334428e+10, 1.334428e+10, 1.333551e+10, 
    1.3318e+10, 1.32918e+10, 1.3257e+10, 1.32137e+10, 1.316203e+10, 
    1.310215e+10, 1.303425e+10, 1.295852e+10, 1.287519e+10, 1.27845e+10, 
    1.268671e+10, 1.258209e+10, 1.247093e+10, 1.235355e+10, 1.223023e+10, 
    1.210132e+10, 1.196713e+10, 1.1828e+10, 1.168427e+10, 1.153626e+10, 
    1.138432e+10, 1.122879e+10, 1.106999e+10, 1.090825e+10, 1.07439e+10, 
    1.057725e+10, 1.040861e+10, 1.023827e+10, 1.006654e+10, 9.893683e+09, 
    9.719975e+09, 9.54567e+09, 9.371016e+09, 9.196247e+09, 9.021585e+09, 
    8.84724e+09, 8.673409e+09, 8.500278e+09, 8.32802e+09, 8.156796e+09, 
    7.986756e+09, 7.818037e+09, 7.650767e+09, 7.485062e+09, 7.321026e+09, 
    7.158754e+09,
  7.157529e+09, 7.319673e+09, 7.483577e+09, 7.649145e+09, 7.816271e+09, 
    7.984841e+09, 8.154726e+09, 8.32579e+09, 8.497883e+09, 8.670843e+09, 
    8.844498e+09, 9.018663e+09, 9.193139e+09, 9.367718e+09, 9.542177e+09, 
    9.716282e+09, 9.88979e+09, 1.006244e+10, 1.023397e+10, 1.040409e+10, 
    1.057252e+10, 1.073895e+10, 1.090309e+10, 1.106461e+10, 1.12232e+10, 
    1.137852e+10, 1.153025e+10, 1.167804e+10, 1.182158e+10, 1.19605e+10, 
    1.209449e+10, 1.222321e+10, 1.234634e+10, 1.246355e+10, 1.257453e+10, 
    1.267899e+10, 1.277663e+10, 1.286718e+10, 1.295038e+10, 1.302599e+10, 
    1.309378e+10, 1.315356e+10, 1.320514e+10, 1.324837e+10, 1.328312e+10, 
    1.330927e+10, 1.332675e+10, 1.333551e+10, 1.333551e+10, 1.332675e+10, 
    1.330927e+10, 1.328312e+10, 1.324837e+10, 1.320514e+10, 1.315356e+10, 
    1.309378e+10, 1.302599e+10, 1.295038e+10, 1.286718e+10, 1.277663e+10, 
    1.267899e+10, 1.257453e+10, 1.246355e+10, 1.234634e+10, 1.222321e+10, 
    1.209449e+10, 1.19605e+10, 1.182158e+10, 1.167804e+10, 1.153025e+10, 
    1.137852e+10, 1.12232e+10, 1.106461e+10, 1.090309e+10, 1.073895e+10, 
    1.057252e+10, 1.040409e+10, 1.023397e+10, 1.006244e+10, 9.88979e+09, 
    9.716282e+09, 9.542177e+09, 9.367718e+09, 9.193139e+09, 9.018663e+09, 
    8.844498e+09, 8.670843e+09, 8.497883e+09, 8.32579e+09, 8.154726e+09, 
    7.984841e+09, 7.816271e+09, 7.649145e+09, 7.483577e+09, 7.319673e+09, 
    7.157529e+09,
  7.155078e+09, 7.316969e+09, 7.480609e+09, 7.645901e+09, 7.812741e+09, 
    7.981012e+09, 8.150589e+09, 8.321333e+09, 8.493095e+09, 8.665715e+09, 
    8.839017e+09, 9.012821e+09, 9.186927e+09, 9.361125e+09, 9.535196e+09, 
    9.708905e+09, 9.882009e+09, 1.005425e+10, 1.022536e+10, 1.039506e+10, 
    1.056306e+10, 1.072907e+10, 1.089278e+10, 1.105388e+10, 1.121203e+10, 
    1.136693e+10, 1.151823e+10, 1.166561e+10, 1.180873e+10, 1.194726e+10, 
    1.208085e+10, 1.220919e+10, 1.233195e+10, 1.24488e+10, 1.255944e+10, 
    1.266358e+10, 1.276091e+10, 1.285118e+10, 1.293411e+10, 1.300948e+10, 
    1.307706e+10, 1.313664e+10, 1.318806e+10, 1.323115e+10, 1.326578e+10, 
    1.329185e+10, 1.330927e+10, 1.3318e+10, 1.3318e+10, 1.330927e+10, 
    1.329185e+10, 1.326578e+10, 1.323115e+10, 1.318806e+10, 1.313664e+10, 
    1.307706e+10, 1.300948e+10, 1.293411e+10, 1.285118e+10, 1.276091e+10, 
    1.266358e+10, 1.255944e+10, 1.24488e+10, 1.233195e+10, 1.220919e+10, 
    1.208085e+10, 1.194726e+10, 1.180873e+10, 1.166561e+10, 1.151823e+10, 
    1.136693e+10, 1.121203e+10, 1.105388e+10, 1.089278e+10, 1.072907e+10, 
    1.056306e+10, 1.039506e+10, 1.022536e+10, 1.005425e+10, 9.882009e+09, 
    9.708905e+09, 9.535196e+09, 9.361125e+09, 9.186927e+09, 9.012821e+09, 
    8.839017e+09, 8.665715e+09, 8.493095e+09, 8.321333e+09, 8.150589e+09, 
    7.981012e+09, 7.812741e+09, 7.645901e+09, 7.480609e+09, 7.316969e+09, 
    7.155078e+09,
  7.151404e+09, 7.312915e+09, 7.476158e+09, 7.641037e+09, 7.807448e+09, 
    7.975273e+09, 8.144387e+09, 8.314652e+09, 8.485919e+09, 8.658028e+09, 
    8.830806e+09, 9.004068e+09, 9.177618e+09, 9.351248e+09, 9.524738e+09, 
    9.697854e+09, 9.870353e+09, 1.004198e+10, 1.021247e+10, 1.038154e+10, 
    1.054891e+10, 1.071428e+10, 1.087735e+10, 1.10378e+10, 1.119532e+10, 
    1.134958e+10, 1.150025e+10, 1.164701e+10, 1.178951e+10, 1.192743e+10, 
    1.206044e+10, 1.218821e+10, 1.231041e+10, 1.242673e+10, 1.253687e+10, 
    1.264052e+10, 1.273739e+10, 1.282723e+10, 1.290977e+10, 1.298478e+10, 
    1.305203e+10, 1.311133e+10, 1.316249e+10, 1.320537e+10, 1.323984e+10, 
    1.326578e+10, 1.328312e+10, 1.32918e+10, 1.32918e+10, 1.328312e+10, 
    1.326578e+10, 1.323984e+10, 1.320537e+10, 1.316249e+10, 1.311133e+10, 
    1.305203e+10, 1.298478e+10, 1.290977e+10, 1.282723e+10, 1.273739e+10, 
    1.264052e+10, 1.253687e+10, 1.242673e+10, 1.231041e+10, 1.218821e+10, 
    1.206044e+10, 1.192743e+10, 1.178951e+10, 1.164701e+10, 1.150025e+10, 
    1.134958e+10, 1.119532e+10, 1.10378e+10, 1.087735e+10, 1.071428e+10, 
    1.054891e+10, 1.038154e+10, 1.021247e+10, 1.004198e+10, 9.870353e+09, 
    9.697854e+09, 9.524738e+09, 9.351248e+09, 9.177618e+09, 9.004068e+09, 
    8.830806e+09, 8.658028e+09, 8.485919e+09, 8.314652e+09, 8.144387e+09, 
    7.975273e+09, 7.807448e+09, 7.641037e+09, 7.476158e+09, 7.312915e+09, 
    7.151404e+09,
  7.146505e+09, 7.307511e+09, 7.470226e+09, 7.634556e+09, 7.800395e+09, 
    7.967627e+09, 8.136126e+09, 8.305754e+09, 8.476363e+09, 8.647793e+09, 
    8.819871e+09, 8.992415e+09, 9.165227e+09, 9.338102e+09, 9.510819e+09, 
    9.683147e+09, 9.854844e+09, 1.002566e+10, 1.019532e+10, 1.036355e+10, 
    1.053008e+10, 1.06946e+10, 1.085682e+10, 1.101642e+10, 1.117309e+10, 
    1.13265e+10, 1.147634e+10, 1.162227e+10, 1.176396e+10, 1.190108e+10, 
    1.203331e+10, 1.216031e+10, 1.228178e+10, 1.23974e+10, 1.250686e+10, 
    1.260987e+10, 1.270614e+10, 1.279542e+10, 1.287743e+10, 1.295196e+10, 
    1.301878e+10, 1.30777e+10, 1.312854e+10, 1.317114e+10, 1.320537e+10, 
    1.323115e+10, 1.324837e+10, 1.3257e+10, 1.3257e+10, 1.324837e+10, 
    1.323115e+10, 1.320537e+10, 1.317114e+10, 1.312854e+10, 1.30777e+10, 
    1.301878e+10, 1.295196e+10, 1.287743e+10, 1.279542e+10, 1.270614e+10, 
    1.260987e+10, 1.250686e+10, 1.23974e+10, 1.228178e+10, 1.216031e+10, 
    1.203331e+10, 1.190108e+10, 1.176396e+10, 1.162227e+10, 1.147634e+10, 
    1.13265e+10, 1.117309e+10, 1.101642e+10, 1.085682e+10, 1.06946e+10, 
    1.053008e+10, 1.036355e+10, 1.019532e+10, 1.002566e+10, 9.854844e+09, 
    9.683147e+09, 9.510819e+09, 9.338102e+09, 9.165227e+09, 8.992415e+09, 
    8.819871e+09, 8.647793e+09, 8.476363e+09, 8.305754e+09, 8.136126e+09, 
    7.967627e+09, 7.800395e+09, 7.634556e+09, 7.470226e+09, 7.307511e+09, 
    7.146505e+09,
  7.140384e+09, 7.30076e+09, 7.462817e+09, 7.626462e+09, 7.791588e+09, 
    7.958081e+09, 8.125813e+09, 8.294647e+09, 8.464436e+09, 8.63502e+09, 
    8.806228e+09, 8.977876e+09, 9.14977e+09, 9.321703e+09, 9.49346e+09, 
    9.664807e+09, 9.835507e+09, 1.00053e+10, 1.017394e+10, 1.034114e+10, 
    1.050662e+10, 1.067009e+10, 1.083124e+10, 1.098979e+10, 1.11454e+10, 
    1.129776e+10, 1.144656e+10, 1.159146e+10, 1.173213e+10, 1.186826e+10, 
    1.199952e+10, 1.212559e+10, 1.224615e+10, 1.236089e+10, 1.246951e+10, 
    1.257172e+10, 1.266725e+10, 1.275582e+10, 1.283719e+10, 1.291113e+10, 
    1.297741e+10, 1.303585e+10, 1.308628e+10, 1.312854e+10, 1.316249e+10, 
    1.318806e+10, 1.320514e+10, 1.32137e+10, 1.32137e+10, 1.320514e+10, 
    1.318806e+10, 1.316249e+10, 1.312854e+10, 1.308628e+10, 1.303585e+10, 
    1.297741e+10, 1.291113e+10, 1.283719e+10, 1.275582e+10, 1.266725e+10, 
    1.257172e+10, 1.246951e+10, 1.236089e+10, 1.224615e+10, 1.212559e+10, 
    1.199952e+10, 1.186826e+10, 1.173213e+10, 1.159146e+10, 1.144656e+10, 
    1.129776e+10, 1.11454e+10, 1.098979e+10, 1.083124e+10, 1.067009e+10, 
    1.050662e+10, 1.034114e+10, 1.017394e+10, 1.00053e+10, 9.835507e+09, 
    9.664807e+09, 9.49346e+09, 9.321703e+09, 9.14977e+09, 8.977876e+09, 
    8.806228e+09, 8.63502e+09, 8.464436e+09, 8.294647e+09, 8.125813e+09, 
    7.958081e+09, 7.791588e+09, 7.626462e+09, 7.462817e+09, 7.30076e+09, 
    7.140384e+09,
  7.133041e+09, 7.292662e+09, 7.453934e+09, 7.616759e+09, 7.781033e+09, 
    7.946641e+09, 8.113456e+09, 8.281342e+09, 8.450151e+09, 8.619724e+09, 
    8.789891e+09, 8.96047e+09, 9.131267e+09, 9.302078e+09, 9.472687e+09, 
    9.642865e+09, 9.812372e+09, 9.980962e+09, 1.014837e+10, 1.031433e+10, 
    1.047856e+10, 1.064077e+10, 1.080067e+10, 1.095795e+10, 1.111231e+10, 
    1.126342e+10, 1.141097e+10, 1.155465e+10, 1.169412e+10, 1.182907e+10, 
    1.195917e+10, 1.208412e+10, 1.220359e+10, 1.231729e+10, 1.242492e+10, 
    1.252618e+10, 1.262082e+10, 1.270856e+10, 1.278916e+10, 1.286239e+10, 
    1.292804e+10, 1.298592e+10, 1.303585e+10, 1.30777e+10, 1.311133e+10, 
    1.313664e+10, 1.315356e+10, 1.316203e+10, 1.316203e+10, 1.315356e+10, 
    1.313664e+10, 1.311133e+10, 1.30777e+10, 1.303585e+10, 1.298592e+10, 
    1.292804e+10, 1.286239e+10, 1.278916e+10, 1.270856e+10, 1.262082e+10, 
    1.252618e+10, 1.242492e+10, 1.231729e+10, 1.220359e+10, 1.208412e+10, 
    1.195917e+10, 1.182907e+10, 1.169412e+10, 1.155465e+10, 1.141097e+10, 
    1.126342e+10, 1.111231e+10, 1.095795e+10, 1.080067e+10, 1.064077e+10, 
    1.047856e+10, 1.031433e+10, 1.014837e+10, 9.980962e+09, 9.812372e+09, 
    9.642865e+09, 9.472687e+09, 9.302078e+09, 9.131267e+09, 8.96047e+09, 
    8.789891e+09, 8.619724e+09, 8.450151e+09, 8.281342e+09, 8.113456e+09, 
    7.946641e+09, 7.781033e+09, 7.616759e+09, 7.453934e+09, 7.292662e+09, 
    7.133041e+09,
  7.124479e+09, 7.283223e+09, 7.443579e+09, 7.605452e+09, 7.768736e+09, 
    7.933316e+09, 8.099066e+09, 8.26585e+09, 8.433522e+09, 8.601922e+09, 
    8.770882e+09, 8.940219e+09, 9.109745e+09, 9.279254e+09, 9.448532e+09, 
    9.617354e+09, 9.785482e+09, 9.95267e+09, 1.011866e+10, 1.028319e+10, 
    1.044597e+10, 1.060673e+10, 1.076517e+10, 1.092099e+10, 1.107389e+10, 
    1.122356e+10, 1.136968e+10, 1.151193e+10, 1.165001e+10, 1.17836e+10, 
    1.191237e+10, 1.203602e+10, 1.215424e+10, 1.226673e+10, 1.237321e+10, 
    1.247338e+10, 1.256699e+10, 1.265377e+10, 1.273348e+10, 1.280589e+10, 
    1.287081e+10, 1.292804e+10, 1.297741e+10, 1.301878e+10, 1.305203e+10, 
    1.307706e+10, 1.309378e+10, 1.310215e+10, 1.310215e+10, 1.309378e+10, 
    1.307706e+10, 1.305203e+10, 1.301878e+10, 1.297741e+10, 1.292804e+10, 
    1.287081e+10, 1.280589e+10, 1.273348e+10, 1.265377e+10, 1.256699e+10, 
    1.247338e+10, 1.237321e+10, 1.226673e+10, 1.215424e+10, 1.203602e+10, 
    1.191237e+10, 1.17836e+10, 1.165001e+10, 1.151193e+10, 1.136968e+10, 
    1.122356e+10, 1.107389e+10, 1.092099e+10, 1.076517e+10, 1.060673e+10, 
    1.044597e+10, 1.028319e+10, 1.011866e+10, 9.95267e+09, 9.785482e+09, 
    9.617354e+09, 9.448532e+09, 9.279254e+09, 9.109745e+09, 8.940219e+09, 
    8.770882e+09, 8.601922e+09, 8.433522e+09, 8.26585e+09, 8.099066e+09, 
    7.933316e+09, 7.768736e+09, 7.605452e+09, 7.443579e+09, 7.283223e+09, 
    7.124479e+09,
  7.1147e+09, 7.272444e+09, 7.431758e+09, 7.592547e+09, 7.754704e+09, 
    7.918115e+09, 8.082655e+09, 8.248187e+09, 8.414565e+09, 8.581632e+09, 
    8.749221e+09, 8.917151e+09, 9.085231e+09, 9.253263e+09, 9.421031e+09, 
    9.588315e+09, 9.754878e+09, 9.920478e+09, 1.008486e+10, 1.024776e+10, 
    1.040891e+10, 1.056802e+10, 1.07248e+10, 1.087898e+10, 1.103023e+10, 
    1.117826e+10, 1.132276e+10, 1.146341e+10, 1.159992e+10, 1.173195e+10, 
    1.185922e+10, 1.198141e+10, 1.209821e+10, 1.220935e+10, 1.231452e+10, 
    1.241347e+10, 1.250591e+10, 1.25916e+10, 1.267031e+10, 1.27418e+10, 
    1.280589e+10, 1.286239e+10, 1.291113e+10, 1.295196e+10, 1.298478e+10, 
    1.300948e+10, 1.302599e+10, 1.303425e+10, 1.303425e+10, 1.302599e+10, 
    1.300948e+10, 1.298478e+10, 1.295196e+10, 1.291113e+10, 1.286239e+10, 
    1.280589e+10, 1.27418e+10, 1.267031e+10, 1.25916e+10, 1.250591e+10, 
    1.241347e+10, 1.231452e+10, 1.220935e+10, 1.209821e+10, 1.198141e+10, 
    1.185922e+10, 1.173195e+10, 1.159992e+10, 1.146341e+10, 1.132276e+10, 
    1.117826e+10, 1.103023e+10, 1.087898e+10, 1.07248e+10, 1.056802e+10, 
    1.040891e+10, 1.024776e+10, 1.008486e+10, 9.920478e+09, 9.754878e+09, 
    9.588315e+09, 9.421031e+09, 9.253263e+09, 9.085231e+09, 8.917151e+09, 
    8.749221e+09, 8.581632e+09, 8.414565e+09, 8.248187e+09, 8.082655e+09, 
    7.918115e+09, 7.754704e+09, 7.592547e+09, 7.431758e+09, 7.272444e+09, 
    7.1147e+09,
  7.103705e+09, 7.260329e+09, 7.418477e+09, 7.578052e+09, 7.738948e+09, 
    7.901051e+09, 8.064236e+09, 8.228367e+09, 8.3933e+09, 8.558878e+09, 
    8.724934e+09, 8.891291e+09, 9.05776e+09, 9.224142e+09, 9.390226e+09, 
    9.555794e+09, 9.720613e+09, 9.884442e+09, 1.004703e+10, 1.020812e+10, 
    1.036744e+10, 1.052472e+10, 1.067967e+10, 1.0832e+10, 1.098142e+10, 
    1.112763e+10, 1.127033e+10, 1.14092e+10, 1.154395e+10, 1.167428e+10, 
    1.179987e+10, 1.192043e+10, 1.203567e+10, 1.214529e+10, 1.224902e+10, 
    1.234659e+10, 1.243775e+10, 1.252223e+10, 1.259983e+10, 1.267031e+10, 
    1.273348e+10, 1.278916e+10, 1.283719e+10, 1.287743e+10, 1.290977e+10, 
    1.293411e+10, 1.295038e+10, 1.295852e+10, 1.295852e+10, 1.295038e+10, 
    1.293411e+10, 1.290977e+10, 1.287743e+10, 1.283719e+10, 1.278916e+10, 
    1.273348e+10, 1.267031e+10, 1.259983e+10, 1.252223e+10, 1.243775e+10, 
    1.234659e+10, 1.224902e+10, 1.214529e+10, 1.203567e+10, 1.192043e+10, 
    1.179987e+10, 1.167428e+10, 1.154395e+10, 1.14092e+10, 1.127033e+10, 
    1.112763e+10, 1.098142e+10, 1.0832e+10, 1.067967e+10, 1.052472e+10, 
    1.036744e+10, 1.020812e+10, 1.004703e+10, 9.884442e+09, 9.720613e+09, 
    9.555794e+09, 9.390226e+09, 9.224142e+09, 9.05776e+09, 8.891291e+09, 
    8.724934e+09, 8.558878e+09, 8.3933e+09, 8.228367e+09, 8.064236e+09, 
    7.901051e+09, 7.738948e+09, 7.578052e+09, 7.418477e+09, 7.260329e+09, 
    7.103705e+09,
  7.091497e+09, 7.246883e+09, 7.403741e+09, 7.561974e+09, 7.721477e+09, 
    7.882135e+09, 8.043825e+09, 8.20641e+09, 8.369748e+09, 8.533684e+09, 
    8.698051e+09, 8.862674e+09, 9.027367e+09, 9.191932e+09, 9.356163e+09, 
    9.519842e+09, 9.68274e+09, 9.844622e+09, 1.000524e+10, 1.016434e+10, 
    1.032166e+10, 1.047692e+10, 1.062985e+10, 1.078017e+10, 1.092757e+10, 
    1.107179e+10, 1.12125e+10, 1.134943e+10, 1.148226e+10, 1.16107e+10, 
    1.173446e+10, 1.185324e+10, 1.196675e+10, 1.207473e+10, 1.217688e+10, 
    1.227295e+10, 1.236269e+10, 1.244586e+10, 1.252223e+10, 1.25916e+10, 
    1.265377e+10, 1.270856e+10, 1.275582e+10, 1.279542e+10, 1.282723e+10, 
    1.285118e+10, 1.286718e+10, 1.287519e+10, 1.287519e+10, 1.286718e+10, 
    1.285118e+10, 1.282723e+10, 1.279542e+10, 1.275582e+10, 1.270856e+10, 
    1.265377e+10, 1.25916e+10, 1.252223e+10, 1.244586e+10, 1.236269e+10, 
    1.227295e+10, 1.217688e+10, 1.207473e+10, 1.196675e+10, 1.185324e+10, 
    1.173446e+10, 1.16107e+10, 1.148226e+10, 1.134943e+10, 1.12125e+10, 
    1.107179e+10, 1.092757e+10, 1.078017e+10, 1.062985e+10, 1.047692e+10, 
    1.032166e+10, 1.016434e+10, 1.000524e+10, 9.844622e+09, 9.68274e+09, 
    9.519842e+09, 9.356163e+09, 9.191932e+09, 9.027367e+09, 8.862674e+09, 
    8.698051e+09, 8.533684e+09, 8.369748e+09, 8.20641e+09, 8.043825e+09, 
    7.882135e+09, 7.721477e+09, 7.561974e+09, 7.403741e+09, 7.246883e+09, 
    7.091497e+09,
  7.078078e+09, 7.23211e+09, 7.387556e+09, 7.544322e+09, 7.702302e+09, 
    7.861382e+09, 8.021437e+09, 8.182336e+09, 8.343933e+09, 8.506077e+09, 
    8.668601e+09, 8.831335e+09, 8.994092e+09, 9.156679e+09, 9.318892e+09, 
    9.480515e+09, 9.641325e+09, 9.801088e+09, 9.959563e+09, 1.01165e+10, 
    1.027164e+10, 1.042471e+10, 1.057545e+10, 1.072358e+10, 1.08688e+10, 
    1.101085e+10, 1.114942e+10, 1.128423e+10, 1.141498e+10, 1.154138e+10, 
    1.166315e+10, 1.178001e+10, 1.189166e+10, 1.199784e+10, 1.209829e+10, 
    1.219274e+10, 1.228095e+10, 1.236269e+10, 1.243775e+10, 1.250591e+10, 
    1.256699e+10, 1.262082e+10, 1.266725e+10, 1.270614e+10, 1.273739e+10, 
    1.276091e+10, 1.277663e+10, 1.27845e+10, 1.27845e+10, 1.277663e+10, 
    1.276091e+10, 1.273739e+10, 1.270614e+10, 1.266725e+10, 1.262082e+10, 
    1.256699e+10, 1.250591e+10, 1.243775e+10, 1.236269e+10, 1.228095e+10, 
    1.219274e+10, 1.209829e+10, 1.199784e+10, 1.189166e+10, 1.178001e+10, 
    1.166315e+10, 1.154138e+10, 1.141498e+10, 1.128423e+10, 1.114942e+10, 
    1.101085e+10, 1.08688e+10, 1.072358e+10, 1.057545e+10, 1.042471e+10, 
    1.027164e+10, 1.01165e+10, 9.959563e+09, 9.801088e+09, 9.641325e+09, 
    9.480515e+09, 9.318892e+09, 9.156679e+09, 8.994092e+09, 8.831335e+09, 
    8.668601e+09, 8.506077e+09, 8.343933e+09, 8.182336e+09, 8.021437e+09, 
    7.861382e+09, 7.702302e+09, 7.544322e+09, 7.387556e+09, 7.23211e+09, 
    7.078078e+09,
  7.063453e+09, 7.216014e+09, 7.36993e+09, 7.525106e+09, 7.681435e+09, 
    7.838806e+09, 7.997093e+09, 8.156166e+09, 8.31588e+09, 8.476086e+09, 
    8.636621e+09, 8.797313e+09, 8.95798e+09, 9.118431e+09, 9.278465e+09, 
    9.437871e+09, 9.596429e+09, 9.753911e+09, 9.910078e+09, 1.006469e+10, 
    1.021748e+10, 1.03682e+10, 1.051658e+10, 1.066235e+10, 1.080523e+10, 
    1.094495e+10, 1.108122e+10, 1.121375e+10, 1.134227e+10, 1.146649e+10, 
    1.158613e+10, 1.170091e+10, 1.181057e+10, 1.191483e+10, 1.201345e+10, 
    1.210616e+10, 1.219274e+10, 1.227295e+10, 1.234659e+10, 1.241347e+10, 
    1.247338e+10, 1.252618e+10, 1.257172e+10, 1.260987e+10, 1.264052e+10, 
    1.266358e+10, 1.267899e+10, 1.268671e+10, 1.268671e+10, 1.267899e+10, 
    1.266358e+10, 1.264052e+10, 1.260987e+10, 1.257172e+10, 1.252618e+10, 
    1.247338e+10, 1.241347e+10, 1.234659e+10, 1.227295e+10, 1.219274e+10, 
    1.210616e+10, 1.201345e+10, 1.191483e+10, 1.181057e+10, 1.170091e+10, 
    1.158613e+10, 1.146649e+10, 1.134227e+10, 1.121375e+10, 1.108122e+10, 
    1.094495e+10, 1.080523e+10, 1.066235e+10, 1.051658e+10, 1.03682e+10, 
    1.021748e+10, 1.006469e+10, 9.910078e+09, 9.753911e+09, 9.596429e+09, 
    9.437871e+09, 9.278465e+09, 9.118431e+09, 8.95798e+09, 8.797313e+09, 
    8.636621e+09, 8.476086e+09, 8.31588e+09, 8.156166e+09, 7.997093e+09, 
    7.838806e+09, 7.681435e+09, 7.525106e+09, 7.36993e+09, 7.216014e+09, 
    7.063453e+09,
  7.047623e+09, 7.198601e+09, 7.350871e+09, 7.504335e+09, 7.65889e+09, 
    7.814423e+09, 7.970811e+09, 8.127923e+09, 8.285618e+09, 8.443745e+09, 
    8.602145e+09, 8.760649e+09, 8.919077e+09, 9.077242e+09, 9.234944e+09, 
    9.391978e+09, 9.548129e+09, 9.703171e+09, 9.856871e+09, 1.000899e+10, 
    1.015928e+10, 1.030749e+10, 1.045336e+10, 1.059662e+10, 1.0737e+10, 
    1.087423e+10, 1.100805e+10, 1.113816e+10, 1.12643e+10, 1.13862e+10, 
    1.150357e+10, 1.161615e+10, 1.172369e+10, 1.182591e+10, 1.192258e+10, 
    1.201345e+10, 1.209829e+10, 1.217688e+10, 1.224902e+10, 1.231452e+10, 
    1.237321e+10, 1.242492e+10, 1.246951e+10, 1.250686e+10, 1.253687e+10, 
    1.255944e+10, 1.257453e+10, 1.258209e+10, 1.258209e+10, 1.257453e+10, 
    1.255944e+10, 1.253687e+10, 1.250686e+10, 1.246951e+10, 1.242492e+10, 
    1.237321e+10, 1.231452e+10, 1.224902e+10, 1.217688e+10, 1.209829e+10, 
    1.201345e+10, 1.192258e+10, 1.182591e+10, 1.172369e+10, 1.161615e+10, 
    1.150357e+10, 1.13862e+10, 1.12643e+10, 1.113816e+10, 1.100805e+10, 
    1.087423e+10, 1.0737e+10, 1.059662e+10, 1.045336e+10, 1.030749e+10, 
    1.015928e+10, 1.000899e+10, 9.856871e+09, 9.703171e+09, 9.548129e+09, 
    9.391978e+09, 9.234944e+09, 9.077242e+09, 8.919077e+09, 8.760649e+09, 
    8.602145e+09, 8.443745e+09, 8.285618e+09, 8.127923e+09, 7.970811e+09, 
    7.814423e+09, 7.65889e+09, 7.504335e+09, 7.350871e+09, 7.198601e+09, 
    7.047623e+09,
  7.030593e+09, 7.179877e+09, 7.330385e+09, 7.482021e+09, 7.634681e+09, 
    7.788252e+09, 7.942612e+09, 8.097633e+09, 8.253174e+09, 8.409087e+09, 
    8.565214e+09, 8.721389e+09, 8.877434e+09, 9.033167e+09, 9.188391e+09, 
    9.342905e+09, 9.496498e+09, 9.64895e+09, 9.800034e+09, 9.949515e+09, 
    1.009715e+10, 1.02427e+10, 1.03859e+10, 1.05265e+10, 1.066424e+10, 
    1.079885e+10, 1.093007e+10, 1.105763e+10, 1.118125e+10, 1.130069e+10, 
    1.141567e+10, 1.152593e+10, 1.163122e+10, 1.17313e+10, 1.182591e+10, 
    1.191483e+10, 1.199784e+10, 1.207473e+10, 1.214529e+10, 1.220935e+10, 
    1.226673e+10, 1.231729e+10, 1.236089e+10, 1.23974e+10, 1.242673e+10, 
    1.24488e+10, 1.246355e+10, 1.247093e+10, 1.247093e+10, 1.246355e+10, 
    1.24488e+10, 1.242673e+10, 1.23974e+10, 1.236089e+10, 1.231729e+10, 
    1.226673e+10, 1.220935e+10, 1.214529e+10, 1.207473e+10, 1.199784e+10, 
    1.191483e+10, 1.182591e+10, 1.17313e+10, 1.163122e+10, 1.152593e+10, 
    1.141567e+10, 1.130069e+10, 1.118125e+10, 1.105763e+10, 1.093007e+10, 
    1.079885e+10, 1.066424e+10, 1.05265e+10, 1.03859e+10, 1.02427e+10, 
    1.009715e+10, 9.949515e+09, 9.800034e+09, 9.64895e+09, 9.496498e+09, 
    9.342905e+09, 9.188391e+09, 9.033167e+09, 8.877434e+09, 8.721389e+09, 
    8.565214e+09, 8.409087e+09, 8.253174e+09, 8.097633e+09, 7.942612e+09, 
    7.788252e+09, 7.634681e+09, 7.482021e+09, 7.330385e+09, 7.179877e+09, 
    7.030593e+09,
  7.012366e+09, 7.159848e+09, 7.308484e+09, 7.458176e+09, 7.608822e+09, 
    7.760311e+09, 7.912521e+09, 8.065324e+09, 8.218582e+09, 8.372148e+09, 
    8.525868e+09, 8.679578e+09, 8.833104e+09, 8.986266e+09, 9.138871e+09, 
    9.290724e+09, 9.441618e+09, 9.591338e+09, 9.739662e+09, 9.886363e+09, 
    1.00312e+10, 1.017395e+10, 1.031435e+10, 1.045215e+10, 1.058711e+10, 
    1.071896e+10, 1.084745e+10, 1.097232e+10, 1.109331e+10, 1.121017e+10, 
    1.132264e+10, 1.143046e+10, 1.153341e+10, 1.163122e+10, 1.172369e+10, 
    1.181057e+10, 1.189166e+10, 1.196675e+10, 1.203567e+10, 1.209821e+10, 
    1.215424e+10, 1.220359e+10, 1.224615e+10, 1.228178e+10, 1.231041e+10, 
    1.233195e+10, 1.234634e+10, 1.235355e+10, 1.235355e+10, 1.234634e+10, 
    1.233195e+10, 1.231041e+10, 1.228178e+10, 1.224615e+10, 1.220359e+10, 
    1.215424e+10, 1.209821e+10, 1.203567e+10, 1.196675e+10, 1.189166e+10, 
    1.181057e+10, 1.172369e+10, 1.163122e+10, 1.153341e+10, 1.143046e+10, 
    1.132264e+10, 1.121017e+10, 1.109331e+10, 1.097232e+10, 1.084745e+10, 
    1.071896e+10, 1.058711e+10, 1.045215e+10, 1.031435e+10, 1.017395e+10, 
    1.00312e+10, 9.886363e+09, 9.739662e+09, 9.591338e+09, 9.441618e+09, 
    9.290724e+09, 9.138871e+09, 8.986266e+09, 8.833104e+09, 8.679578e+09, 
    8.525868e+09, 8.372148e+09, 8.218582e+09, 8.065324e+09, 7.912521e+09, 
    7.760311e+09, 7.608822e+09, 7.458176e+09, 7.308484e+09, 7.159848e+09, 
    7.012366e+09,
  6.992947e+09, 7.138521e+09, 7.285175e+09, 7.432813e+09, 7.581331e+09, 
    7.73062e+09, 7.880559e+09, 8.031022e+09, 8.181873e+09, 8.332967e+09, 
    8.484152e+09, 8.635267e+09, 8.786142e+09, 8.936601e+09, 9.086456e+09, 
    9.235513e+09, 9.383574e+09, 9.530426e+09, 9.675857e+09, 9.819643e+09, 
    9.961556e+09, 1.010136e+10, 1.023883e+10, 1.037371e+10, 1.050575e+10, 
    1.063472e+10, 1.076036e+10, 1.088243e+10, 1.100067e+10, 1.111483e+10, 
    1.122468e+10, 1.132997e+10, 1.143046e+10, 1.152593e+10, 1.161615e+10, 
    1.170091e+10, 1.178001e+10, 1.185324e+10, 1.192043e+10, 1.198141e+10, 
    1.203602e+10, 1.208412e+10, 1.212559e+10, 1.216031e+10, 1.218821e+10, 
    1.220919e+10, 1.222321e+10, 1.223023e+10, 1.223023e+10, 1.222321e+10, 
    1.220919e+10, 1.218821e+10, 1.216031e+10, 1.212559e+10, 1.208412e+10, 
    1.203602e+10, 1.198141e+10, 1.192043e+10, 1.185324e+10, 1.178001e+10, 
    1.170091e+10, 1.161615e+10, 1.152593e+10, 1.143046e+10, 1.132997e+10, 
    1.122468e+10, 1.111483e+10, 1.100067e+10, 1.088243e+10, 1.076036e+10, 
    1.063472e+10, 1.050575e+10, 1.037371e+10, 1.023883e+10, 1.010136e+10, 
    9.961556e+09, 9.819643e+09, 9.675857e+09, 9.530426e+09, 9.383574e+09, 
    9.235513e+09, 9.086456e+09, 8.936601e+09, 8.786142e+09, 8.635267e+09, 
    8.484152e+09, 8.332967e+09, 8.181873e+09, 8.031022e+09, 7.880559e+09, 
    7.73062e+09, 7.581331e+09, 7.432813e+09, 7.285175e+09, 7.138521e+09, 
    6.992947e+09,
  6.972339e+09, 7.115902e+09, 7.260469e+09, 7.405943e+09, 7.552224e+09, 
    7.699199e+09, 7.846753e+09, 7.994759e+09, 8.143084e+09, 8.291585e+09, 
    8.440113e+09, 8.58851e+09, 8.736609e+09, 8.884238e+09, 9.031216e+09, 
    9.177352e+09, 9.322452e+09, 9.466312e+09, 9.608722e+09, 9.749469e+09, 
    9.88833e+09, 1.002508e+10, 1.015949e+10, 1.029132e+10, 1.042034e+10, 
    1.054631e+10, 1.066899e+10, 1.078814e+10, 1.090352e+10, 1.10149e+10, 
    1.112203e+10, 1.122468e+10, 1.132264e+10, 1.141567e+10, 1.150357e+10, 
    1.158613e+10, 1.166315e+10, 1.173446e+10, 1.179987e+10, 1.185922e+10, 
    1.191237e+10, 1.195917e+10, 1.199952e+10, 1.203331e+10, 1.206044e+10, 
    1.208085e+10, 1.209449e+10, 1.210132e+10, 1.210132e+10, 1.209449e+10, 
    1.208085e+10, 1.206044e+10, 1.203331e+10, 1.199952e+10, 1.195917e+10, 
    1.191237e+10, 1.185922e+10, 1.179987e+10, 1.173446e+10, 1.166315e+10, 
    1.158613e+10, 1.150357e+10, 1.141567e+10, 1.132264e+10, 1.122468e+10, 
    1.112203e+10, 1.10149e+10, 1.090352e+10, 1.078814e+10, 1.066899e+10, 
    1.054631e+10, 1.042034e+10, 1.029132e+10, 1.015949e+10, 1.002508e+10, 
    9.88833e+09, 9.749469e+09, 9.608722e+09, 9.466312e+09, 9.322452e+09, 
    9.177352e+09, 9.031216e+09, 8.884238e+09, 8.736609e+09, 8.58851e+09, 
    8.440113e+09, 8.291585e+09, 8.143084e+09, 7.994759e+09, 7.846753e+09, 
    7.699199e+09, 7.552224e+09, 7.405943e+09, 7.260469e+09, 7.115902e+09, 
    6.972339e+09,
  6.950547e+09, 7.092e+09, 7.234377e+09, 7.377583e+09, 7.521518e+09, 
    7.666072e+09, 7.811129e+09, 7.956566e+09, 8.10225e+09, 8.248043e+09, 
    8.393798e+09, 8.539359e+09, 8.684566e+09, 8.829247e+09, 8.973229e+09, 
    9.116325e+09, 9.258346e+09, 9.399095e+09, 9.53837e+09, 9.67596e+09, 
    9.811654e+09, 9.945231e+09, 1.007647e+10, 1.020515e+10, 1.033104e+10, 
    1.045391e+10, 1.057352e+10, 1.068966e+10, 1.080209e+10, 1.091057e+10, 
    1.10149e+10, 1.111483e+10, 1.121017e+10, 1.130069e+10, 1.13862e+10, 
    1.146649e+10, 1.154138e+10, 1.16107e+10, 1.167428e+10, 1.173195e+10, 
    1.17836e+10, 1.182907e+10, 1.186826e+10, 1.190108e+10, 1.192743e+10, 
    1.194726e+10, 1.19605e+10, 1.196713e+10, 1.196713e+10, 1.19605e+10, 
    1.194726e+10, 1.192743e+10, 1.190108e+10, 1.186826e+10, 1.182907e+10, 
    1.17836e+10, 1.173195e+10, 1.167428e+10, 1.16107e+10, 1.154138e+10, 
    1.146649e+10, 1.13862e+10, 1.130069e+10, 1.121017e+10, 1.111483e+10, 
    1.10149e+10, 1.091057e+10, 1.080209e+10, 1.068966e+10, 1.057352e+10, 
    1.045391e+10, 1.033104e+10, 1.020515e+10, 1.007647e+10, 9.945231e+09, 
    9.811654e+09, 9.67596e+09, 9.53837e+09, 9.399095e+09, 9.258346e+09, 
    9.116325e+09, 8.973229e+09, 8.829247e+09, 8.684566e+09, 8.539359e+09, 
    8.393798e+09, 8.248043e+09, 8.10225e+09, 7.956566e+09, 7.811129e+09, 
    7.666072e+09, 7.521518e+09, 7.377583e+09, 7.234377e+09, 7.092e+09, 
    6.950547e+09,
  6.927576e+09, 7.066821e+09, 7.206909e+09, 7.347746e+09, 7.489233e+09, 
    7.631261e+09, 7.773715e+09, 7.916475e+09, 8.059411e+09, 8.202386e+09, 
    8.345257e+09, 8.487873e+09, 8.630074e+09, 8.771699e+09, 8.912572e+09, 
    9.052518e+09, 9.191351e+09, 9.32888e+09, 9.464909e+09, 9.599237e+09, 
    9.731658e+09, 9.861961e+09, 9.989933e+09, 1.011536e+10, 1.023802e+10, 
    1.035769e+10, 1.047415e+10, 1.058718e+10, 1.069657e+10, 1.080209e+10, 
    1.090352e+10, 1.100067e+10, 1.109331e+10, 1.118125e+10, 1.12643e+10, 
    1.134227e+10, 1.141498e+10, 1.148226e+10, 1.154395e+10, 1.159992e+10, 
    1.165001e+10, 1.169412e+10, 1.173213e+10, 1.176396e+10, 1.178951e+10, 
    1.180873e+10, 1.182158e+10, 1.1828e+10, 1.1828e+10, 1.182158e+10, 
    1.180873e+10, 1.178951e+10, 1.176396e+10, 1.173213e+10, 1.169412e+10, 
    1.165001e+10, 1.159992e+10, 1.154395e+10, 1.148226e+10, 1.141498e+10, 
    1.134227e+10, 1.12643e+10, 1.118125e+10, 1.109331e+10, 1.100067e+10, 
    1.090352e+10, 1.080209e+10, 1.069657e+10, 1.058718e+10, 1.047415e+10, 
    1.035769e+10, 1.023802e+10, 1.011536e+10, 9.989933e+09, 9.861961e+09, 
    9.731658e+09, 9.599237e+09, 9.464909e+09, 9.32888e+09, 9.191351e+09, 
    9.052518e+09, 8.912572e+09, 8.771699e+09, 8.630074e+09, 8.487873e+09, 
    8.345257e+09, 8.202386e+09, 8.059411e+09, 7.916475e+09, 7.773715e+09, 
    7.631261e+09, 7.489233e+09, 7.347746e+09, 7.206909e+09, 7.066821e+09, 
    6.927576e+09,
  6.903431e+09, 7.040374e+09, 7.178077e+09, 7.316448e+09, 7.455388e+09, 
    7.594789e+09, 7.734541e+09, 7.874522e+09, 8.014606e+09, 8.15466e+09, 
    8.294543e+09, 8.434108e+09, 8.573202e+09, 8.711665e+09, 8.849328e+09, 
    8.986021e+09, 9.121564e+09, 9.255772e+09, 9.388457e+09, 9.519426e+09, 
    9.648477e+09, 9.775411e+09, 9.900023e+09, 1.00221e+10, 1.014144e+10, 
    1.025783e+10, 1.037106e+10, 1.048091e+10, 1.058718e+10, 1.068966e+10, 
    1.078814e+10, 1.088243e+10, 1.097232e+10, 1.105763e+10, 1.113816e+10, 
    1.121375e+10, 1.128423e+10, 1.134943e+10, 1.14092e+10, 1.146341e+10, 
    1.151193e+10, 1.155465e+10, 1.159146e+10, 1.162227e+10, 1.164701e+10, 
    1.166561e+10, 1.167804e+10, 1.168427e+10, 1.168427e+10, 1.167804e+10, 
    1.166561e+10, 1.164701e+10, 1.162227e+10, 1.159146e+10, 1.155465e+10, 
    1.151193e+10, 1.146341e+10, 1.14092e+10, 1.134943e+10, 1.128423e+10, 
    1.121375e+10, 1.113816e+10, 1.105763e+10, 1.097232e+10, 1.088243e+10, 
    1.078814e+10, 1.068966e+10, 1.058718e+10, 1.048091e+10, 1.037106e+10, 
    1.025783e+10, 1.014144e+10, 1.00221e+10, 9.900023e+09, 9.775411e+09, 
    9.648477e+09, 9.519426e+09, 9.388457e+09, 9.255772e+09, 9.121564e+09, 
    8.986021e+09, 8.849328e+09, 8.711665e+09, 8.573202e+09, 8.434108e+09, 
    8.294543e+09, 8.15466e+09, 8.014606e+09, 7.874522e+09, 7.734541e+09, 
    7.594789e+09, 7.455388e+09, 7.316448e+09, 7.178077e+09, 7.040374e+09, 
    6.903431e+09,
  6.878117e+09, 7.012667e+09, 7.147894e+09, 7.283705e+09, 7.420003e+09, 
    7.556683e+09, 7.693634e+09, 7.830739e+09, 7.967875e+09, 8.10491e+09, 
    8.241709e+09, 8.378128e+09, 8.514017e+09, 8.649221e+09, 8.78358e+09, 
    8.916924e+09, 9.049084e+09, 9.17988e+09, 9.309132e+09, 9.436652e+09, 
    9.562249e+09, 9.68573e+09, 9.806899e+09, 9.925557e+09, 1.00415e+10, 
    1.015454e+10, 1.026446e+10, 1.037106e+10, 1.047415e+10, 1.057352e+10, 
    1.066899e+10, 1.076036e+10, 1.084745e+10, 1.093007e+10, 1.100805e+10, 
    1.108122e+10, 1.114942e+10, 1.12125e+10, 1.127033e+10, 1.132276e+10, 
    1.136968e+10, 1.141097e+10, 1.144656e+10, 1.147634e+10, 1.150025e+10, 
    1.151823e+10, 1.153025e+10, 1.153626e+10, 1.153626e+10, 1.153025e+10, 
    1.151823e+10, 1.150025e+10, 1.147634e+10, 1.144656e+10, 1.141097e+10, 
    1.136968e+10, 1.132276e+10, 1.127033e+10, 1.12125e+10, 1.114942e+10, 
    1.108122e+10, 1.100805e+10, 1.093007e+10, 1.084745e+10, 1.076036e+10, 
    1.066899e+10, 1.057352e+10, 1.047415e+10, 1.037106e+10, 1.026446e+10, 
    1.015454e+10, 1.00415e+10, 9.925557e+09, 9.806899e+09, 9.68573e+09, 
    9.562249e+09, 9.436652e+09, 9.309132e+09, 9.17988e+09, 9.049084e+09, 
    8.916924e+09, 8.78358e+09, 8.649221e+09, 8.514017e+09, 8.378128e+09, 
    8.241709e+09, 8.10491e+09, 7.967875e+09, 7.830739e+09, 7.693634e+09, 
    7.556683e+09, 7.420003e+09, 7.283705e+09, 7.147894e+09, 7.012667e+09, 
    6.878117e+09,
  6.851641e+09, 6.98371e+09, 7.116371e+09, 7.249533e+09, 7.383099e+09, 
    7.516966e+09, 7.651027e+09, 7.785166e+09, 7.919261e+09, 8.053188e+09, 
    8.186811e+09, 8.319992e+09, 8.452588e+09, 8.584445e+09, 8.715411e+09, 
    8.845323e+09, 8.974015e+09, 9.101317e+09, 9.227054e+09, 9.351046e+09, 
    9.473112e+09, 9.593066e+09, 9.710721e+09, 9.825887e+09, 9.938373e+09, 
    1.004799e+10, 1.015454e+10, 1.025783e+10, 1.035769e+10, 1.045391e+10, 
    1.054631e+10, 1.063472e+10, 1.071896e+10, 1.079885e+10, 1.087423e+10, 
    1.094495e+10, 1.101085e+10, 1.107179e+10, 1.112763e+10, 1.117826e+10, 
    1.122356e+10, 1.126342e+10, 1.129776e+10, 1.13265e+10, 1.134958e+10, 
    1.136693e+10, 1.137852e+10, 1.138432e+10, 1.138432e+10, 1.137852e+10, 
    1.136693e+10, 1.134958e+10, 1.13265e+10, 1.129776e+10, 1.126342e+10, 
    1.122356e+10, 1.117826e+10, 1.112763e+10, 1.107179e+10, 1.101085e+10, 
    1.094495e+10, 1.087423e+10, 1.079885e+10, 1.071896e+10, 1.063472e+10, 
    1.054631e+10, 1.045391e+10, 1.035769e+10, 1.025783e+10, 1.015454e+10, 
    1.004799e+10, 9.938373e+09, 9.825887e+09, 9.710721e+09, 9.593066e+09, 
    9.473112e+09, 9.351046e+09, 9.227054e+09, 9.101317e+09, 8.974015e+09, 
    8.845323e+09, 8.715411e+09, 8.584445e+09, 8.452588e+09, 8.319992e+09, 
    8.186811e+09, 8.053188e+09, 7.919261e+09, 7.785166e+09, 7.651027e+09, 
    7.516966e+09, 7.383099e+09, 7.249533e+09, 7.116371e+09, 6.98371e+09, 
    6.851641e+09,
  6.824007e+09, 6.953512e+09, 7.083523e+09, 7.21395e+09, 7.344698e+09, 
    7.475667e+09, 7.606751e+09, 7.737838e+09, 7.868808e+09, 7.99954e+09, 
    8.129904e+09, 8.259766e+09, 8.388985e+09, 8.517416e+09, 8.64491e+09, 
    8.771312e+09, 8.896461e+09, 9.020195e+09, 9.142345e+09, 9.262742e+09, 
    9.381209e+09, 9.497571e+09, 9.61165e+09, 9.723264e+09, 9.832232e+09, 
    9.938373e+09, 1.00415e+10, 1.014144e+10, 1.023802e+10, 1.033104e+10, 
    1.042034e+10, 1.050575e+10, 1.058711e+10, 1.066424e+10, 1.0737e+10, 
    1.080523e+10, 1.08688e+10, 1.092757e+10, 1.098142e+10, 1.103023e+10, 
    1.107389e+10, 1.111231e+10, 1.11454e+10, 1.117309e+10, 1.119532e+10, 
    1.121203e+10, 1.12232e+10, 1.122879e+10, 1.122879e+10, 1.12232e+10, 
    1.121203e+10, 1.119532e+10, 1.117309e+10, 1.11454e+10, 1.111231e+10, 
    1.107389e+10, 1.103023e+10, 1.098142e+10, 1.092757e+10, 1.08688e+10, 
    1.080523e+10, 1.0737e+10, 1.066424e+10, 1.058711e+10, 1.050575e+10, 
    1.042034e+10, 1.033104e+10, 1.023802e+10, 1.014144e+10, 1.00415e+10, 
    9.938373e+09, 9.832232e+09, 9.723264e+09, 9.61165e+09, 9.497571e+09, 
    9.381209e+09, 9.262742e+09, 9.142345e+09, 9.020195e+09, 8.896461e+09, 
    8.771312e+09, 8.64491e+09, 8.517416e+09, 8.388985e+09, 8.259766e+09, 
    8.129904e+09, 7.99954e+09, 7.868808e+09, 7.737838e+09, 7.606751e+09, 
    7.475667e+09, 7.344698e+09, 7.21395e+09, 7.083523e+09, 6.953512e+09, 
    6.824007e+09,
  6.795221e+09, 6.922081e+09, 7.049361e+09, 7.176973e+09, 7.304823e+09, 
    7.432814e+09, 7.56084e+09, 7.688794e+09, 7.816561e+09, 7.94402e+09, 
    8.071048e+09, 8.197513e+09, 8.323282e+09, 8.448214e+09, 8.572165e+09, 
    8.694987e+09, 8.816526e+09, 8.936627e+09, 9.055129e+09, 9.171869e+09, 
    9.286681e+09, 9.399396e+09, 9.509846e+09, 9.61786e+09, 9.723264e+09, 
    9.825887e+09, 9.925557e+09, 1.00221e+10, 1.011536e+10, 1.020515e+10, 
    1.029132e+10, 1.037371e+10, 1.045215e+10, 1.05265e+10, 1.059662e+10, 
    1.066235e+10, 1.072358e+10, 1.078017e+10, 1.0832e+10, 1.087898e+10, 
    1.092099e+10, 1.095795e+10, 1.098979e+10, 1.101642e+10, 1.10378e+10, 
    1.105388e+10, 1.106461e+10, 1.106999e+10, 1.106999e+10, 1.106461e+10, 
    1.105388e+10, 1.10378e+10, 1.101642e+10, 1.098979e+10, 1.095795e+10, 
    1.092099e+10, 1.087898e+10, 1.0832e+10, 1.078017e+10, 1.072358e+10, 
    1.066235e+10, 1.059662e+10, 1.05265e+10, 1.045215e+10, 1.037371e+10, 
    1.029132e+10, 1.020515e+10, 1.011536e+10, 1.00221e+10, 9.925557e+09, 
    9.825887e+09, 9.723264e+09, 9.61786e+09, 9.509846e+09, 9.399396e+09, 
    9.286681e+09, 9.171869e+09, 9.055129e+09, 8.936627e+09, 8.816526e+09, 
    8.694987e+09, 8.572165e+09, 8.448214e+09, 8.323282e+09, 8.197513e+09, 
    8.071048e+09, 7.94402e+09, 7.816561e+09, 7.688794e+09, 7.56084e+09, 
    7.432814e+09, 7.304823e+09, 7.176973e+09, 7.049361e+09, 6.922081e+09, 
    6.795221e+09,
  6.76529e+09, 6.889429e+09, 7.013901e+09, 7.13862e+09, 7.263496e+09, 
    7.388432e+09, 7.513327e+09, 7.638074e+09, 7.762563e+09, 7.886679e+09, 
    8.010299e+09, 8.133301e+09, 8.255552e+09, 8.37692e+09, 8.497266e+09, 
    8.616447e+09, 8.734319e+09, 8.85073e+09, 8.96553e+09, 9.078562e+09, 
    9.18967e+09, 9.298694e+09, 9.405474e+09, 9.509846e+09, 9.61165e+09, 
    9.710721e+09, 9.806899e+09, 9.900023e+09, 9.989933e+09, 1.007647e+10, 
    1.015949e+10, 1.023883e+10, 1.031435e+10, 1.03859e+10, 1.045336e+10, 
    1.051658e+10, 1.057545e+10, 1.062985e+10, 1.067967e+10, 1.07248e+10, 
    1.076517e+10, 1.080067e+10, 1.083124e+10, 1.085682e+10, 1.087735e+10, 
    1.089278e+10, 1.090309e+10, 1.090825e+10, 1.090825e+10, 1.090309e+10, 
    1.089278e+10, 1.087735e+10, 1.085682e+10, 1.083124e+10, 1.080067e+10, 
    1.076517e+10, 1.07248e+10, 1.067967e+10, 1.062985e+10, 1.057545e+10, 
    1.051658e+10, 1.045336e+10, 1.03859e+10, 1.031435e+10, 1.023883e+10, 
    1.015949e+10, 1.007647e+10, 9.989933e+09, 9.900023e+09, 9.806899e+09, 
    9.710721e+09, 9.61165e+09, 9.509846e+09, 9.405474e+09, 9.298694e+09, 
    9.18967e+09, 9.078562e+09, 8.96553e+09, 8.85073e+09, 8.734319e+09, 
    8.616447e+09, 8.497266e+09, 8.37692e+09, 8.255552e+09, 8.133301e+09, 
    8.010299e+09, 7.886679e+09, 7.762563e+09, 7.638074e+09, 7.513327e+09, 
    7.388432e+09, 7.263496e+09, 7.13862e+09, 7.013901e+09, 6.889429e+09, 
    6.76529e+09,
  6.734221e+09, 6.855565e+09, 6.977157e+09, 7.098912e+09, 7.220742e+09, 
    7.342552e+09, 7.464245e+09, 7.585717e+09, 7.706863e+09, 7.827569e+09, 
    7.94772e+09, 8.067195e+09, 8.18587e+09, 8.303616e+09, 8.420301e+09, 
    8.53579e+09, 8.649944e+09, 8.762619e+09, 8.873673e+09, 8.982957e+09, 
    9.090322e+09, 9.195619e+09, 9.298694e+09, 9.399396e+09, 9.497571e+09, 
    9.593066e+09, 9.68573e+09, 9.775411e+09, 9.861961e+09, 9.945231e+09, 
    1.002508e+10, 1.010136e+10, 1.017395e+10, 1.02427e+10, 1.030749e+10, 
    1.03682e+10, 1.042471e+10, 1.047692e+10, 1.052472e+10, 1.056802e+10, 
    1.060673e+10, 1.064077e+10, 1.067009e+10, 1.06946e+10, 1.071428e+10, 
    1.072907e+10, 1.073895e+10, 1.07439e+10, 1.07439e+10, 1.073895e+10, 
    1.072907e+10, 1.071428e+10, 1.06946e+10, 1.067009e+10, 1.064077e+10, 
    1.060673e+10, 1.056802e+10, 1.052472e+10, 1.047692e+10, 1.042471e+10, 
    1.03682e+10, 1.030749e+10, 1.02427e+10, 1.017395e+10, 1.010136e+10, 
    1.002508e+10, 9.945231e+09, 9.861961e+09, 9.775411e+09, 9.68573e+09, 
    9.593066e+09, 9.497571e+09, 9.399396e+09, 9.298694e+09, 9.195619e+09, 
    9.090322e+09, 8.982957e+09, 8.873673e+09, 8.762619e+09, 8.649944e+09, 
    8.53579e+09, 8.420301e+09, 8.303616e+09, 8.18587e+09, 8.067195e+09, 
    7.94772e+09, 7.827569e+09, 7.706863e+09, 7.585717e+09, 7.464245e+09, 
    7.342552e+09, 7.220742e+09, 7.098912e+09, 6.977157e+09, 6.855565e+09, 
    6.734221e+09,
  6.702019e+09, 6.8205e+09, 6.939143e+09, 7.057866e+09, 7.176583e+09, 
    7.295202e+09, 7.41363e+09, 7.531766e+09, 7.649507e+09, 7.766745e+09, 
    7.883369e+09, 7.999264e+09, 8.11431e+09, 8.228386e+09, 8.341364e+09, 
    8.453116e+09, 8.563511e+09, 8.672412e+09, 8.779684e+09, 8.885187e+09, 
    8.988781e+09, 9.090322e+09, 9.18967e+09, 9.286681e+09, 9.381209e+09, 
    9.473112e+09, 9.562249e+09, 9.648477e+09, 9.731658e+09, 9.811654e+09, 
    9.88833e+09, 9.961556e+09, 1.00312e+10, 1.009715e+10, 1.015928e+10, 
    1.021748e+10, 1.027164e+10, 1.032166e+10, 1.036744e+10, 1.040891e+10, 
    1.044597e+10, 1.047856e+10, 1.050662e+10, 1.053008e+10, 1.054891e+10, 
    1.056306e+10, 1.057252e+10, 1.057725e+10, 1.057725e+10, 1.057252e+10, 
    1.056306e+10, 1.054891e+10, 1.053008e+10, 1.050662e+10, 1.047856e+10, 
    1.044597e+10, 1.040891e+10, 1.036744e+10, 1.032166e+10, 1.027164e+10, 
    1.021748e+10, 1.015928e+10, 1.009715e+10, 1.00312e+10, 9.961556e+09, 
    9.88833e+09, 9.811654e+09, 9.731658e+09, 9.648477e+09, 9.562249e+09, 
    9.473112e+09, 9.381209e+09, 9.286681e+09, 9.18967e+09, 9.090322e+09, 
    8.988781e+09, 8.885187e+09, 8.779684e+09, 8.672412e+09, 8.563511e+09, 
    8.453116e+09, 8.341364e+09, 8.228386e+09, 8.11431e+09, 7.999264e+09, 
    7.883369e+09, 7.766745e+09, 7.649507e+09, 7.531766e+09, 7.41363e+09, 
    7.295202e+09, 7.176583e+09, 7.057866e+09, 6.939143e+09, 6.8205e+09, 
    6.702019e+09,
  6.668692e+09, 6.784244e+09, 6.899874e+09, 7.015503e+09, 7.131045e+09, 
    7.246414e+09, 7.361518e+09, 7.47626e+09, 7.590542e+09, 7.704261e+09, 
    7.817309e+09, 7.929576e+09, 8.04095e+09, 8.151313e+09, 8.260545e+09, 
    8.368525e+09, 8.475127e+09, 8.580225e+09, 8.683688e+09, 8.785385e+09, 
    8.885187e+09, 8.982957e+09, 9.078562e+09, 9.171869e+09, 9.262742e+09, 
    9.351046e+09, 9.436652e+09, 9.519426e+09, 9.599237e+09, 9.67596e+09, 
    9.749469e+09, 9.819643e+09, 9.886363e+09, 9.949515e+09, 1.000899e+10, 
    1.006469e+10, 1.01165e+10, 1.016434e+10, 1.020812e+10, 1.024776e+10, 
    1.028319e+10, 1.031433e+10, 1.034114e+10, 1.036355e+10, 1.038154e+10, 
    1.039506e+10, 1.040409e+10, 1.040861e+10, 1.040861e+10, 1.040409e+10, 
    1.039506e+10, 1.038154e+10, 1.036355e+10, 1.034114e+10, 1.031433e+10, 
    1.028319e+10, 1.024776e+10, 1.020812e+10, 1.016434e+10, 1.01165e+10, 
    1.006469e+10, 1.000899e+10, 9.949515e+09, 9.886363e+09, 9.819643e+09, 
    9.749469e+09, 9.67596e+09, 9.599237e+09, 9.519426e+09, 9.436652e+09, 
    9.351046e+09, 9.262742e+09, 9.171869e+09, 9.078562e+09, 8.982957e+09, 
    8.885187e+09, 8.785385e+09, 8.683688e+09, 8.580225e+09, 8.475127e+09, 
    8.368525e+09, 8.260545e+09, 8.151313e+09, 8.04095e+09, 7.929576e+09, 
    7.817309e+09, 7.704261e+09, 7.590542e+09, 7.47626e+09, 7.361518e+09, 
    7.246414e+09, 7.131045e+09, 7.015503e+09, 6.899874e+09, 6.784244e+09, 
    6.668692e+09,
  6.634248e+09, 6.74681e+09, 6.859367e+09, 6.971842e+09, 7.084154e+09, 
    7.196217e+09, 7.307944e+09, 7.419243e+09, 7.530018e+09, 7.640172e+09, 
    7.749601e+09, 7.858201e+09, 7.965864e+09, 8.072481e+09, 8.177936e+09, 
    8.282116e+09, 8.384902e+09, 8.486173e+09, 8.585809e+09, 8.683688e+09, 
    8.779684e+09, 8.873673e+09, 8.96553e+09, 9.055129e+09, 9.142345e+09, 
    9.227054e+09, 9.309132e+09, 9.388457e+09, 9.464909e+09, 9.53837e+09, 
    9.608722e+09, 9.675857e+09, 9.739662e+09, 9.800034e+09, 9.856871e+09, 
    9.910078e+09, 9.959563e+09, 1.000524e+10, 1.004703e+10, 1.008486e+10, 
    1.011866e+10, 1.014837e+10, 1.017394e+10, 1.019532e+10, 1.021247e+10, 
    1.022536e+10, 1.023397e+10, 1.023827e+10, 1.023827e+10, 1.023397e+10, 
    1.022536e+10, 1.021247e+10, 1.019532e+10, 1.017394e+10, 1.014837e+10, 
    1.011866e+10, 1.008486e+10, 1.004703e+10, 1.000524e+10, 9.959563e+09, 
    9.910078e+09, 9.856871e+09, 9.800034e+09, 9.739662e+09, 9.675857e+09, 
    9.608722e+09, 9.53837e+09, 9.464909e+09, 9.388457e+09, 9.309132e+09, 
    9.227054e+09, 9.142345e+09, 9.055129e+09, 8.96553e+09, 8.873673e+09, 
    8.779684e+09, 8.683688e+09, 8.585809e+09, 8.486173e+09, 8.384902e+09, 
    8.282116e+09, 8.177936e+09, 8.072481e+09, 7.965864e+09, 7.858201e+09, 
    7.749601e+09, 7.640172e+09, 7.530018e+09, 7.419243e+09, 7.307944e+09, 
    7.196217e+09, 7.084154e+09, 6.971842e+09, 6.859367e+09, 6.74681e+09, 
    6.634248e+09,
  6.598693e+09, 6.708208e+09, 6.817636e+09, 6.926904e+09, 7.035934e+09, 
    7.144643e+09, 7.252946e+09, 7.360757e+09, 7.467984e+09, 7.574533e+09, 
    7.680307e+09, 7.785207e+09, 7.889131e+09, 7.991974e+09, 8.093629e+09, 
    8.193989e+09, 8.292941e+09, 8.390374e+09, 8.486173e+09, 8.580225e+09, 
    8.672412e+09, 8.762619e+09, 8.85073e+09, 8.936627e+09, 9.020195e+09, 
    9.101317e+09, 9.17988e+09, 9.255772e+09, 9.32888e+09, 9.399095e+09, 
    9.466312e+09, 9.530426e+09, 9.591338e+09, 9.64895e+09, 9.703171e+09, 
    9.753911e+09, 9.801088e+09, 9.844622e+09, 9.884442e+09, 9.920478e+09, 
    9.95267e+09, 9.980962e+09, 1.00053e+10, 1.002566e+10, 1.004198e+10, 
    1.005425e+10, 1.006244e+10, 1.006654e+10, 1.006654e+10, 1.006244e+10, 
    1.005425e+10, 1.004198e+10, 1.002566e+10, 1.00053e+10, 9.980962e+09, 
    9.95267e+09, 9.920478e+09, 9.884442e+09, 9.844622e+09, 9.801088e+09, 
    9.753911e+09, 9.703171e+09, 9.64895e+09, 9.591338e+09, 9.530426e+09, 
    9.466312e+09, 9.399095e+09, 9.32888e+09, 9.255772e+09, 9.17988e+09, 
    9.101317e+09, 9.020195e+09, 8.936627e+09, 8.85073e+09, 8.762619e+09, 
    8.672412e+09, 8.580225e+09, 8.486173e+09, 8.390374e+09, 8.292941e+09, 
    8.193989e+09, 8.093629e+09, 7.991974e+09, 7.889131e+09, 7.785207e+09, 
    7.680307e+09, 7.574533e+09, 7.467984e+09, 7.360757e+09, 7.252946e+09, 
    7.144643e+09, 7.035934e+09, 6.926904e+09, 6.817636e+09, 6.708208e+09, 
    6.598693e+09,
  6.562035e+09, 6.668449e+09, 6.774699e+09, 6.880711e+09, 6.986412e+09, 
    7.091722e+09, 7.196561e+09, 7.300845e+09, 7.404488e+09, 7.5074e+09, 
    7.60949e+09, 7.710664e+09, 7.810825e+09, 7.909876e+09, 8.007716e+09, 
    8.104243e+09, 8.199353e+09, 8.292941e+09, 8.384902e+09, 8.475127e+09, 
    8.563511e+09, 8.649944e+09, 8.734319e+09, 8.816526e+09, 8.896461e+09, 
    8.974015e+09, 9.049084e+09, 9.121564e+09, 9.191351e+09, 9.258346e+09, 
    9.322452e+09, 9.383574e+09, 9.441618e+09, 9.496498e+09, 9.548129e+09, 
    9.596429e+09, 9.641325e+09, 9.68274e+09, 9.720613e+09, 9.754878e+09, 
    9.785482e+09, 9.812372e+09, 9.835507e+09, 9.854844e+09, 9.870353e+09, 
    9.882009e+09, 9.88979e+09, 9.893683e+09, 9.893683e+09, 9.88979e+09, 
    9.882009e+09, 9.870353e+09, 9.854844e+09, 9.835507e+09, 9.812372e+09, 
    9.785482e+09, 9.754878e+09, 9.720613e+09, 9.68274e+09, 9.641325e+09, 
    9.596429e+09, 9.548129e+09, 9.496498e+09, 9.441618e+09, 9.383574e+09, 
    9.322452e+09, 9.258346e+09, 9.191351e+09, 9.121564e+09, 9.049084e+09, 
    8.974015e+09, 8.896461e+09, 8.816526e+09, 8.734319e+09, 8.649944e+09, 
    8.563511e+09, 8.475127e+09, 8.384902e+09, 8.292941e+09, 8.199353e+09, 
    8.104243e+09, 8.007716e+09, 7.909876e+09, 7.810825e+09, 7.710664e+09, 
    7.60949e+09, 7.5074e+09, 7.404488e+09, 7.300845e+09, 7.196561e+09, 
    7.091722e+09, 6.986412e+09, 6.880711e+09, 6.774699e+09, 6.668449e+09, 
    6.562035e+09,
  6.524282e+09, 6.627547e+09, 6.730571e+09, 6.833284e+09, 6.935614e+09, 
    7.037487e+09, 7.138825e+09, 7.23955e+09, 7.339579e+09, 7.438829e+09, 
    7.537212e+09, 7.634641e+09, 7.731025e+09, 7.826271e+09, 7.920287e+09, 
    8.012976e+09, 8.104243e+09, 8.193989e+09, 8.282116e+09, 8.368525e+09, 
    8.453116e+09, 8.53579e+09, 8.616447e+09, 8.694987e+09, 8.771312e+09, 
    8.845323e+09, 8.916924e+09, 8.986021e+09, 9.052518e+09, 9.116325e+09, 
    9.177352e+09, 9.235513e+09, 9.290724e+09, 9.342905e+09, 9.391978e+09, 
    9.437871e+09, 9.480515e+09, 9.519842e+09, 9.555794e+09, 9.588315e+09, 
    9.617354e+09, 9.642865e+09, 9.664807e+09, 9.683147e+09, 9.697854e+09, 
    9.708905e+09, 9.716282e+09, 9.719975e+09, 9.719975e+09, 9.716282e+09, 
    9.708905e+09, 9.697854e+09, 9.683147e+09, 9.664807e+09, 9.642865e+09, 
    9.617354e+09, 9.588315e+09, 9.555794e+09, 9.519842e+09, 9.480515e+09, 
    9.437871e+09, 9.391978e+09, 9.342905e+09, 9.290724e+09, 9.235513e+09, 
    9.177352e+09, 9.116325e+09, 9.052518e+09, 8.986021e+09, 8.916924e+09, 
    8.845323e+09, 8.771312e+09, 8.694987e+09, 8.616447e+09, 8.53579e+09, 
    8.453116e+09, 8.368525e+09, 8.282116e+09, 8.193989e+09, 8.104243e+09, 
    8.012976e+09, 7.920287e+09, 7.826271e+09, 7.731025e+09, 7.634641e+09, 
    7.537212e+09, 7.438829e+09, 7.339579e+09, 7.23955e+09, 7.138825e+09, 
    7.037487e+09, 6.935614e+09, 6.833284e+09, 6.730571e+09, 6.627547e+09, 
    6.524282e+09,
  6.485442e+09, 6.585513e+09, 6.685269e+09, 6.784643e+09, 6.883567e+09, 
    6.981969e+09, 7.079777e+09, 7.176916e+09, 7.273309e+09, 7.368877e+09, 
    7.463537e+09, 7.557208e+09, 7.649805e+09, 7.741242e+09, 7.831433e+09, 
    7.920287e+09, 8.007716e+09, 8.093629e+09, 8.177936e+09, 8.260545e+09, 
    8.341364e+09, 8.420301e+09, 8.497266e+09, 8.572165e+09, 8.64491e+09, 
    8.715411e+09, 8.78358e+09, 8.849328e+09, 8.912572e+09, 8.973229e+09, 
    9.031216e+09, 9.086456e+09, 9.138871e+09, 9.188391e+09, 9.234944e+09, 
    9.278465e+09, 9.318892e+09, 9.356163e+09, 9.390226e+09, 9.421031e+09, 
    9.448532e+09, 9.472687e+09, 9.49346e+09, 9.510819e+09, 9.524738e+09, 
    9.535196e+09, 9.542177e+09, 9.54567e+09, 9.54567e+09, 9.542177e+09, 
    9.535196e+09, 9.524738e+09, 9.510819e+09, 9.49346e+09, 9.472687e+09, 
    9.448532e+09, 9.421031e+09, 9.390226e+09, 9.356163e+09, 9.318892e+09, 
    9.278465e+09, 9.234944e+09, 9.188391e+09, 9.138871e+09, 9.086456e+09, 
    9.031216e+09, 8.973229e+09, 8.912572e+09, 8.849328e+09, 8.78358e+09, 
    8.715411e+09, 8.64491e+09, 8.572165e+09, 8.497266e+09, 8.420301e+09, 
    8.341364e+09, 8.260545e+09, 8.177936e+09, 8.093629e+09, 8.007716e+09, 
    7.920287e+09, 7.831433e+09, 7.741242e+09, 7.649805e+09, 7.557208e+09, 
    7.463537e+09, 7.368877e+09, 7.273309e+09, 7.176916e+09, 7.079777e+09, 
    6.981969e+09, 6.883567e+09, 6.784643e+09, 6.685269e+09, 6.585513e+09, 
    6.485442e+09,
  6.445522e+09, 6.54236e+09, 6.638811e+09, 6.734811e+09, 6.830297e+09, 
    6.925201e+09, 7.019455e+09, 7.112987e+09, 7.205726e+09, 7.297597e+09, 
    7.388526e+09, 7.478433e+09, 7.567242e+09, 7.654872e+09, 7.741242e+09, 
    7.826271e+09, 7.909876e+09, 7.991974e+09, 8.072481e+09, 8.151313e+09, 
    8.228386e+09, 8.303616e+09, 8.37692e+09, 8.448214e+09, 8.517416e+09, 
    8.584445e+09, 8.649221e+09, 8.711665e+09, 8.771699e+09, 8.829247e+09, 
    8.884238e+09, 8.936601e+09, 8.986266e+09, 9.033167e+09, 9.077242e+09, 
    9.118431e+09, 9.156679e+09, 9.191932e+09, 9.224142e+09, 9.253263e+09, 
    9.279254e+09, 9.302078e+09, 9.321703e+09, 9.338102e+09, 9.351248e+09, 
    9.361125e+09, 9.367718e+09, 9.371016e+09, 9.371016e+09, 9.367718e+09, 
    9.361125e+09, 9.351248e+09, 9.338102e+09, 9.321703e+09, 9.302078e+09, 
    9.279254e+09, 9.253263e+09, 9.224142e+09, 9.191932e+09, 9.156679e+09, 
    9.118431e+09, 9.077242e+09, 9.033167e+09, 8.986266e+09, 8.936601e+09, 
    8.884238e+09, 8.829247e+09, 8.771699e+09, 8.711665e+09, 8.649221e+09, 
    8.584445e+09, 8.517416e+09, 8.448214e+09, 8.37692e+09, 8.303616e+09, 
    8.228386e+09, 8.151313e+09, 8.072481e+09, 7.991974e+09, 7.909876e+09, 
    7.826271e+09, 7.741242e+09, 7.654872e+09, 7.567242e+09, 7.478433e+09, 
    7.388526e+09, 7.297597e+09, 7.205726e+09, 7.112987e+09, 7.019455e+09, 
    6.925201e+09, 6.830297e+09, 6.734811e+09, 6.638811e+09, 6.54236e+09, 
    6.445522e+09,
  6.404531e+09, 6.4981e+09, 6.591213e+09, 6.683811e+09, 6.775833e+09, 
    6.867216e+09, 6.957896e+09, 7.047806e+09, 7.136881e+09, 7.225049e+09, 
    7.312241e+09, 7.398386e+09, 7.483411e+09, 7.567242e+09, 7.649805e+09, 
    7.731025e+09, 7.810825e+09, 7.889131e+09, 7.965864e+09, 8.04095e+09, 
    8.11431e+09, 8.18587e+09, 8.255552e+09, 8.323282e+09, 8.388985e+09, 
    8.452588e+09, 8.514017e+09, 8.573202e+09, 8.630074e+09, 8.684566e+09, 
    8.736609e+09, 8.786142e+09, 8.833104e+09, 8.877434e+09, 8.919077e+09, 
    8.95798e+09, 8.994092e+09, 9.027367e+09, 9.05776e+09, 9.085231e+09, 
    9.109745e+09, 9.131267e+09, 9.14977e+09, 9.165227e+09, 9.177618e+09, 
    9.186927e+09, 9.193139e+09, 9.196247e+09, 9.196247e+09, 9.193139e+09, 
    9.186927e+09, 9.177618e+09, 9.165227e+09, 9.14977e+09, 9.131267e+09, 
    9.109745e+09, 9.085231e+09, 9.05776e+09, 9.027367e+09, 8.994092e+09, 
    8.95798e+09, 8.919077e+09, 8.877434e+09, 8.833104e+09, 8.786142e+09, 
    8.736609e+09, 8.684566e+09, 8.630074e+09, 8.573202e+09, 8.514017e+09, 
    8.452588e+09, 8.388985e+09, 8.323282e+09, 8.255552e+09, 8.18587e+09, 
    8.11431e+09, 8.04095e+09, 7.965864e+09, 7.889131e+09, 7.810825e+09, 
    7.731025e+09, 7.649805e+09, 7.567242e+09, 7.483411e+09, 7.398386e+09, 
    7.312241e+09, 7.225049e+09, 7.136881e+09, 7.047806e+09, 6.957896e+09, 
    6.867216e+09, 6.775833e+09, 6.683811e+09, 6.591213e+09, 6.4981e+09, 
    6.404531e+09,
  6.362479e+09, 6.452746e+09, 6.542493e+09, 6.631664e+09, 6.720201e+09, 
    6.808046e+09, 6.895139e+09, 6.981418e+09, 7.066822e+09, 7.151286e+09, 
    7.234745e+09, 7.317134e+09, 7.398386e+09, 7.478433e+09, 7.557208e+09, 
    7.634641e+09, 7.710664e+09, 7.785207e+09, 7.858201e+09, 7.929576e+09, 
    7.999264e+09, 8.067195e+09, 8.133301e+09, 8.197513e+09, 8.259766e+09, 
    8.319992e+09, 8.378128e+09, 8.434108e+09, 8.487873e+09, 8.539359e+09, 
    8.58851e+09, 8.635267e+09, 8.679578e+09, 8.721389e+09, 8.760649e+09, 
    8.797313e+09, 8.831335e+09, 8.862674e+09, 8.891291e+09, 8.917151e+09, 
    8.940219e+09, 8.96047e+09, 8.977876e+09, 8.992415e+09, 9.004068e+09, 
    9.012821e+09, 9.018663e+09, 9.021585e+09, 9.021585e+09, 9.018663e+09, 
    9.012821e+09, 9.004068e+09, 8.992415e+09, 8.977876e+09, 8.96047e+09, 
    8.940219e+09, 8.917151e+09, 8.891291e+09, 8.862674e+09, 8.831335e+09, 
    8.797313e+09, 8.760649e+09, 8.721389e+09, 8.679578e+09, 8.635267e+09, 
    8.58851e+09, 8.539359e+09, 8.487873e+09, 8.434108e+09, 8.378128e+09, 
    8.319992e+09, 8.259766e+09, 8.197513e+09, 8.133301e+09, 8.067195e+09, 
    7.999264e+09, 7.929576e+09, 7.858201e+09, 7.785207e+09, 7.710664e+09, 
    7.634641e+09, 7.557208e+09, 7.478433e+09, 7.398386e+09, 7.317134e+09, 
    7.234745e+09, 7.151286e+09, 7.066822e+09, 6.981418e+09, 6.895139e+09, 
    6.808046e+09, 6.720201e+09, 6.631664e+09, 6.542493e+09, 6.452746e+09, 
    6.362479e+09,
  6.319373e+09, 6.406312e+09, 6.492669e+09, 6.578392e+09, 6.663429e+09, 
    6.747724e+09, 6.831222e+09, 6.913867e+09, 6.9956e+09, 7.076365e+09, 
    7.1561e+09, 7.234745e+09, 7.312241e+09, 7.388526e+09, 7.463537e+09, 
    7.537212e+09, 7.60949e+09, 7.680307e+09, 7.749601e+09, 7.817309e+09, 
    7.883369e+09, 7.94772e+09, 8.010299e+09, 8.071048e+09, 8.129904e+09, 
    8.186811e+09, 8.241709e+09, 8.294543e+09, 8.345257e+09, 8.393798e+09, 
    8.440113e+09, 8.484152e+09, 8.525868e+09, 8.565214e+09, 8.602145e+09, 
    8.636621e+09, 8.668601e+09, 8.698051e+09, 8.724934e+09, 8.749221e+09, 
    8.770882e+09, 8.789891e+09, 8.806228e+09, 8.819871e+09, 8.830806e+09, 
    8.839017e+09, 8.844498e+09, 8.84724e+09, 8.84724e+09, 8.844498e+09, 
    8.839017e+09, 8.830806e+09, 8.819871e+09, 8.806228e+09, 8.789891e+09, 
    8.770882e+09, 8.749221e+09, 8.724934e+09, 8.698051e+09, 8.668601e+09, 
    8.636621e+09, 8.602145e+09, 8.565214e+09, 8.525868e+09, 8.484152e+09, 
    8.440113e+09, 8.393798e+09, 8.345257e+09, 8.294543e+09, 8.241709e+09, 
    8.186811e+09, 8.129904e+09, 8.071048e+09, 8.010299e+09, 7.94772e+09, 
    7.883369e+09, 7.817309e+09, 7.749601e+09, 7.680307e+09, 7.60949e+09, 
    7.537212e+09, 7.463537e+09, 7.388526e+09, 7.312241e+09, 7.234745e+09, 
    7.1561e+09, 7.076365e+09, 6.9956e+09, 6.913867e+09, 6.831222e+09, 
    6.747724e+09, 6.663429e+09, 6.578392e+09, 6.492669e+09, 6.406312e+09, 
    6.319373e+09,
  6.275223e+09, 6.35881e+09, 6.441759e+09, 6.52402e+09, 6.605544e+09, 
    6.686283e+09, 6.766183e+09, 6.845195e+09, 6.923265e+09, 7.000339e+09, 
    7.076365e+09, 7.151286e+09, 7.225049e+09, 7.297597e+09, 7.368877e+09, 
    7.438829e+09, 7.5074e+09, 7.574533e+09, 7.640172e+09, 7.704261e+09, 
    7.766745e+09, 7.827569e+09, 7.886679e+09, 7.94402e+09, 7.99954e+09, 
    8.053188e+09, 8.10491e+09, 8.15466e+09, 8.202386e+09, 8.248043e+09, 
    8.291585e+09, 8.332967e+09, 8.372148e+09, 8.409087e+09, 8.443745e+09, 
    8.476086e+09, 8.506077e+09, 8.533684e+09, 8.558878e+09, 8.581632e+09, 
    8.601922e+09, 8.619724e+09, 8.63502e+09, 8.647793e+09, 8.658028e+09, 
    8.665715e+09, 8.670843e+09, 8.673409e+09, 8.673409e+09, 8.670843e+09, 
    8.665715e+09, 8.658028e+09, 8.647793e+09, 8.63502e+09, 8.619724e+09, 
    8.601922e+09, 8.581632e+09, 8.558878e+09, 8.533684e+09, 8.506077e+09, 
    8.476086e+09, 8.443745e+09, 8.409087e+09, 8.372148e+09, 8.332967e+09, 
    8.291585e+09, 8.248043e+09, 8.202386e+09, 8.15466e+09, 8.10491e+09, 
    8.053188e+09, 7.99954e+09, 7.94402e+09, 7.886679e+09, 7.827569e+09, 
    7.766745e+09, 7.704261e+09, 7.640172e+09, 7.574533e+09, 7.5074e+09, 
    7.438829e+09, 7.368877e+09, 7.297597e+09, 7.225049e+09, 7.151286e+09, 
    7.076365e+09, 7.000339e+09, 6.923265e+09, 6.845195e+09, 6.766183e+09, 
    6.686283e+09, 6.605544e+09, 6.52402e+09, 6.441759e+09, 6.35881e+09, 
    6.275223e+09,
  6.230037e+09, 6.310255e+09, 6.38978e+09, 6.468569e+09, 6.546576e+09, 
    6.623755e+09, 6.700061e+09, 6.775447e+09, 6.849864e+09, 6.923265e+09, 
    6.9956e+09, 7.066822e+09, 7.136881e+09, 7.205726e+09, 7.273309e+09, 
    7.339579e+09, 7.404488e+09, 7.467984e+09, 7.530018e+09, 7.590542e+09, 
    7.649507e+09, 7.706863e+09, 7.762563e+09, 7.816561e+09, 7.868808e+09, 
    7.919261e+09, 7.967875e+09, 8.014606e+09, 8.059411e+09, 8.10225e+09, 
    8.143084e+09, 8.181873e+09, 8.218582e+09, 8.253174e+09, 8.285618e+09, 
    8.31588e+09, 8.343933e+09, 8.369748e+09, 8.3933e+09, 8.414565e+09, 
    8.433522e+09, 8.450151e+09, 8.464436e+09, 8.476363e+09, 8.485919e+09, 
    8.493095e+09, 8.497883e+09, 8.500278e+09, 8.500278e+09, 8.497883e+09, 
    8.493095e+09, 8.485919e+09, 8.476363e+09, 8.464436e+09, 8.450151e+09, 
    8.433522e+09, 8.414565e+09, 8.3933e+09, 8.369748e+09, 8.343933e+09, 
    8.31588e+09, 8.285618e+09, 8.253174e+09, 8.218582e+09, 8.181873e+09, 
    8.143084e+09, 8.10225e+09, 8.059411e+09, 8.014606e+09, 7.967875e+09, 
    7.919261e+09, 7.868808e+09, 7.816561e+09, 7.762563e+09, 7.706863e+09, 
    7.649507e+09, 7.590542e+09, 7.530018e+09, 7.467984e+09, 7.404488e+09, 
    7.339579e+09, 7.273309e+09, 7.205726e+09, 7.136881e+09, 7.066822e+09, 
    6.9956e+09, 6.923265e+09, 6.849864e+09, 6.775447e+09, 6.700061e+09, 
    6.623755e+09, 6.546576e+09, 6.468569e+09, 6.38978e+09, 6.310255e+09, 
    6.230037e+09,
  6.183825e+09, 6.260659e+09, 6.336752e+09, 6.412062e+09, 6.486551e+09, 
    6.560175e+09, 6.632894e+09, 6.704666e+09, 6.775447e+09, 6.845195e+09, 
    6.913867e+09, 6.981418e+09, 7.047806e+09, 7.112987e+09, 7.176916e+09, 
    7.23955e+09, 7.300845e+09, 7.360757e+09, 7.419243e+09, 7.47626e+09, 
    7.531766e+09, 7.585717e+09, 7.638074e+09, 7.688794e+09, 7.737838e+09, 
    7.785166e+09, 7.830739e+09, 7.874522e+09, 7.916475e+09, 7.956566e+09, 
    7.994759e+09, 8.031022e+09, 8.065324e+09, 8.097633e+09, 8.127923e+09, 
    8.156166e+09, 8.182336e+09, 8.20641e+09, 8.228367e+09, 8.248187e+09, 
    8.26585e+09, 8.281342e+09, 8.294647e+09, 8.305754e+09, 8.314652e+09, 
    8.321333e+09, 8.32579e+09, 8.32802e+09, 8.32802e+09, 8.32579e+09, 
    8.321333e+09, 8.314652e+09, 8.305754e+09, 8.294647e+09, 8.281342e+09, 
    8.26585e+09, 8.248187e+09, 8.228367e+09, 8.20641e+09, 8.182336e+09, 
    8.156166e+09, 8.127923e+09, 8.097633e+09, 8.065324e+09, 8.031022e+09, 
    7.994759e+09, 7.956566e+09, 7.916475e+09, 7.874522e+09, 7.830739e+09, 
    7.785166e+09, 7.737838e+09, 7.688794e+09, 7.638074e+09, 7.585717e+09, 
    7.531766e+09, 7.47626e+09, 7.419243e+09, 7.360757e+09, 7.300845e+09, 
    7.23955e+09, 7.176916e+09, 7.112987e+09, 7.047806e+09, 6.981418e+09, 
    6.913867e+09, 6.845195e+09, 6.775447e+09, 6.704666e+09, 6.632894e+09, 
    6.560175e+09, 6.486551e+09, 6.412062e+09, 6.336752e+09, 6.260659e+09, 
    6.183825e+09,
  6.136596e+09, 6.210038e+09, 6.282692e+09, 6.354524e+09, 6.425497e+09, 
    6.495574e+09, 6.564719e+09, 6.632894e+09, 6.700061e+09, 6.766183e+09, 
    6.831222e+09, 6.895139e+09, 6.957896e+09, 7.019455e+09, 7.079777e+09, 
    7.138825e+09, 7.196561e+09, 7.252946e+09, 7.307944e+09, 7.361518e+09, 
    7.41363e+09, 7.464245e+09, 7.513327e+09, 7.56084e+09, 7.606751e+09, 
    7.651027e+09, 7.693634e+09, 7.734541e+09, 7.773715e+09, 7.811129e+09, 
    7.846753e+09, 7.880559e+09, 7.912521e+09, 7.942612e+09, 7.970811e+09, 
    7.997093e+09, 8.021437e+09, 8.043825e+09, 8.064236e+09, 8.082655e+09, 
    8.099066e+09, 8.113456e+09, 8.125813e+09, 8.136126e+09, 8.144387e+09, 
    8.150589e+09, 8.154726e+09, 8.156796e+09, 8.156796e+09, 8.154726e+09, 
    8.150589e+09, 8.144387e+09, 8.136126e+09, 8.125813e+09, 8.113456e+09, 
    8.099066e+09, 8.082655e+09, 8.064236e+09, 8.043825e+09, 8.021437e+09, 
    7.997093e+09, 7.970811e+09, 7.942612e+09, 7.912521e+09, 7.880559e+09, 
    7.846753e+09, 7.811129e+09, 7.773715e+09, 7.734541e+09, 7.693634e+09, 
    7.651027e+09, 7.606751e+09, 7.56084e+09, 7.513327e+09, 7.464245e+09, 
    7.41363e+09, 7.361518e+09, 7.307944e+09, 7.252946e+09, 7.196561e+09, 
    7.138825e+09, 7.079777e+09, 7.019455e+09, 6.957896e+09, 6.895139e+09, 
    6.831222e+09, 6.766183e+09, 6.700061e+09, 6.632894e+09, 6.564719e+09, 
    6.495574e+09, 6.425497e+09, 6.354524e+09, 6.282692e+09, 6.210038e+09, 
    6.136596e+09,
  6.088361e+09, 6.158404e+09, 6.227619e+09, 6.295976e+09, 6.363442e+09, 
    6.429985e+09, 6.495574e+09, 6.560175e+09, 6.623755e+09, 6.686283e+09, 
    6.747724e+09, 6.808046e+09, 6.867216e+09, 6.925201e+09, 6.981969e+09, 
    7.037487e+09, 7.091722e+09, 7.144643e+09, 7.196217e+09, 7.246414e+09, 
    7.295202e+09, 7.342552e+09, 7.388432e+09, 7.432814e+09, 7.475667e+09, 
    7.516966e+09, 7.556683e+09, 7.594789e+09, 7.631261e+09, 7.666072e+09, 
    7.699199e+09, 7.73062e+09, 7.760311e+09, 7.788252e+09, 7.814423e+09, 
    7.838806e+09, 7.861382e+09, 7.882135e+09, 7.901051e+09, 7.918115e+09, 
    7.933316e+09, 7.946641e+09, 7.958081e+09, 7.967627e+09, 7.975273e+09, 
    7.981012e+09, 7.984841e+09, 7.986756e+09, 7.986756e+09, 7.984841e+09, 
    7.981012e+09, 7.975273e+09, 7.967627e+09, 7.958081e+09, 7.946641e+09, 
    7.933316e+09, 7.918115e+09, 7.901051e+09, 7.882135e+09, 7.861382e+09, 
    7.838806e+09, 7.814423e+09, 7.788252e+09, 7.760311e+09, 7.73062e+09, 
    7.699199e+09, 7.666072e+09, 7.631261e+09, 7.594789e+09, 7.556683e+09, 
    7.516966e+09, 7.475667e+09, 7.432814e+09, 7.388432e+09, 7.342552e+09, 
    7.295202e+09, 7.246414e+09, 7.196217e+09, 7.144643e+09, 7.091722e+09, 
    7.037487e+09, 6.981969e+09, 6.925201e+09, 6.867216e+09, 6.808046e+09, 
    6.747724e+09, 6.686283e+09, 6.623755e+09, 6.560175e+09, 6.495574e+09, 
    6.429985e+09, 6.363442e+09, 6.295976e+09, 6.227619e+09, 6.158404e+09, 
    6.088361e+09,
  6.039129e+09, 6.105772e+09, 6.171552e+09, 6.236442e+09, 6.300414e+09, 
    6.363442e+09, 6.425497e+09, 6.486551e+09, 6.546576e+09, 6.605544e+09, 
    6.663429e+09, 6.720201e+09, 6.775833e+09, 6.830297e+09, 6.883567e+09, 
    6.935614e+09, 6.986412e+09, 7.035934e+09, 7.084154e+09, 7.131045e+09, 
    7.176583e+09, 7.220742e+09, 7.263496e+09, 7.304823e+09, 7.344698e+09, 
    7.383099e+09, 7.420003e+09, 7.455388e+09, 7.489233e+09, 7.521518e+09, 
    7.552224e+09, 7.581331e+09, 7.608822e+09, 7.634681e+09, 7.65889e+09, 
    7.681435e+09, 7.702302e+09, 7.721477e+09, 7.738948e+09, 7.754704e+09, 
    7.768736e+09, 7.781033e+09, 7.791588e+09, 7.800395e+09, 7.807448e+09, 
    7.812741e+09, 7.816271e+09, 7.818037e+09, 7.818037e+09, 7.816271e+09, 
    7.812741e+09, 7.807448e+09, 7.800395e+09, 7.791588e+09, 7.781033e+09, 
    7.768736e+09, 7.754704e+09, 7.738948e+09, 7.721477e+09, 7.702302e+09, 
    7.681435e+09, 7.65889e+09, 7.634681e+09, 7.608822e+09, 7.581331e+09, 
    7.552224e+09, 7.521518e+09, 7.489233e+09, 7.455388e+09, 7.420003e+09, 
    7.383099e+09, 7.344698e+09, 7.304823e+09, 7.263496e+09, 7.220742e+09, 
    7.176583e+09, 7.131045e+09, 7.084154e+09, 7.035934e+09, 6.986412e+09, 
    6.935614e+09, 6.883567e+09, 6.830297e+09, 6.775833e+09, 6.720201e+09, 
    6.663429e+09, 6.605544e+09, 6.546576e+09, 6.486551e+09, 6.425497e+09, 
    6.363442e+09, 6.300414e+09, 6.236442e+09, 6.171552e+09, 6.105772e+09, 
    6.039129e+09,
  5.988909e+09, 6.052155e+09, 6.114508e+09, 6.175945e+09, 6.236442e+09, 
    6.295976e+09, 6.354524e+09, 6.412062e+09, 6.468569e+09, 6.52402e+09, 
    6.578392e+09, 6.631664e+09, 6.683811e+09, 6.734811e+09, 6.784643e+09, 
    6.833284e+09, 6.880711e+09, 6.926904e+09, 6.971842e+09, 7.015503e+09, 
    7.057866e+09, 7.098912e+09, 7.13862e+09, 7.176973e+09, 7.21395e+09, 
    7.249533e+09, 7.283705e+09, 7.316448e+09, 7.347746e+09, 7.377583e+09, 
    7.405943e+09, 7.432813e+09, 7.458176e+09, 7.482021e+09, 7.504335e+09, 
    7.525106e+09, 7.544322e+09, 7.561974e+09, 7.578052e+09, 7.592547e+09, 
    7.605452e+09, 7.616759e+09, 7.626462e+09, 7.634556e+09, 7.641037e+09, 
    7.645901e+09, 7.649145e+09, 7.650767e+09, 7.650767e+09, 7.649145e+09, 
    7.645901e+09, 7.641037e+09, 7.634556e+09, 7.626462e+09, 7.616759e+09, 
    7.605452e+09, 7.592547e+09, 7.578052e+09, 7.561974e+09, 7.544322e+09, 
    7.525106e+09, 7.504335e+09, 7.482021e+09, 7.458176e+09, 7.432813e+09, 
    7.405943e+09, 7.377583e+09, 7.347746e+09, 7.316448e+09, 7.283705e+09, 
    7.249533e+09, 7.21395e+09, 7.176973e+09, 7.13862e+09, 7.098912e+09, 
    7.057866e+09, 7.015503e+09, 6.971842e+09, 6.926904e+09, 6.880711e+09, 
    6.833284e+09, 6.784643e+09, 6.734811e+09, 6.683811e+09, 6.631664e+09, 
    6.578392e+09, 6.52402e+09, 6.468569e+09, 6.412062e+09, 6.354524e+09, 
    6.295976e+09, 6.236442e+09, 6.175945e+09, 6.114508e+09, 6.052155e+09, 
    5.988909e+09,
  5.937712e+09, 5.99757e+09, 6.056508e+09, 6.114508e+09, 6.171552e+09, 
    6.227619e+09, 6.282692e+09, 6.336752e+09, 6.38978e+09, 6.441759e+09, 
    6.492669e+09, 6.542493e+09, 6.591213e+09, 6.638811e+09, 6.685269e+09, 
    6.730571e+09, 6.774699e+09, 6.817636e+09, 6.859367e+09, 6.899874e+09, 
    6.939143e+09, 6.977157e+09, 7.013901e+09, 7.049361e+09, 7.083523e+09, 
    7.116371e+09, 7.147894e+09, 7.178077e+09, 7.206909e+09, 7.234377e+09, 
    7.260469e+09, 7.285175e+09, 7.308484e+09, 7.330385e+09, 7.350871e+09, 
    7.36993e+09, 7.387556e+09, 7.403741e+09, 7.418477e+09, 7.431758e+09, 
    7.443579e+09, 7.453934e+09, 7.462817e+09, 7.470226e+09, 7.476158e+09, 
    7.480609e+09, 7.483577e+09, 7.485062e+09, 7.485062e+09, 7.483577e+09, 
    7.480609e+09, 7.476158e+09, 7.470226e+09, 7.462817e+09, 7.453934e+09, 
    7.443579e+09, 7.431758e+09, 7.418477e+09, 7.403741e+09, 7.387556e+09, 
    7.36993e+09, 7.350871e+09, 7.330385e+09, 7.308484e+09, 7.285175e+09, 
    7.260469e+09, 7.234377e+09, 7.206909e+09, 7.178077e+09, 7.147894e+09, 
    7.116371e+09, 7.083523e+09, 7.049361e+09, 7.013901e+09, 6.977157e+09, 
    6.939143e+09, 6.899874e+09, 6.859367e+09, 6.817636e+09, 6.774699e+09, 
    6.730571e+09, 6.685269e+09, 6.638811e+09, 6.591213e+09, 6.542493e+09, 
    6.492669e+09, 6.441759e+09, 6.38978e+09, 6.336752e+09, 6.282692e+09, 
    6.227619e+09, 6.171552e+09, 6.114508e+09, 6.056508e+09, 5.99757e+09, 
    5.937712e+09,
  5.885548e+09, 5.942029e+09, 5.99757e+09, 6.052155e+09, 6.105772e+09, 
    6.158404e+09, 6.210038e+09, 6.260659e+09, 6.310255e+09, 6.35881e+09, 
    6.406312e+09, 6.452746e+09, 6.4981e+09, 6.54236e+09, 6.585513e+09, 
    6.627547e+09, 6.668449e+09, 6.708208e+09, 6.74681e+09, 6.784244e+09, 
    6.8205e+09, 6.855565e+09, 6.889429e+09, 6.922081e+09, 6.953512e+09, 
    6.98371e+09, 7.012667e+09, 7.040374e+09, 7.066821e+09, 7.092e+09, 
    7.115902e+09, 7.138521e+09, 7.159848e+09, 7.179877e+09, 7.198601e+09, 
    7.216014e+09, 7.23211e+09, 7.246883e+09, 7.260329e+09, 7.272444e+09, 
    7.283223e+09, 7.292662e+09, 7.30076e+09, 7.307511e+09, 7.312915e+09, 
    7.316969e+09, 7.319673e+09, 7.321026e+09, 7.321026e+09, 7.319673e+09, 
    7.316969e+09, 7.312915e+09, 7.307511e+09, 7.30076e+09, 7.292662e+09, 
    7.283223e+09, 7.272444e+09, 7.260329e+09, 7.246883e+09, 7.23211e+09, 
    7.216014e+09, 7.198601e+09, 7.179877e+09, 7.159848e+09, 7.138521e+09, 
    7.115902e+09, 7.092e+09, 7.066821e+09, 7.040374e+09, 7.012667e+09, 
    6.98371e+09, 6.953512e+09, 6.922081e+09, 6.889429e+09, 6.855565e+09, 
    6.8205e+09, 6.784244e+09, 6.74681e+09, 6.708208e+09, 6.668449e+09, 
    6.627547e+09, 6.585513e+09, 6.54236e+09, 6.4981e+09, 6.452746e+09, 
    6.406312e+09, 6.35881e+09, 6.310255e+09, 6.260659e+09, 6.210038e+09, 
    6.158404e+09, 6.105772e+09, 6.052155e+09, 5.99757e+09, 5.942029e+09, 
    5.885548e+09,
  5.832426e+09, 5.885548e+09, 5.937712e+09, 5.988909e+09, 6.039129e+09, 
    6.088361e+09, 6.136596e+09, 6.183825e+09, 6.230037e+09, 6.275223e+09, 
    6.319373e+09, 6.362479e+09, 6.404531e+09, 6.445522e+09, 6.485442e+09, 
    6.524282e+09, 6.562035e+09, 6.598693e+09, 6.634248e+09, 6.668692e+09, 
    6.702019e+09, 6.734221e+09, 6.76529e+09, 6.795221e+09, 6.824007e+09, 
    6.851641e+09, 6.878117e+09, 6.903431e+09, 6.927576e+09, 6.950547e+09, 
    6.972339e+09, 6.992947e+09, 7.012366e+09, 7.030593e+09, 7.047623e+09, 
    7.063453e+09, 7.078078e+09, 7.091497e+09, 7.103705e+09, 7.1147e+09, 
    7.124479e+09, 7.133041e+09, 7.140384e+09, 7.146505e+09, 7.151404e+09, 
    7.155078e+09, 7.157529e+09, 7.158754e+09, 7.158754e+09, 7.157529e+09, 
    7.155078e+09, 7.151404e+09, 7.146505e+09, 7.140384e+09, 7.133041e+09, 
    7.124479e+09, 7.1147e+09, 7.103705e+09, 7.091497e+09, 7.078078e+09, 
    7.063453e+09, 7.047623e+09, 7.030593e+09, 7.012366e+09, 6.992947e+09, 
    6.972339e+09, 6.950547e+09, 6.927576e+09, 6.903431e+09, 6.878117e+09, 
    6.851641e+09, 6.824007e+09, 6.795221e+09, 6.76529e+09, 6.734221e+09, 
    6.702019e+09, 6.668692e+09, 6.634248e+09, 6.598693e+09, 6.562035e+09, 
    6.524282e+09, 6.485442e+09, 6.445522e+09, 6.404531e+09, 6.362479e+09, 
    6.319373e+09, 6.275223e+09, 6.230037e+09, 6.183825e+09, 6.136596e+09, 
    6.088361e+09, 6.039129e+09, 5.988909e+09, 5.937712e+09, 5.885548e+09, 
    5.832426e+09 ;

 bk = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.01253, 0.04887, 0.10724, 0.18455, 0.27461, 0.36914, 
    0.46103, 0.54623, 0.62305, 0.69099, 0.75016, 0.8011, 0.84453, 0.88125, 
    0.9121, 0.93766, 0.95849, 0.97495, 0.98743, 0.9958, 1 ;

 pk = 1, 2.69722, 5.17136, 8.89455, 14.2479, 22.07157, 33.61283, 50.48096, 
    74.79993, 109.4006, 158.0046, 225.4411, 317.8956, 443.1935, 611.1156, 
    833.7439, 1125.834, 1505.208, 1993.158, 2614.863, 3399.784, 4382.062, 
    5600.87, 7100.731, 8931.782, 11149.97, 13817.17, 17001.21, 20775.82, 
    23967.34, 25527.65, 25671.22, 24609.3, 22640.51, 20147.13, 17477.63, 
    14859.86, 12414.93, 10201.44, 8241.503, 6534.432, 5066.179, 3815.607, 
    2758.603, 1880.646, 1169.339, 618.4799, 225, 10, 0 ;

 sftlf =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01177494, 
    0.2004458, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01095872, 0, 0.003575196, 0, 
    0.04133711, 0.4170527, 0.86152, 0.830821, 0.6877613,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1264342, 0.5097121, 0.8753754, 
    0.7817355, 0.2817629, 0.5366528, 0.9293424, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1668709, 0.9869201, 1, 1, 1, 
    0.9988317, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.06910358, 0.8185359, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.08511406, 0.7756319, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.5162452, 0.9977401, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.3129568, 0.9959389, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.02861756, 0.6951866, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1453591, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1453354, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.6664422, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0.02644386, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.175007, 0.9126859, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1,
  0.6233622, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2911646, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1,
  0.6379205, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.7788954, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1,
  0.6378774, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.005386431, 0.309769, 0.4789902, 
    0.1082563, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.7179049, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0.6374285, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01172521, 1, 1, 0.7862632, 
    0.2317922, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.6998634, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0.06200648, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2357621, 1, 1, 1, 0.9253088, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.8606739, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.5966171, 1, 1, 1, 0.9915225, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.519107, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1,
  0.3754489, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.5966566, 1, 1, 1, 0.9932248, 
    0.07400899, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.2909555, 1, 0.9996659, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0.9468521, 0.2389454, 0, 0, 0, 0, 0, 0, 0, 0, 0.1795021, 1, 1, 1, 1, 
    0.5510066, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1121078, 
    0.2244427, 0.2677908, 0.8841233, 0.9811913, 0.7802478, 0.9785666, 
    0.8345276, 0.9690673, 0.8673143, 1, 1, 1, 1,
  1, 0.9377849, 0.1510155, 0, 0, 0, 0, 0, 0, 0, 0.004869109, 0.7091162, 1, 1, 
    1, 0.7690508, 0.04686088, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.08630638, 0.05072459, 0.00715183, 0.05010708, 0.0435742, 
    0.04084156, 0.4005074, 1, 1, 1, 1,
  1, 1, 0.5535783, 0, 0, 0, 0, 0, 0, 0, 0.0003298247, 0.4347998, 1, 1, 1, 1, 
    0.1105905, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.1101263, 0.8236522, 1, 1, 1,
  1, 1, 0.9985871, 0.7174072, 0.04896508, 0, 0, 0, 0, 0, 0.0117381, 
    0.9759874, 1, 1, 1, 1, 0.5814301, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.5950869, 0.9525636, 
    0.9839157, 1,
  1, 1, 1, 1, 0.9804606, 0.1933275, 0, 0, 0, 0, 0.01173972, 1, 1, 1, 1, 1, 
    0.6657338, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.0211766, 0.02256984, 0.21058, 0.6582654,
  1, 1, 1, 1, 1, 0.8694932, 0.1387404, 0, 0, 0, 0.01174129, 1, 1, 1, 1, 1, 
    0.9328697, 0.1643069, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.3509133,
  1, 1, 1, 1, 1, 1, 0.8173901, 0, 0, 0, 4.984859e-05, 0.3204487, 0.9584024, 
    1, 1, 1, 1, 0.3567966, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 0.8408963, 0, 0, 0, 0, 0, 0.2506884, 0.7998602, 1, 1, 1, 
    0.7708181, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 0.8408804, 0, 0, 0, 0, 0, 0, 0.002590244, 0.3868952, 1, 
    1, 0.9516376, 0.2383268, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 0.8408653, 0, 0, 0, 0, 0, 0, 0, 0.00495693, 0.7948567, 1, 
    0.7986782, 0.05182758, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 0.8408509, 0, 0, 0, 0, 0, 0, 0, 0, 0.2693094, 0.9602194, 
    0.7707613, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 0.8408375, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.6405759, 
    0.6084861, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 0.8408248, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01842676, 
    0.01816703, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.004960603, 0, 0, 0, 0.4832949, 0.5081044,
  1, 1, 1, 1, 1, 0.822592, 0.252383, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1190309, 
    0.4765593, 0.5912097, 0, 0, 0, 0.1877966, 0.5820142,
  1, 1, 1, 1, 1, 0.6266645, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.07368479, 0, 
    0.06970806, 0.1497295, 0.2323898, 0.3694812, 0.09263787, 0.1388984, 
    0.02827013, 0,
  1, 1, 1, 1, 1, 0.6266469, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01073292, 0.03063297, 0.5991629, 
    0.6986423, 0.8001084, 0.4512461, 0.2554947, 0.185261, 0.05334708, 0, 
    0.08976555, 0.01147698, 0,
  1, 1, 1, 1, 1, 0.6266309, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.04137734, 0.2410906, 0.3296587, 0.6321196, 
    0.8407705, 0.5324757, 0.1355897, 0.1754358, 0.02694144, 0.0008469501, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 0.3423578, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.005920551, 0.2284444, 0.6276525, 0.7197345, 0.8359697, 1, 
    1, 0.8431623, 0.505213, 0.04540349, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 0.01733314, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.284229, 0.6896634, 1, 0.8693293, 0.349668, 0.3810897, 
    0.6086794, 0.240112, 0.01585283, 0.1599976, 0, 0, 0, 0, 0, 0, 0, 
    1.805722e-05, 0, 0.03666643, 0.119504, 0, 0,
  1, 1, 1, 1, 1, 0.03475345, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.1117143, 0.4876121, 0.4447544, 0.2373162, 0.01928726, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.7862673, 0.3681437, 0.1774964, 0.787069, 
    0.4654977, 0, 0,
  1, 1, 1, 1, 1, 0.6265825, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.3158722, 0.9526677, 0.9008846, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.8407551, 0.3746317, 0.4537332, 0.9686775, 0.3652169, 0, 0,
  1, 1, 1, 1, 1, 0.8866345, 0.1598364, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.03936394, 0.6387691, 0.9943234, 1, 0.9008874, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.01252412, 0.4860564, 0.5318119, 0.2620075, 0, 0, 0.1320914, 
    0.8908585, 0.3907566, 1, 0.8389638, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 0.4656247, 0.0110646, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.6010675, 1, 1, 1, 0.9167563, 0.07269689, 0.2391122, 0.2968679, 0, 
    0.2234619, 0.3493941, 0.8015904, 0.8455765, 0.9577049, 1, 1, 0.4179517, 
    0, 0, 0.4412683, 1, 0.6472766, 1, 0.3203639, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 0.6503397, 0.01531898, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.2558588, 0.9597831, 1, 1, 0.972702, 0.9489372, 0.4348444, 0.1722408, 
    0.04735889, 0, 0.7706258, 1, 1, 1, 1, 1, 1, 0.5972056, 0, 0, 0.1294438, 
    0.8859251, 1, 0.8678412, 0.2493258, 0.1075096, 0.1135316, 0.3466776,
  1, 1, 1, 1, 1, 1, 1, 1, 0.287686, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1325035, 0, 
    0.8317441, 1, 1, 0.9539555, 0.2448101, 0.2613218, 0, 0, 0.1152575, 
    0.2170084, 0.900425, 1, 1, 1, 1, 1, 1, 0.8761324, 0.1775864, 0, 0, 
    0.8103314, 0.4596019, 0.6510904, 0.7820377, 0.592761, 0.06109875, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 0.920251, 0.1775966, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.3923621, 0.987651, 1, 1, 0.3509198, 0.2281306, 0, 0, 0, 0, 0.7061847, 
    1, 1, 1, 1, 1, 1, 1, 1, 0.7719379, 0, 0, 0.6054041, 0, 0, 0.02613228, 
    0.1559717, 0.01388168, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 0.7677791, 0.09293438, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.1779837, 0.3241267, 0.9822798, 1, 1, 0.9843383, 0.2598756, 0.01625016, 
    0, 0, 0, 0, 0.866449, 1, 1, 1, 1, 1, 1, 1, 1, 0.8224034, 0.07974907, 0, 
    0.2945428, 0.6333175, 0.5063159, 0.446091, 0.3369552, 0.4868954, 0.174956,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9503866, 0.2001637, 0.005799863, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.1038464, 0.6664168, 1, 1, 0.8380957, 0.2760953, 0.4406356, 
    0.1536544, 0, 0, 0, 0, 0.8664498, 0.9701261, 0.9560779, 1, 1, 1, 1, 1, 1, 
    1, 0.9252388, 0.3537527, 0.03041064, 0.3419223, 0.4810721, 0.4459109, 
    0.1816519, 0.1972405, 0.5183649,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.6181571, 0.04856747, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.6580371, 1, 0.8227324, 0.4224875, 0.510656, 0.9363688, 0.6996492, 0, 0, 
    0, 0, 0, 0.1081687, 0.109901, 0.5228179, 1, 1, 1, 1, 1, 1, 1, 0.3901491, 
    0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8356921, 0.1330075, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.005403113, 
    0.4351665, 0.9745526, 0.7136913, 0.2152697, 0.3135631, 0.9907392, 1, 
    0.2640299, 0, 0, 0, 0, 0, 0, 0, 0.03659684, 0.3494267, 0.8000365, 
    0.9991509, 1, 1, 1, 0.8337656, 0.1029233, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8476309, 0.1004762, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002844633, 
    0.6518675, 1, 0.7256781, 0.03523427, 0, 0.6580248, 1, 1, 0.2640252, 0, 0, 
    0, 0, 0.3051819, 0, 0, 0, 0, 0, 0.8034117, 1, 1, 1, 0.9529892, 0.2843654, 
    0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.7001464, 0.03844476, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.1336879, 0.05886054, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.2070477, 0.4348271, 0.2998562, 0.06389595, 0, 0.1970171, 0.9302663, 1, 
    0.8744631, 0.138245, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1508173, 0.772752, 
    0.9572471, 1, 1, 0.8470377, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.3652858, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 0.7193018, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.5087034, 0.9593135, 0.7576354, 0.1099733, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.318427, 0.9950952, 1, 0.9854341, 0.3656026, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.7283692, 0.04570163, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.06553631, 0.005726846, 0, 1, 0.448386, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.2178526, 0.8641504, 0.4405744, 0.03868152, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.7589623, 0.9413608, 0.3499206, 
    0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.5236878, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.2793671, 0.9727733, 0.3410493, 0.004538658, 0.9128425, 0.1045216, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2580416, 0.9425887, 0.64642, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1441312, 0.3183418, 0, 
    0, 0, 0, 0.1504084, 0.08207643, 0, 0.1264589, 0.6360483,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8886915, 0.171717, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.4181546, 1, 1, 0.2572959, 0.09995186, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.2655529, 0.9644211, 0.5325517, 0, 0, 0, 0, 0.09022734, 
    0.2022693, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.5111119, 0.0366355, 0.2737309, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.7781987, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0143113, 
    0.8599525, 1, 1, 0.8562455, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.1380162, 0.923599, 0.1353773, 0, 0, 0, 0.03968213, 0.2221394, 
    0.7275295, 0.3227897, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1441023, 
    0.2176893, 0, 0, 0, 0, 0.1160006, 0.885816, 0.6751633, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8664993, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.4873159, 
    1, 1, 1, 0.68866, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.1955505, 0.939324, 0.3395239, 0, 0, 0.1328799, 0.7831334, 1, 1, 
    0.7539828, 0.4905147, 0.03082606, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.04012534, 
    0.5083878, 0, 0, 0, 0, 0, 0.1388984, 0.256223, 0.6417912,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9953002, 0.5326272, 0.519923, 0.4552467, 
    0.5700993, 0.8583444, 0.7375726, 0.923451, 0.9061459, 0.1658801, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1702366, 
    0.9217622, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1872573, 0, 
    0, 0, 0, 0.3864902, 1, 0.6463704, 0, 0.1308702, 0.7559305, 1, 1, 1, 1, 1, 
    0.8225404, 0.1237965, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.084927, 0.5631165, 
    0.1094015, 0, 0, 0.08819825, 0.6943044, 0.07551906, 0.006831904,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.4421961, 0, 0, 0, 0, 0, 0, 0.01769246, 
    0.1738239, 0, 0, 0.1787293, 0.04062913, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.3148586, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0808153, 0.9058402, 0.6547354, 0.2428028, 
    0.7843866, 1, 1, 1, 1, 1, 1, 1, 0.6807549, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.2588764, 0.1009072, 0, 0, 0.2429036, 0.7849156, 0.4656103, 0.169591,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9108992, 0.188346, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.7856974, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.3914096, 1, 1, 0.9854771, 1, 1, 1, 1, 1, 1, 1, 1, 0.6807355, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.7825689, 0.6956174, 0.09677283, 
    0.1274765,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 0.7852127, 0.4266168, 0.8433919, 0.4879982, 
    0.2553098, 0.4059382, 0.1131723, 0.02167348, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2218162, 0.963348, 1, 1, 
    1, 1, 1, 0.688597, 0.09377675, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.01462167, 0.002184577, 0, 0, 0.8908938, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 0.3777061, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.003051978, 
    0.07014503, 0.1355046, 0.1359438, 0.006367458, 0.6373758,
  1, 1, 1, 1, 1, 1, 1, 1, 0.8328858, 0.2307329, 0.8818867, 1, 1, 1, 1, 1, 
    0.691934, 0.4109589, 0.2119478, 0.1284744, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.5544662, 1, 1, 1, 1, 1, 1, 1, 
    0.946013, 0.1113746, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.3114816, 0.7581814, 
    0.5352249, 0.1977297, 0.9311432, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.1334493, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.181796, 0.5997484, 0, 0, 
    0.3158956, 0.500448,
  1, 1, 1, 1, 1, 1, 1, 1, 0.1062542, 0.1823296, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.9209124, 0.0554863, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.7544572, 1, 1, 1, 1, 1, 1, 1, 1, 0.9121619, 0.5140178, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.8938125, 1, 0.7836286, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 0.9445137, 0.6255063, 0.02327494, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.316875, 0.3196791, 0.2422916, 0.0662774, 0.6194771, 0,
  1, 1, 1, 1, 1, 1, 0.8702384, 0.2501028, 0.005983606, 0.5771939, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 0.8631834, 0.8403694, 0.5729032, 0.2040605, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.00724657, 0.7643476, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0.9984289, 0.3873025, 0, 0, 0, 0, 0, 0, 0, 0, 0.2322503, 
    0.9433986, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9763494, 0.1368165, 
    0.0004370618, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1078297, 0.7730162, 
    1, 0.6829644, 0.4463389, 0.2076392, 0.1887735,
  1, 1, 1, 1, 1, 0.8587388, 0.1308349, 0, 0, 0.4788192, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 0.9391835, 0.775203, 0.1979599, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.239585, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9413478, 
    0.3537645, 0.05398361, 0, 0, 0, 0, 0, 0, 0.8853288, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0.9915676, 0.4714071, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.2355691, 1, 0.7928132, 0.1206847, 0, 0, 0,
  1, 1, 1, 1, 1, 0.4860172, 0, 0, 0, 0.7716876, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0.9360449, 0.2212868, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.1080709, 0.2082748, 0.2002707, 0.8915246, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 0.6313275, 0, 0, 0, 0, 0.0001691831, 0.5004879, 0.9755507, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 0.6524076, 0, 0, 0.2558733, 0.5018113, 0.2678142, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.136077, 0.8694932, 0.7911853, 0.08738397, 
    0, 0, 0,
  1, 1, 1, 1, 1, 0.01735635, 0, 0, 0.1874817, 0.9048839, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 0.5105418, 0.01035661, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.1085859, 0.8962955, 1, 0.9106531, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 0.8520856, 0.3672015, 0.313609, 0.2533256, 0.03519395, 0.3614787, 
    0.9965006, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9207106, 0.068037, 0, 
    0.3333627, 0.9408049, 0.8420026, 0.07602482, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.6269207, 1, 0.3631722, 0, 0, 0,
  1, 1, 1, 1, 0.7065716, 0.007449343, 0, 0, 0.8899581, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9990095, 0.6469289, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.302171, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 0.2509532, 0.7259984, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.4962145, 0.009399206, 0, 0.163563, 0.8311784, 0.2532057, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.6269538, 1, 0.7403622, 0, 0, 0,
  1, 1, 1, 0.9591063, 0.2903444, 0, 0, 0.3821371, 0.9899979, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8423643, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.1113189, 0.9288797, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 0.9148951, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.7166897, 0.193198, 0.378679, 0.7709084, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.2623808, 0.6417641, 0.1763478, 0, 0, 0,
  1, 1, 1, 0.4600145, 0, 0, 0.06470905, 0.7741343, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9729096, 0.4085401, 0, 0, 0, 0, 0, 0, 0, 
    0.09763272, 0.8372439, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.8914483, 0.9574527, 0.9569234, 0.6728632, 0.2309492, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 0.9083645, 0.1139706, 0, 0.006719753, 0.6425024, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.6623873, 0.3399824, 0, 0, 0, 0, 0, 
    0.01343901, 0.1122996, 0.2740395, 0.8126243, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9409829, 0.4917598, 0.01190909, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 0.5350372, 0, 0, 0.3691856, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.9817434, 0.7555508, 0.5806262, 0.721405, 0.9975661, 0.7792664, 
    0.03027645, 0, 0.05746033, 0.4528793, 0.6003847, 0.7402431, 0.8724493, 
    0.9833708, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0.9409539, 0.3217609, 0.0036727, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  1, 1, 0.5350789, 0, 0, 0.8339525, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.5068051, 4.62555e-05, 0, 0.01343513, 0.4826073, 0.6908599, 0.1210046, 
    0.6430895, 0.8287125, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9063402, 0.1092877, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 0.5351219, 0, 0, 0.9826248, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.6957842, 0.4102102, 0, 0, 0, 0.04356555, 0.1127979, 0.72868, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 0.9970281, 0.3331997, 0, 0, 0, 0.3913397, 0, 0, 
    0, 0, 0,
  1, 0.952481, 0.2011694, 0, 0, 0.9826218, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.8811629, 0.2063091, 0.1352319, 0.007285898, 0.3884326, 0.8899049, 
    0.8934386, 0.7892479, 0.9770009, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.9107391, 0.1889964, 0, 0.1838041, 0.8709035, 0.1881444, 0, 0, 0, 0,
  0.9999014, 0.380338, 0, 0, 0.4566294, 0.9974383, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 0.6904973, 0.03093301, 0.01432722, 0.6824431, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8582283, 0.03906883, 0.08034394, 
    0.7920045, 0.5992478, 0, 0, 0, 0,
  0.6594298, 0, 0, 0.3033189, 0.9943448, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.8270786, 0.08996841, 0.002212425, 0.4717253, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.7097963, 0.03884534, 0.4686598, 
    0.7735896, 0.07057529, 0, 0, 0,
  0.6233622, 0, 0.156587, 0.9117836, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.4757935, 0, 0.1331947, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 0.4924225, 0.007284605, 0.6021019, 0.1786143, 0, 0, 0,
  0.02644386, 0, 0.4743553, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9506161, 
    0.08966529, 0.03939142, 0.6957731, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8284553, 0.06092081, 0, 0, 0, 0, 0,
  0, 0.07934966, 0.98106, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.5513756, 0, 
    0.5253358, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 0.3725595, 0, 0, 0, 0, 0,
  0, 0.4350433, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9976279, 0.3553158, 
    0.6696817, 0.9791158, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 0.8894136, 0.02892898, 0, 0, 0, 0,
  0.01680065, 0.7740205, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9978701, 
    0.8976342, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 0.5902183, 0, 0, 0, 0,
  0.5105151, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8744972, 
    0.1220256, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9973416, 
    0.2167705, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9901414, 0.2867822, 
    0.3897793, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.816124, 
    0.1255585, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9809267, 0.9553849, 
    0.3948242, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.2193899, 0.1200667, 0, 
    0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.4875835, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.1584725, 0, 0, 0, 0, 0, 0,
  0.5802633, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.6097519, 0, 0, 
    0, 0, 0, 0,
  0.08221136, 0.7452577, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9897885, 
    0.9358599, 0.9987948, 0.7364435, 0, 0, 0, 0, 0,
  0, 0.7250001, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9684403, 0.774133, 
    0.3314505, 0.8281783, 0.9904674, 0.221187, 0, 0, 0, 0 ;

 orog =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.007482118, 
    4.885016, 6.027729, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.712759, 58.8956, 
    114.3027, 105.147, 66.36284,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.754428, 58.17822, 103.8941, 
    76.19964, 51.16923, 83.5846, 145.4227, 210.3575, 222.043, 166.9021, 
    138.0394,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12.60223, 150.9446, 238.0754, 281.3481, 
    288.7326, 300.3335, 276.3248, 277.1753, 296.433, 282.2253, 207.1847, 
    170.1954,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.971491, 107.903, 253.5528, 311.8893, 
    314.664, 349.46, 376.1395, 363.9048, 328.7521, 316.8185, 308.9201, 
    249.6144, 213.1554,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1077713, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.728832, 54.67075, 280.7457, 
    309.0462, 322.4052, 368.6298, 412.7725, 423.5071, 379.2067, 346.22, 
    351.7698, 329.3646, 274.3772,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.078801, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17.70223, 257.5212, 295.4054, 
    313.6127, 373.5954, 422.1055, 435.1128, 393.682, 374.0881, 409.6835, 
    409.2048, 354.9377,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26.2593, 246.0138, 296.1431, 348.5571, 
    410.7598, 429.6357, 435.3861, 395.7879, 402.5177, 442.4218, 430.7854, 
    398.5805,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 113.7163, 268.1346, 336.5029, 392.1589, 
    444.2632, 443.9155, 420.9473, 421.8472, 452.1077, 471.5658, 444.4251, 
    418.9319,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.859579, 200.0244, 305.7336, 330.6553, 
    391.9315, 444.2378, 439.8025, 441.541, 463.3921, 503.8092, 497.416, 
    462.6526, 441.0611,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14.25746, 228.6333, 312.2241, 361.2495, 
    416.0756, 482.3185, 484.5522, 484.6867, 507.3547, 509.7314, 483.8749, 
    461.7263, 442.7195,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.007934935, 91.5881, 260.8788, 351.2304, 
    404.0062, 456.2148, 509.2211, 528.7908, 527.3947, 511.4882, 494.72, 
    462.9256, 467.0975, 450.041,
  7.299402, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8.026843, 190.214, 291.695, 351.6114, 
    434.4432, 470.4533, 537.1084, 567.7097, 561.1059, 537.2833, 494.2285, 
    457.0371, 454.9888, 443.677,
  46.47058, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32.85493, 192.2326, 276.3241, 346.8046, 
    419.9743, 473.221, 539.5166, 587.4988, 579.1885, 551.3723, 502.3163, 
    438.6668, 426.6781, 416.2831,
  56.36044, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2935236, 29.53243, 141.496, 253.5633, 
    345.4431, 426.5362, 485.1349, 548.7592, 600.852, 588.0337, 535.9756, 
    460.5315, 394.231, 382.3351, 380.9086,
  39.45049, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32.83228, 53.73461, 1.585332, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3.041326, 10.00888, 
    106.9153, 227.8007, 348.7626, 445.4996, 478.5939, 575.4977, 600.4197, 
    570.2203, 506.0541, 415.3415, 330.4285, 332.2667, 343.1945,
  13.59347, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26.08635, 195.4105, 256.4257, 146.537, 
    55.481, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.186994, 
    18.06586, 130.0469, 253.3653, 363.8199, 394.896, 513.6748, 590.4353, 
    558.9642, 518.7917, 454.3615, 363.8717, 303.3865, 300.713, 321.3069,
  0.9656757, 0, 0, 0, 0, 0, 0.03586638, 0, 0, 0, 49.68565, 326.9774, 
    455.3936, 576.6316, 425.3625, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.01508173, 21.43529, 144.3786, 255.7441, 319.1965, 459.2542, 
    569.7118, 604.0175, 513.782, 425.8328, 371.0454, 316.678, 281.3964, 
    295.9887, 312.7417,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 188.9793, 461.0893, 744.1964, 857.3239, 
    577.0432, 10.22077, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    28.41998, 89.48728, 170.1808, 341.458, 487.3284, 552.6357, 471.7288, 
    351.3307, 336.5912, 295.8323, 257.3056, 256.7657, 275.5327, 266.8901,
  14.46666, 0, 0, 0, 0, 0, 0, 0, 0, 0, 98.10371, 430.0524, 658.2639, 
    869.6558, 593.5727, 27.91763, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 28.79319, 27.47902, 102.3828, 250.1567, 353.9292, 297.6356, 
    194.349, 196.082, 204.2073, 194.9052, 184.4335, 186.8029, 202.2491, 
    201.6232,
  63.77672, 3.367655, 0, 0, 0, 0, 0, 0, 0, 0, 20.47009, 226.3262, 481.9063, 
    847.3206, 850.9589, 97.98926, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 5.864242, 1.030459, 11.5586, 92.8717, 81.6533, 37.3248, 
    45.25832, 55.12968, 71.40536, 80.22321, 109.8221, 156.4528, 158.7244, 
    139.6773,
  92.77831, 10.55024, 0.7231424, 0, 0, 0, 0, 0, 0, 0, 0.06683189, 88.24445, 
    325.958, 897.7953, 1142.866, 334.1817, 0.2153307, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.6444512, 1.022004, 0.2444094, 0, 
    0.1744056, 0, 0, 11.61093, 95.71937, 140.5593, 109.8717, 89.47809,
  148.8612, 111.2776, 10.43683, 0.2487843, 0, 0, 0, 0, 0, 0, 0, 26.9947, 
    302.4542, 900.6857, 1410.459, 722.3347, 26.92253, 0, 0, 0, 0, 0, 0, 
    0.2948902, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.04675792, 32.30137, 73.17574, 45.04506, 113.3446,
  356.8611, 272.9169, 144.0292, 36.66886, 4.051232, 0, 0, 0, 0, 0, 
    0.00622688, 95.44665, 402.4702, 1000.551, 1468.909, 1068.681, 138.7007, 
    0, 0, 0, 0, 0, 0, 224.4563, 0.7204035, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 40.79513, 46.98636, 44.90553, 135.4555,
  607.5697, 617.0065, 415.9779, 222.5245, 82.16385, 13.76159, 0, 0, 0, 0, 
    0.7036354, 167.195, 549.0036, 865.797, 1297.997, 1084.883, 386.271, 0, 0, 
    0, 0, 0, 0, 0, 0, 38.47579, 1.349345, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.05735796, 3.489815, 17.0652, 91.46315,
  805.8144, 689.3148, 665.8074, 521.1199, 295.9792, 99.36646, 9.087084, 0, 0, 
    0.005802704, 0.3102686, 111.6922, 363.4742, 565.2116, 806.0615, 1016.094, 
    629.3563, 16.26268, 0, 0, 0, 0, 0, 0, 0, 0, 0.02296036, 0, 0, 0, 0, 
    1.214581, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002000303, 0.005462797, 
    18.32721,
  760.7727, 661.396, 709.6733, 604.6326, 464.2514, 283.1679, 79.76301, 
    0.1074248, 0, 0, 0, 17.74922, 148.9407, 173.6682, 402.7549, 729.6694, 
    723.2713, 46.89246, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1074003,
  860.9228, 736.6833, 628.5461, 564.9741, 466.655, 335.0508, 169.4657, 
    9.562907, 0, 0, 0, 0, 7.39888, 15.74615, 103.3149, 461.4926, 652.2623, 
    214.472, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, -0.0001159482, 0, 0,
  954.5076, 825.0037, 642.887, 541.5004, 467.5988, 374.7963, 167.8485, 
    1.774008, 0, 0, 0, 0, 0, 0.3348222, 19.11695, 171.6814, 741.9515, 
    374.4197, 25.98872, 0, 0, 0, 0.0003252521, 0, 0, 0, 0, 0.001458651, 
    7.516816e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  858.3884, 673.0359, 533.1504, 448.0885, 424.8119, 345.4697, 166.7318, 0, 0, 
    0, 0, 0, 0, 0, 0.567318, 193.9483, 883.2621, 655.3737, 12.50792, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.0002288724, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.005102882, 0, 0,
  765.3333, 667.6134, 488.7987, 363.019, 313.4333, 341.2213, 122.4717, 0, 0, 
    0, 0, 0, 5.00687, 0, 0, 60.76902, 616.8209, 406.96, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  892.0968, 795.8924, 625.4323, 432.2025, 321.9835, 331.9277, 130.2014, 
    0.004251794, 0, 0, 57.24534, 20.8572, 0.7291545, 0, 0, 0, 119.2905, 
    99.81622, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 13.85986, 0.004370535, 0,
  1001.771, 792.1298, 674.5222, 541.9408, 384.3335, 350.6531, 103.3347, 
    0.1868827, 0, 0, 18.48727, 0, 0, 0, 0, 0, 9.2637, 4.286283, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.02841037, 
    1.063279, 1.850597, 3.574715, 3.295839, 153.8647, 199.7177,
  1318.781, 598.8708, 526.7117, 510.9486, 354.2004, 223.6784, 15.55483, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.01238247, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10.38296, 174.51, 148.3694, 0, 0, 0, 
    148.5062, 285.8834,
  1220.16, 848.2032, 380.6071, 390.465, 259.5177, 95.94141, 0, 0, 0, 0, 0, 0, 
    0, 0.01723676, 0.0002739781, 0.009286015, 0, 0, 0, 0.006633122, 0, 0, 0, 
    0, 0.003201818, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001933358, 
    0, 0, 0, 0, 0, 0, 0, 0, 2.528343, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.01048129, 0, 35.29255, 81.26061, 161.3701, 172.8166, 125.7769, 
    60.08969, 51.96622, 164.8291,
  1338.663, 964.2402, 591.19, 291.6062, 139.8224, 33.77381, 0.002896692, 0, 
    0, 0, 0, 0, 0, 0.09759907, 0, 0, 0, 0, 0.003041361, 0, 0, 0, 0, 0, 
    0.003417519, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.214117, 10.05566, 31.4626, 
    198.6635, 257.3435, 200.3842, 110.9841, 79.73378, 263.6654, 36.78745, 
    1.378057, 31.15954, 8.130059, 1.005422,
  1026.086, 1045.23, 716.394, 366.1234, 142.9799, 30.33171, 0.4619157, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10.88786, 
    115.5257, 170.2808, 339.2503, 395.8933, 151.5352, 149.8366, 27.3561, 
    4.022614, 20.95062, 0, 0, 3.260029, 1.872875, 0.0508271, 0, 0, 0,
  974.4459, 1067.982, 927.8552, 494.0284, 130.0466, 22.65291, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.899872, 139.8198, 
    115.3161, 168.5896, 352.7554, 266.0829, 177.1721, 131.6926, 43.10759, 
    1.240668, 4.394837, 0.006916575, 0.0003986534, 0.0104446, 0.0172614, 0, 
    2.609623, 0, 0.001365404, 0.09803439, 0.2262536, 0.004817449,
  1204.486, 1237.256, 1141.603, 688.0075, 263.0531, 10.36784, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001947393, 0, 0, 0, 0.01043915, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01680503, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.04407993, 32.09272, 400.8964, 597.5397, 333.6716, 124.2354, 104.7639, 
    67.59129, 23.81756, 3.731113, 1.087241, 0, 0, 0, 0, 0, 0, 4.881635, 
    10.31701, 0, 6.561506, 40.6811, 3.38201, 0.01358287,
  1440.196, 1303.7, 1187.572, 799.9657, 447.4943, 28.87032, 0.287935, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.008367683, 0, 0.0005597501, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.006913288, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 17.87501, 27.6564, 41.68385, 40.07766, 2.412819, 0, 0.3703949, 0, 0, 
    2.694052, 0, 0.06298108, 0, 0, 0.007401017, 0.01018163, 0.5245222, 
    314.3598, 25.13958, 10.84065, 64.80965, 69.94651, 0.2126305, 0,
  1507.507, 1338.634, 1162.16, 895.2739, 556.3425, 113.5388, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.003531589, 0, 0.3608332, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.645804e-05, 0.008660849, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.399279, 1.708197, 228.0259, 260.7763, 73.72216, 0.01350134, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.04154294, 0.6853305, 0.0007041242, 0, 0, 0, 222.6289, 
    19.51247, 152.801, 98.75947, 68.60026, 0, 0,
  1593.552, 1288.948, 1293.234, 1037.663, 604.3491, 220.0716, 11.92896, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3.231213, 0.1002754, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.003929192, 0.06615317, 
    326.9998, 382.6881, 215.296, 6.51867, 0, 0, 0.0005210711, 0, 0, 0, 
    0.00945402, 0, 0.04497931, 26.08819, 57.13885, 7.390703, 0, 0, 69.87069, 
    559.0273, 111.9894, 624.2891, 262.6683, 1.642632, 0, 0,
  1658.693, 1261.843, 1404.586, 1067.003, 563.8726, 182.1493, 36.27239, 
    0.3323672, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002778716, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3.277349, 3.089526, 
    220.2578, 271.9154, 232.9942, 11.41514, 6.090748, 2.68348, 5.510962, 
    3.529593, 0, 1.621469, 5.491666, 9.77548, 7.35185, 3.514773, 53.89715, 
    161.2589, 24.12606, 0, 0.007201126, 433.8056, 1036.646, 400.0064, 
    500.544, 149.6249, 0, 0, 0,
  1645.619, 1472.14, 1404.025, 1096.18, 483.7211, 188.2313, 50.92135, 
    15.02244, 0.3012842, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9.016459, 125.5137, 
    477.9677, 315.6645, 11.36371, 6.38086, 10.82686, 9.825094, 2.584005, 
    0.8772991, 0, 14.4698, 70.73858, 64.99486, 20.69061, 17.08455, 32.61346, 
    164.0018, 34.12597, 0.002215982, 0, 41.34579, 1159.648, 903.4078, 
    550.6257, 25.76042, 12.09169, 7.678148, 124.0715,
  1967.175, 1791.275, 1808.567, 1089.094, 523.5789, 218.3327, 97.51249, 
    52.39918, 11.84871, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26.70954, 0.01252906, 
    573.1802, 456.6572, 67.73898, 16.5005, 4.31343, 5.305326, 0.0450154, 0, 
    0.8252385, 6.159415, 65.49741, 194.1909, 179.5106, 157.9093, 77.64091, 
    91.67677, 141.2131, 99.64323, 8.659935, 0, 4.571824, 614.8233, 532.0992, 
    483.2188, 457.6458, 209.052, 8.435591, 0,
  2024.533, 2181.229, 2001.106, 1283.735, 528.7686, 242.7618, 136.9167, 
    79.82225, 23.44122, 3.95113, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.004921097, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.6401625, 
    6.308005, 158.2323, 422.013, 185.8305, 17.01043, 4.866463, 8.841109, 
    0.001300426, 0, 0, 0, 11.91, 84.76138, 176.0108, 242.7657, 291.476, 
    330.5183, 200.2534, 138.5459, 34.58592, 22.24334, 0, 0, 144.1948, 0, 
    6.173299, 15.85019, 45.24471, 0.213134, 0,
  1923.579, 1771.256, 1778.076, 1070.793, 505.6136, 241.9928, 148.163, 
    76.44843, 32.30178, 17.09214, 7.496256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01376197, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.004098975, 22.05864, 72.32189, 406.9106, 296.7709, 13.30871, 10.29677, 
    4.396094, 1.765978, 0, 0.01962267, 0.09792335, 0.3374118, 51.71622, 
    88.17578, 76.92102, 159.3824, 380.0949, 535.228, 499.3378, 330.4606, 
    165.3464, 41.27188, 2.509667, 0.02632017, 117.6165, 245.3032, 188.3384, 
    112.4978, 172.8582, 310.4585, 94.6843,
  1794.133, 1276.998, 1319.927, 847.228, 358.8172, 233.8158, 187.9514, 
    116.8452, 68.52618, 71.37233, 45.78811, 16.83432, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.009340961, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2.670939, 25.97792, 355.1271, 272.5902, 27.50756, 10.82965, 
    10.10394, 20.80869, 2.207196, 0, 0.004632319, 0.4954259, 0, 54.69146, 
    103.1393, 87.46021, 162.231, 378.5865, 622.8563, 789.714, 748.1737, 
    514.2153, 211.2245, 106.0069, 43.93421, 0, 117.153, 217.9034, 176.2699, 
    56.00568, 72.75879, 291.925,
  1122.184, 817.0998, 942.5208, 629.3625, 367.3386, 319.362, 310.6506, 
    233.7132, 219.4219, 172.6176, 170.9612, 87.88506, 52.56012, 6.837942, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.01282556, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.003567874, 9.907857, 7.509503, 341.4931, 669.8797, 266.7873, 
    11.2073, 57.75204, 56.43156, 49.87582, 0.7429065, 0.01104457, 0.2828173, 
    0, 0.04069449, 4.1862, 0.06066301, 11.07728, 86.06728, 187.3697, 
    479.2986, 762.8614, 937.4857, 601.6578, 195.3882, 27.83612, 0.1914168, 0, 
    0, 0, 0, 0, 0, 11.51637,
  846.5782, 504.4499, 654.7703, 570.2628, 501.0254, 542.6677, 483.9015, 
    424.1021, 332.9808, 314.234, 333.5416, 253.9334, 130.1149, 111.9619, 
    7.31144, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.0009155833, 0.003754308, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.204808, 504.0269, 598.7817, 428.9163, 
    11.3934, 12.47365, 231.9589, 136.3775, 6.838151, 0, 2.634708, 3.781463, 
    0.1162148, 0.6912898, 0.01993117, 0, 0.4706172, 7.387184, 44.55817, 
    244.1146, 594.9794, 933.8558, 513.5035, 77.61767, 4.361522, 0, 0, 0, 0, 
    0, 0, 0, 0,
  681.6527, 442.5084, 578.8173, 717.4026, 922.1249, 813.6738, 759.1872, 
    525.2695, 321.9953, 302.5872, 458.9889, 403.1359, 243.0368, 181.6122, 
    107.4319, 9.799197, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.0001312634, 0.006848679, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.3214408, 335.2546, 813.2599, 438.9796, 
    1.541609, 0.004860971, 141.2879, 433.2815, 256.4115, 14.89001, 0, 0, 0, 
    0.1404909, 6.80957, 0, 0, 0, 0, 0.4797853, 35.22785, 388.0224, 854.2148, 
    528.0695, 83.28231, 2.967625, 0, 0, 0, 0, 0, 0, 0, 0,
  545.9903, 500.1561, 701.9286, 1102.757, 1219.171, 1147.172, 956.5318, 
    675.6527, 331.725, 351.9229, 475.9785, 420.0756, 313.623, 228.7287, 
    180.0209, 134.015, 0.3182439, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01651771, 0, 0, 0, 0, 0, 0, 22.53872, 
    0.65847, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30.20723, 195.3939, 
    90.67072, 4.860431, 0, 5.169554, 264.6625, 416.897, 223.7468, 2.467426, 
    0, 0, 0, 0.01299047, 0.1073577, 0, 0, 0, 0, 0, 2.723956, 80.23975, 
    657.4532, 634.125, 285.9821, 125.6809, 2.169004, 0.1452292, 0, 0, 0, 0, 
    0, 0,
  575.7665, 549.1124, 1004.394, 1257.504, 1520.269, 1214.792, 1053.349, 
    760.7601, 506.7095, 417.5125, 432.6968, 399.7943, 364.9707, 304.9736, 
    209.8668, 138.7341, 27.90703, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001978899, 0.02694878, 0, 0, 0, 0, 0, 
    7.94479, 361.0423, 148.2079, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3.387879, 
    0.004412269, 0, 0, 0, 1.012016, 28.95815, 159.6374, 162.7487, 6.871452, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002113436, 123.6737, 502.31, 
    321.5427, 69.19288, 34.57666, 4.016514, 0.6476752, 0, 0, 0, 0, 0,
  771.0378, 731.9822, 1232.212, 1579.218, 1810.72, 1665.98, 1247.325, 
    891.9006, 552.7863, 534.0606, 470.0626, 487.2615, 500.9968, 399.5934, 
    301.6216, 216.2957, 101.2677, 1.366401, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7.578414, 0, 10.02934, 
    217.377, 48.73487, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2398228, 7.076045, 0, 
    0, 0, 0.5435731, 5.565549, 79.59003, 18.13072, 1.341174, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.07269884, 342.0459, 154.1556, 9.21379, 
    0.01240786, 0.0236598, 5.468072, 10.2199, 0.1744068, 0, 0, 1.12455,
  1005.523, 1089.269, 1428.493, 1729.941, 2157.611, 2366.877, 1791.208, 
    1172.936, 789.075, 679.2053, 769.5369, 774.6565, 661.5249, 538.7116, 
    499.1805, 452.9259, 318.8668, 107.7354, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.003257784, 0, 0, 14.33969, 
    269.4527, 18.4388, 2.629723, 63.20306, 3.818854, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.4436082, 0.4391197, 0, 0, 0, 11.42085, 94.30405, 98.075, 
    0.03083581, 0, 0, 0, 0.03971905, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9.149135e-05, 
    0, 0, 9.795963, 11.95197, 0.4926467, 0.0001121615, 0, 0.0542269, 
    0.1652767, 35.90819, 0, 61.54511, 395.5136,
  1443.506, 1620.422, 1765.2, 1789.817, 2168.043, 2356.399, 1999.072, 
    1344.355, 974.863, 966.6523, 1036.74, 970.4948, 807.8265, 729.062, 
    640.0353, 622.3807, 558.9814, 343.8018, 29.92353, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0003971517, 0.002529405, 0, 0, 
    121.7922, 429.6986, 193.016, 6.398975, 3.334329, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.2867806, 0, 0, 0, 0, 3.61325, 129.9913, 54.15724, 0, 0, 0, 
    0.1055335, 0.3423316, 0.3816859, 0.8894814, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3.002282, 0, 0, 0, 0, 0, 91.78906, 15.18766, 64.01128, 362.9198,
  1620.956, 2030.3, 1884.991, 2049.509, 2068.68, 2175.013, 1586.164, 
    1522.586, 1346.341, 1360.391, 1342.486, 1150.649, 1009.675, 798.4236, 
    803.64, 793.613, 751.2167, 539.5749, 185.2117, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.00889502, 0.008948714, 0, 1.305878, 
    327.1373, 460.4203, 183.9435, 19.73282, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.001868226, 3.177953, 0, 0, 0, 0, 5.91536, 94.78001, 1.925256, 0, 0, 
    0.02996243, 4.757724, 2.262005, 0.8893167, 0.6945848, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 38.47111, 40.73141, 0, 0, 0, 0, 68.93193, 198.6472, 
    337.3564, 558.7494,
  1649.085, 1708.983, 1942.575, 2064.672, 2304.163, 2042.305, 1346.739, 
    1341.973, 1536.301, 1614.115, 1351.418, 1085.79, 943.1578, 900.9448, 
    952.3292, 1066.381, 834.631, 657.6016, 280.5684, 3.45371, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001200154, 0.001476862, 0, 
    152.6915, 685.7798, 660.864, 391.5136, 81.102, 0.08322787, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.1983324, 8.214144, 0, 0, 0, 0, 7.976196, 96.0976, 
    32.68804, 0, 0, 11.5986, 136.4807, 24.27074, 1.852875, 7.053572, 
    56.97015, 4.038934, 0.03956408, 0, 0, 0, 0, 0, 9.457328e-05, 0, 0, 
    0.1137195, 89.28968, 12.82965, 0, 0.000534966, 0, 0, 46.44008, 85.76493, 
    411.291,
  1466.144, 1621.266, 1631.515, 2122.453, 2175.795, 2267.993, 1097.97, 
    824.9056, 896.3997, 932.9909, 568.8134, 122.1493, 139.7222, 230.9751, 
    585.2339, 743.4264, 595.6318, 653.7233, 457.3597, 15.86434, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.980672, 440.7948, 
    848.3855, 797.6866, 593.3608, 199.7116, 8.479733, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 11.56622, 0.1151541, 0, 0, 0, 11.44357, 154.1412, 126.2073, 
    0.02027015, 0.8643358, 204.4469, 257.3035, 118.653, 15.25982, 90.17926, 
    348.3282, 451.6818, 20.03893, 0, 0, 0, 0, 0, 0.0003784416, 0, 0, 0, 
    0.3295275, 73.48798, 1.209638, 0.001240408, 0.04867897, 35.55901, 
    205.4684, 37.47905, 55.50045,
  1265.107, 1271.335, 1965.781, 1997.247, 2257.103, 2371.452, 1157.836, 
    568.8094, 507.9307, 527.9256, 61.88685, 0, 0, 0, 0, 0, 0, 0, 25.08505, 
    2.611548, 1.012719, 54.77631, 55.46979, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 56.8435, 558.8643, 753.3204, 685.9753, 529.2399, 
    221.9993, 6.638701, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.390496, 0.1437027, 
    0, 0, 0, 5.025319, 296.0272, 133.192, 26.48146, 105.7203, 124.3082, 
    133.4471, 18.79172, 41.91351, 168.925, 502.5459, 687.1468, 145.1467, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 9.612703, 23.07717, 0.1670243, 0.3258666, 
    40.60841, 178.4189, 98.15704, 58.47993,
  935.9797, 1371.701, 1933.655, 2314.278, 2206.839, 2331.325, 1047.749, 
    519.5513, 454.4148, 405.1205, 26.92118, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 244.4359, 
    576.6982, 579.9873, 438.5885, 334.7599, 131.4858, 3.241302, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.0453538, 0.0158177, 0, 0, 0, 75.12135, 375.2448, 
    88.78672, 19.92136, 145.9868, 126.3988, 55.09162, 79.25726, 93.2966, 
    89.02313, 311.1271, 517.6355, 122.5172, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.03161435, 9.429642, 0.6056394, 0.146424, 207.0213, 126.4081, 45.91529, 
    85.9324,
  705.9424, 1077.602, 1789.276, 2157.059, 2121.644, 2145.599, 927.7297, 
    349.9645, 414.1831, 239.4039, 205.0616, 535.8789, 337.7988, 224.2843, 
    93.21812, 12.07225, 4.108486, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21.81651, 480.2482, 616.3601, 509.2854, 
    411.6318, 353.8981, 172.9756, 23.66262, 1.744636, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.001127199, 0.426254, 0.06272013, 0, 158.0811, 521.639, 
    141.0725, 99.96737, 247.5734, 203.0635, 144.6472, 146.9874, 146.9239, 
    291.5794, 505.7589, 561.468, 82.04576, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7.754673, 7.457764, 24.7692, 42.12467, 9.055123, 4.078703, 80.82257,
  560.522, 873.38, 1472.261, 1866.38, 1992.183, 1959.356, 668.1165, 250.8919, 
    291.7672, 17.91137, 626.5022, 1631.719, 1588.758, 1237.268, 972.5966, 
    822.8162, 666.3598, 231.6238, 95.20377, 24.35091, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 93.28631, 598.2587, 574.9574, 
    508.1927, 475.7988, 445.4901, 244.6739, 75.22868, 59.67073, 26.13394, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 7.006592, 9.506021, 2.820326, 1.543359, 
    144.5288, 485.7056, 157.8752, 139.0608, 306.2983, 182.6353, 140.4857, 
    150.7803, 237.6682, 550.9364, 811.1963, 598.2958, 25.34849, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 140.1268, 241.5589, 39.90154, 11.41144, 38.09826, 
    75.28021,
  520.9725, 685.0739, 1104.142, 1548.977, 1849.273, 1977.533, 530.145, 
    203.5752, 23.72789, 27.13107, 956.7662, 2034.414, 1627.404, 1195.415, 
    1080.397, 1104.885, 1093.357, 887.1946, 732.5614, 442.7809, 42.32203, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 227.5572, 
    614.1383, 604.0764, 532.1347, 527.2681, 501.3772, 266.3045, 197.5267, 
    319.5226, 439.0925, 52.55056, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01218646, 
    68.76542, 10.88835, 49.6851, 244.7333, 434.6059, 156.4234, 331.7645, 
    396.8661, 241.47, 169.5624, 150.5604, 254.91, 544.6859, 578.8292, 
    122.1243, 0.04935317, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.776042, 
    88.48724, 86.04845, 37.06418, 36.67148, 83.62952, 1.168923,
  520.364, 623.9707, 845.1304, 1182.964, 1794.826, 1631.395, 245.3956, 
    30.59338, 0.1295522, 65.68732, 1191.472, 1929.175, 1380.801, 898.722, 
    945.2995, 1004.129, 951.7753, 889.402, 807.7346, 725.3493, 650.4291, 
    576.4832, 399.0143, 189.4995, 1.069616, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 290.6859, 650.6129, 587.6777, 538.5913, 469.5362, 
    367.0397, 239.3359, 267.2038, 520.4188, 582.6263, 354.7753, 95.80848, 0, 
    0, 0, 0, 0, 0, 0, 0, 10.50261, 205.8622, 156.8265, 367.9012, 536.3768, 
    554.2907, 339.4029, 439.8899, 418.0555, 214.6228, 185.1647, 265.1077, 
    310.9288, 294.0193, 49.32493, 0, 0, 0, 0.0004447775, 0.0008141641, 
    0.0001843075, 0, 0, 0, 0, 0, 0.00153388, 0, 9.762164, 91.66759, 151.5858, 
    43.30084, 69.43888, 56.62251, 23.58093,
  527.755, 558.0959, 777.8425, 1038.259, 1442.285, 857.6389, 34.7822, 
    0.06794915, 0.1317989, 65.86896, 1226.782, 1676.783, 1155.866, 959.6856, 
    863.8164, 851.5259, 757.8932, 699.1624, 691.1156, 647.6199, 588.8004, 
    448.2683, 337.8521, 251.0181, 128.1548, 0.6675929, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1.583894, 274.4207, 587.1978, 539.9442, 498.1378, 
    401.8043, 324.701, 235.9535, 351.3758, 472.5636, 586.2536, 372.6698, 
    260.64, 20.91498, 0.5449734, 0, 0, 0, 0, 0, 0.1160287, 111.142, 209.0083, 
    276.4948, 646.7979, 765.1041, 724.9354, 477.4805, 577.1857, 463.0179, 
    431.689, 425.1302, 450.4791, 382.4208, 78.48548, 0, 0, 0, 0, 0, 
    0.003998051, 0.002220947, 0, 0, 0, 0, 0, 0, 0, 105.1281, 169.7474, 
    236.0875, 9.81155, 0.1445957, 0, 0,
  489.275, 506.2431, 635.707, 891.2947, 1140.819, 104.9125, 0.5735672, 
    0.0001255112, 2.393601, 199.3139, 1536.486, 1511.392, 1079.511, 820.4056, 
    728.9279, 624.3528, 521.0572, 428.4595, 417.1996, 391.4514, 321.5363, 
    234.6511, 206.3434, 187.8103, 161.0246, 103.9707, 3.567678, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 4.888042, 22.56903, 1.230958, 202.7648, 429.525, 
    412.595, 342.0215, 395.2505, 348.6987, 285.1621, 336.5508, 375.4762, 
    287.4457, 307.1478, 204.0902, 144.1289, 12.40784, 0, 0, 0, 0, 0.09297946, 
    48.31137, 410.1348, 219.7555, 321.0481, 912.0163, 957.0075, 782.5162, 
    689.6246, 672.2351, 803.3319, 900.5595, 921.7489, 653.4254, 113.7043, 0, 
    0, 14.97981, 163.9573, 16.21266, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34.01518, 
    399.7357, 415.947, 11.40101, 0, 0, 0,
  423.9285, 419.6786, 540.4236, 810.2414, 880.0971, 25.37736, 0, 0, 43.69834, 
    958.8488, 1720.627, 1412.165, 928.663, 770.8799, 633.066, 510.455, 
    402.9467, 319.4293, 278.5269, 235.3018, 194.7553, 149.0402, 112.7481, 
    124.9141, 133.1899, 112.3536, 20.9965, 2.64545, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2.267793, 70.71137, 122.5515, 31.54795, 87.75684, 313.0298, 326.2078, 
    392.7047, 459.9867, 517.2142, 481.4169, 442.511, 390.7699, 276.8941, 
    289.5733, 344.4179, 305.1668, 167.0574, 9.916601, 1.032431, 1.048887, 
    0.2411555, 23.19702, 397.0361, 721.8358, 320.7461, 332.2949, 979.869, 
    1030.202, 931.765, 809.9, 823.1024, 793.5685, 951.8102, 1033.525, 
    719.0648, 119.1517, 0.833892, 0, 14.80536, 271.7417, 152.8016, 
    0.00275539, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 621.5582, 558.1843, 245.3577, 
    0, 0, 0,
  389.9949, 432.4892, 525.9587, 618.4981, 485.3033, 0.03390811, 0, 1.35604, 
    605.9611, 1549.469, 1794.849, 1175.007, 871.842, 714.1773, 567.928, 
    445.1647, 359.2397, 288.548, 230.5943, 181.9214, 144.2462, 113.5117, 
    92.68795, 83.6313, 99.99515, 113.782, 90.98781, 80.63214, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 10.24857, 59.58021, 91.44401, 35.23301, 92.64501, 269.2377, 
    433.9703, 408.1391, 449.0736, 489.8803, 490.6386, 587.921, 538.6768, 
    542.0423, 504.0613, 493.4232, 387.6947, 149.3013, 21.24825, 2.08333, 
    3.27737, 3.702941, 63.49332, 591.3827, 870.5641, 260.2408, 218.9506, 
    877.173, 980.9655, 1040.86, 1143.761, 991.8488, 921.4819, 835.4803, 
    934.3461, 614.5713, 122.0434, 14.56706, 2.029026, 0, 21.34945, 37.91715, 
    4.003912, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 419.2063, 402.9444, 268.8748, 0, 
    0, 0,
  431.8418, 536.3006, 574.058, 315.8998, 41.75761, 0, 0, 59.75841, 954.189, 
    1557.024, 1298.473, 942.2996, 752.2569, 616.2059, 486.4283, 377.0709, 
    312.1561, 255.6407, 198.0654, 142.262, 116.617, 107.7247, 90.60133, 
    80.00478, 98.95425, 307.284, 343.9886, 272.9455, 6.16348, 0, 0, 0, 0, 0, 
    0, 0, 2.050448, 40.84933, 34.03916, 33.79316, 71.37947, 217.7432, 
    315.7126, 443.3457, 437.9484, 458.0936, 444.2867, 431.0873, 447.9553, 
    504.2306, 471.0587, 559.8055, 493.2112, 392.4747, 196.1293, 47.81644, 
    8.629056, 4.509862, 7.082555, 123.9592, 629.7461, 843.9626, 281.6333, 
    305.7295, 690.8347, 1054.628, 1119.722, 1335.16, 1190.468, 1065.214, 
    984.9171, 869.7607, 546.3845, 225.0289, 150.4363, 163.5934, 3.164987, 
    1.992715, 22.49724, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 167.7594, 192.5879, 
    127.9389, 0, 0, 0,
  464.4328, 710.1633, 619.1936, 47.74748, 0.006608745, 0, 1.039034, 425.7875, 
    1205.512, 1296.795, 937.6955, 818.3823, 688.7088, 615.1889, 470.3323, 
    343.0821, 270.3759, 214.7289, 163.605, 112.6529, 104.0565, 122.8048, 
    107.724, 95.03403, 378.6848, 553.5956, 557.1316, 213.1545, 0, 0, 0, 0, 0, 
    0, 0, 3.253178, 4.987194, 15.42553, 23.11442, 53.14434, 198.1807, 
    390.6396, 476.5912, 416.6757, 370.3962, 423.6606, 388.2758, 315.9665, 
    300.9809, 279.9049, 272.6179, 240.4554, 254.8682, 231.5103, 158.6761, 
    75.81209, 21.71908, 9.130775, 31.90206, 180.6022, 519.5223, 818.9929, 
    367.1069, 232.1573, 540.9075, 1020.897, 1331.289, 1515.057, 1429.161, 
    1326.372, 1300.804, 1167.494, 857.9363, 537.9557, 430.6571, 235.6319, 
    105.8424, 52.64319, 52.60298, 48.16794, 5.177803, 0.0127918, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 7.925615, 7.623189, 0, 0, 0,
  541.9563, 702.7642, 525.0195, 0.008912559, 0, 0.7958623, 220.1246, 
    1012.623, 1381.692, 1054.735, 911.1928, 865.9833, 754.9418, 683.0833, 
    507.5714, 339.2844, 241.6909, 185.5594, 133.8963, 81.90056, 93.08733, 
    116.5835, 104.0461, 220.4304, 362.2358, 272.5128, 22.4466, 0, 0, 0, 0, 0, 
    0.464163, 2.217875, 1.132218, 118.9751, 48.45937, 24.96659, 68.75862, 
    119.5871, 168.0666, 359.0999, 420.4307, 372.978, 292.5229, 326.5298, 
    261.4095, 174.0229, 145.3442, 113.1015, 90.15494, 74.61478, 49.53991, 
    51.27683, 45.57203, 19.36777, 16.3014, 20.58949, 212.4812, 371.5741, 
    567.3152, 837.6189, 773.0519, 254.7844, 402.2862, 1117.507, 1593.182, 
    1713.899, 1657.007, 1585.993, 1660.75, 1626.9, 1297.729, 1008.488, 
    628.0763, 368.5419, 180.6032, 125.0678, 198.4454, 235.6197, 149.7811, 
    32.02615, 2.138504, 0.001609906, 0, 0.0001999206, 0, 0, 0, 0, 0, 
    0.04724865, 3.110864, 0, 0, 0,
  549.2347, 686.2816, 401.375, 0, 0, 65.01826, 822.366, 1329.428, 1219.403, 
    975.2758, 969.5549, 932.9362, 803.3354, 731.2571, 572.4413, 387.7809, 
    255.709, 181.6068, 113.3861, 42.95264, 32.65179, 33.98416, 38.83173, 
    138.7656, 318.7718, 0.7992804, 0, 4.0433, 27.02569, 43.15045, 65.88136, 
    171.93, 328.6717, 326.6402, 310.495, 300.1921, 112.6526, 39.34247, 
    116.7174, 196.2544, 210.7351, 281.5956, 376.5725, 369.3636, 290.0414, 
    245.2731, 172.5113, 134.9192, 115.1656, 85.47749, 72.11951, 66.97635, 
    58.92198, 81.27972, 173.3912, 214.537, 108.2215, 198.1225, 218.5382, 
    378.2805, 263.0815, 752.1837, 870.6851, 687.0273, 413.0518, 1141.952, 
    1943.944, 2054.098, 1926.115, 1828.285, 1968.703, 1788.26, 1402.79, 
    904.152, 675.1245, 442.3218, 270.6985, 164.4036, 201.3591, 233.2095, 
    139.005, 55.39569, 31.88385, 19.8936, 0, 0, 0, 0, 0, 0, 0, 0.36459, 
    2.782869, 0, 0, 0,
  535.8906, 600.8014, 335.9744, 0, 0, 154.2405, 912.732, 1109.16, 989.4586, 
    950.7682, 958.7252, 936.9157, 774.5905, 743.4534, 586.5957, 444.2589, 
    308.8711, 197.4996, 96.48969, 12.3244, 0.1483047, 0.03790293, 0.1436228, 
    37.92851, 155.9851, 30.76747, 221.6138, 252.8131, 416.8718, 624.1976, 
    699.0229, 728.5979, 841.8627, 953.5579, 886.6041, 601.1133, 92.53477, 
    32.85394, 103.7375, 188.0701, 216.8431, 268.9015, 362.442, 393.7513, 
    334.8778, 224.5274, 158.4746, 126.387, 112.2802, 112.7532, 257.5196, 
    397.1968, 538.8138, 1240.1, 2032.906, 2200.138, 2236.536, 1966.697, 
    1706.219, 1459.807, 783.1836, 362.6883, 642.8234, 493.0027, 840.9872, 
    1130.427, 2271.913, 2496.004, 2172.94, 1901.212, 2118.338, 2085.24, 
    1574.87, 1081.068, 810.9539, 635.4389, 423.6662, 250.8699, 288.964, 
    307.7717, 284.6146, 159.4874, 139.9633, 136.567, 123.2743, 19.75318, 0, 
    0, 0, 0, 0, 0, 0.3498602, 0, 0, 0,
  617.859, 478.8044, 162.5502, 0, 0.316467, 273.1028, 967.5567, 1024.078, 
    960.9479, 962.3912, 987.4086, 923.9738, 816.1489, 736.3137, 601.2943, 
    460.8235, 324.0718, 168.9982, 49.51987, 10.05844, 0.003400783, 0, 
    0.6139406, 3.471415, 65.67765, 299.1868, 664.0464, 680.472, 861.0681, 
    1173.805, 1176.411, 882.2818, 935.2615, 1119.443, 1414.621, 875.902, 
    96.9949, 90.53958, 68.45934, 107.9565, 151.2383, 211.1697, 253.7371, 
    301.2069, 273.2981, 195.7737, 154.6178, 177.9713, 194.5825, 716.4048, 
    1805.13, 2597.123, 3127.537, 3920.587, 4658.365, 4768.674, 4483.495, 
    4462.699, 4175.957, 3900.408, 2836.106, 1404.504, 405.8325, 765.2993, 
    1341.417, 1822.338, 2584.409, 2872.491, 2385.164, 1991.338, 2122.929, 
    2156.027, 1849.882, 1308.424, 1070.509, 911.2019, 667.9567, 410.6019, 
    468.2829, 439.6035, 464.8657, 421.4958, 294.738, 311.5735, 259.9264, 
    141.5647, 14.46012, 0, 0, 0, 196.0959, 1.784637, 0, 0, 0, 0,
  589.6921, 369.2813, 29.13641, 0, 10.16494, 462.0075, 953.4734, 992.8953, 
    961.825, 980.4223, 959.9498, 878.5264, 782.0342, 714.8068, 590.7191, 
    438.146, 255.681, 89.16268, 4.204259, 2.031146, 0, 103.8879, 350.6954, 
    283.9107, 257.0193, 369.5965, 704.6323, 645.6995, 1036.557, 1464.105, 
    1060.085, 778.238, 741.6763, 1037.683, 1462.557, 1146.481, 278.6887, 
    344.5007, 247.6657, 85.39928, 122.3622, 162.2269, 193.9326, 217.9708, 
    211.0545, 208.4449, 336.8265, 831.7836, 1583.831, 2516.133, 3871.765, 
    4676.438, 4954.179, 5109.451, 5170.38, 4871.32, 4830.958, 4825.001, 
    4712.904, 4750.763, 4316.47, 2986.506, 1810.279, 1907.389, 3094.098, 
    3158.578, 3400.082, 3428.866, 3037.146, 2417.081, 2381.95, 2137.81, 
    1823.436, 1536.647, 1236.298, 1032.425, 829.5073, 612.1199, 627.1792, 
    549.0421, 514.0405, 437.2412, 523.9689, 332.4905, 376.6574, 324.6547, 
    278.9478, 18.89644, 0.006937383, 11.19048, 622.1964, 266.2146, 0, 0, 0, 0,
  418.7992, 35.6242, 0, 0.003005615, 134.9476, 670.2584, 953.2305, 938.2223, 
    913.4232, 907.8433, 847.9294, 775.7874, 707.1496, 637.6665, 506.9577, 
    328.1991, 144.9271, 21.72296, 0.001061579, 0, 193.2861, 655.1348, 
    890.2563, 1015.931, 1077.46, 1348.436, 1022.688, 766.3108, 1302.777, 
    1343.477, 1030.237, 887.298, 1036.799, 1030.548, 1415.412, 1369.234, 
    954.7562, 897.3719, 604.0056, 161.5459, 117.0032, 160.0316, 186.1864, 
    199.844, 234.4324, 490.8765, 1452.577, 2787.096, 3704.978, 4565.677, 
    5041.605, 5282.9, 5283.827, 5293.211, 5223.339, 5147.862, 5045.44, 
    5014.276, 4810.225, 4833.973, 4828.4, 4279.334, 3368.46, 3630.062, 
    4304.909, 4239.586, 3954.809, 3997.183, 3638.99, 3208.818, 2409.19, 
    1711.776, 1245.757, 1107.457, 1129.331, 956.4644, 789.5651, 568.699, 
    588.8917, 465.5713, 293.4032, 391.9729, 524.9534, 425.9501, 367.7643, 
    501.6449, 504.5149, 232.682, 5.703031, 0.4608422, 517.0116, 853.5552, 0, 
    0, 0, 0,
  208.9919, 0.07399444, 0, 86.20094, 452.0786, 852.0658, 1002.409, 962.3193, 
    888.443, 812.5153, 720.5767, 644.718, 631.5153, 512.2603, 381.4651, 
    213.2256, 41.59562, 0.2816853, 0, 124.2844, 722.3979, 1113.143, 1471.473, 
    1611.769, 2112.062, 2108.031, 1182.046, 772.6594, 1133.844, 1030.302, 
    594.0649, 781.9883, 976.3713, 996.936, 1344.194, 1913.446, 1758.966, 
    1584.213, 828.5089, 218.7474, 120.6228, 168.4115, 186.3442, 204.9695, 
    454.7095, 1957.652, 3490.757, 4445.193, 5092.852, 5200.075, 5270.465, 
    5072.342, 5013.149, 4973.931, 4979.826, 5028.506, 4968.484, 5000.479, 
    4901.846, 4918.038, 5056.896, 4726.156, 4305.746, 4395.774, 4665.846, 
    4441.66, 4191.952, 4342.861, 4170.3, 3571.407, 2256.272, 978.5087, 
    515.0765, 648.3031, 832.2507, 1023.514, 805.8867, 528.6307, 476.446, 
    414.0162, 249.9183, 179.4859, 455.012, 263.6515, 333.0435, 479.9664, 
    632.377, 499.215, 167.3804, 1.14105, 187.7418, 1096.691, 4.065651, 0, 0, 0,
  217.0772, 0.0330215, 14.08818, 507.184, 689.6525, 956.0153, 1135.08, 
    1068.822, 935.9532, 833.0918, 700.9478, 584.4554, 511.998, 405.4882, 
    298.7473, 151.3782, 10.5746, 0, 13.38639, 627.0316, 1415.375, 1796.191, 
    1776.488, 2020.439, 2216.457, 1986.079, 824.9573, 609.1418, 1088.619, 
    704.4744, 531.5552, 655.2637, 836.7814, 991.5665, 1400.434, 1907.079, 
    2138.898, 1730.733, 856.8054, 192.3337, 187.5201, 182.8071, 191.2734, 
    306.0225, 1638.453, 3471.865, 4649.002, 5009.791, 4932.093, 5040.752, 
    4961.458, 4920.357, 4891.655, 4887.036, 4862.397, 4830.989, 4769.84, 
    4764.334, 4749.213, 4840.669, 4871.838, 4824.714, 4635.75, 4551.147, 
    4447.096, 4367.069, 4249.624, 4367.218, 4152.088, 3556.254, 2167.627, 
    517.2781, 330.44, 333.8921, 615.7012, 814.1959, 880.6069, 573.7075, 
    426.0545, 368.3916, 209.4412, 130.0882, 280.0025, 206.5527, 246.2915, 
    389.107, 555.9575, 505.8926, 402.7588, 39.14849, 0.2409696, 211.2308, 
    10.10999, 0.2490215, 8.65174, 0.6303881,
  32.38083, 0, 51.82127, 560.3418, 760.4517, 1012.509, 1175.754, 1092.682, 
    990.1829, 844.8569, 664.1961, 527.9617, 436.3003, 353.342, 264.007, 
    111.6445, 0.1420982, 0, 120.9445, 1149.31, 1999.209, 1945.943, 1973.386, 
    1762.449, 1950.817, 1315.04, 577.0366, 879.3376, 1191.386, 623.9373, 
    548.0479, 722.4045, 1082.094, 1262.284, 1544.662, 2178.558, 2164.37, 
    1978.036, 1035.92, 460.3963, 275.0108, 282.9265, 595.8168, 1425.515, 
    3292.09, 4695.376, 5096.314, 4968.224, 4930.162, 4852.206, 4795.105, 
    4827.783, 4907.193, 5035.4, 4982.63, 5017.723, 4947.738, 4862.034, 
    4921.563, 4884.641, 4879.072, 4878.018, 4793.002, 4559.51, 4386.215, 
    4295.125, 4247.954, 4282.634, 4102.235, 3924.184, 2823.693, 1224.186, 
    358.0084, 332.7956, 348.9137, 678.3985, 848.0242, 821.4729, 618.2599, 
    296.2792, 78.22495, 69.06935, 236.8286, 218.569, 131.588, 226.8546, 
    405.3286, 521.6719, 575.6138, 185.445, 0.1386309, 0, 0.01035178, 0, 0, 
    0.3566946,
  0, 3.552063, 321.7133, 849.3109, 976.9869, 1078, 1041.034, 971.9257, 
    896.7177, 738.8071, 609.843, 479.6385, 370.4907, 299.6009, 196.0335, 
    43.93956, 1.847782, 58.31754, 820.1542, 1913.927, 2158.314, 2047.404, 
    1703.193, 1653.195, 1413.601, 1037.866, 736.9638, 1415.212, 1414.237, 
    810.8496, 802.1318, 1344.746, 1755.177, 1950.15, 2215.817, 2564.552, 
    2719.364, 2259.201, 1462.947, 672.4842, 476.5094, 949.2522, 1674.35, 
    3053.793, 4114.063, 4946.655, 5076.482, 5097.934, 5060.518, 5084.558, 
    5115.013, 5053.414, 5074.056, 5093.611, 5064.592, 5146.818, 5095.178, 
    5143.528, 5132.971, 5072.526, 4904.224, 4783.976, 4806.5, 4586.318, 
    4403.593, 4429.247, 4359.3, 4282.01, 4076.977, 3919.891, 3721.054, 
    2170.56, 812.0792, 348.9857, 379.0044, 509.2384, 835.6813, 1042.576, 
    981.3938, 473.188, 59.4187, 54.51209, 257.2173, 304.478, 147.0937, 
    83.89629, 318.8223, 480.2112, 706.43, 507.7156, 43.1609, 0, 0, 0, 
    0.06568222, 0,
  0, 74.23603, 787.8488, 1047.875, 1021.896, 987.5112, 943.1434, 865.201, 
    751.0483, 636.3491, 527.4158, 403.2906, 282.5342, 179.8925, 87.43723, 
    3.748239, 13.04159, 420.638, 1624.73, 2216.099, 2128.865, 1733.536, 
    1583.128, 1268.357, 1247.077, 910.689, 1149.7, 1639.568, 1381.821, 
    977.155, 1235.957, 1915.405, 2513.842, 2519.291, 2726.454, 3145.376, 
    2913.469, 2521.798, 1770.634, 1137.481, 1062.631, 1737.886, 2865.038, 
    3579.866, 4525.335, 4868.795, 5310.432, 5363.74, 5347.537, 5387.418, 
    5274.167, 5170.409, 5133.905, 5203.841, 5101.455, 5070.62, 5106.412, 
    5089.334, 5089.588, 4879.959, 4693.276, 4713.932, 4758.439, 4678.091, 
    4520.184, 4536.472, 4453.167, 4362.481, 4144.474, 3822.403, 3798.529, 
    3049.53, 1477.426, 703.8835, 612.568, 658.7606, 819.6526, 1062.141, 
    1055.71, 575.3791, 73.42055, 27.57079, 103.5562, 207.4734, 120.4412, 
    30.39635, 148.8998, 383.1422, 591.7628, 532.1869, 174.8339, 1.234607, 0, 
    0, 0, 0,
  6.758009, 487.5991, 1021.831, 1115.679, 886.489, 892.4991, 847.3696, 
    758.7397, 623.5787, 508.0063, 426.4549, 305.7114, 158.1539, 48.50787, 
    5.502139, 5.127207, 40.45427, 1082.158, 2018.84, 2095.057, 1691.412, 
    1381.58, 1191.657, 1015.282, 1019.028, 1079.314, 1296.271, 1340.825, 
    1178.45, 832.3215, 1319.656, 1844.028, 2394.739, 2776.184, 3035.285, 
    3199.43, 3069.708, 2704.726, 3048.322, 2788.972, 2680.07, 3130.915, 
    3342.005, 4203.668, 4655.496, 5272.828, 5415.704, 5200.595, 5129.409, 
    5031.954, 5205.507, 5085.389, 5081.525, 5094.905, 5042.618, 5019.026, 
    4992.753, 5047.111, 5006.662, 4865.849, 4714.873, 4635.37, 4685.44, 
    4620.996, 4597.202, 4502.657, 4462.631, 4332.861, 4098.364, 3766.416, 
    3657.072, 3297.008, 2097.184, 1253.378, 1089.461, 1061.64, 1174.932, 
    1281.606, 1266.194, 835.1642, 263.9403, 79.5519, 32.27344, 68.0872, 
    131.0868, 118.724, 164.2968, 321.6274, 409.3891, 379.2769, 350.8774, 
    57.88399, 0.000805264, 0, 0, 0,
  238.1623, 791.4998, 1109.681, 899.7229, 803.0744, 786.03, 737.5471, 
    634.7917, 498.6732, 393.5605, 324.9799, 180.8011, 45.09904, 5.052932, 
    12.10084, 59.62862, 665.7957, 1742.159, 2304.37, 1936.526, 1518.453, 
    1209.02, 957.4006, 869.3815, 823.4235, 999.6229, 1120.257, 1287.387, 
    1058.116, 943.8759, 842.4662, 1182.286, 1637.921, 2097.368, 2345.563, 
    2374.775, 1990.883, 2252.895, 3334.049, 3940.562, 4061.273, 4010.166, 
    4178.608, 4529.894, 4820.277, 4816.019, 4359.409, 3582.755, 3025.995, 
    3098.254, 3615.333, 4245.46, 4695.494, 5053.856, 5057.838, 5040.737, 
    4995.706, 4951.887, 5012.489, 4828.667, 4652.396, 4480.73, 4422.274, 
    4482.873, 4418.603, 4365.641, 4435.617, 4158.283, 3927.431, 3744.359, 
    3460.329, 3134.216, 2236.319, 1473.672, 1232.209, 1085.229, 938.4994, 
    930.7794, 780.1253, 518.0501, 171.889, 131.0825, 128.4954, 145.3723, 
    306.1799, 273.0995, 216.7841, 302.7602, 352.1556, 292.1012, 300.0482, 
    151.9467, 1.769033, 0, 0, 0,
  762.3385, 958.6488, 967.5426, 836.1221, 672.2523, 743.9036, 705.8074, 
    585.7993, 412.0986, 315.1353, 220.0953, 76.00178, 7.931051, 19.07306, 
    352.5095, 807.7217, 1467.913, 2206.177, 2116.3, 1479.32, 1129.964, 
    788.2949, 807.8799, 715.9404, 766.021, 992.697, 1301.655, 1434.707, 
    1353.936, 786.4489, 618.7448, 572.2695, 753.1136, 781.6061, 869.8459, 
    807.5753, 789.2447, 793.95, 2282.462, 3481.706, 4177.188, 4562.651, 
    4439.226, 4581.507, 3711.448, 2810.206, 2234.735, 1677.431, 1388.387, 
    1278.489, 1672.559, 2128.335, 3001.532, 3830.48, 4550.405, 4801.908, 
    4633.007, 4499.204, 4535.861, 4201.199, 3729.332, 3460.189, 3439.621, 
    3560.627, 3621.553, 3831.16, 4091.066, 3848.02, 3584.761, 3534.397, 
    3254.213, 2773.562, 2217.112, 1683.945, 1579.851, 1373.786, 1237.948, 
    1035.855, 892.402, 538.7142, 249.4172, 148.4552, 154.6931, 130.894, 
    219.8244, 191.3214, 59.69934, 129.1412, 212.872, 166.6351, 130.7894, 
    118.5202, 14.56528, 0, 0, 0,
  989.5663, 927.1322, 930.0528, 724.9628, 672.3023, 786.1067, 760.7014, 
    580.4506, 387.8854, 255.2157, 132.3959, 20.43845, 25.85789, 478.4587, 
    1034.186, 1562.984, 1919.749, 2048.771, 1455.002, 993.2492, 1055.018, 
    1015.837, 1037.239, 1008.556, 891.994, 1129.969, 1403.661, 1486.652, 
    921.8677, 453.2355, 336.5799, 424.1663, 397.4917, 279.882, 307.3911, 
    629.627, 392.5599, 732.6076, 1854.792, 3292.929, 4316.049, 4438.208, 
    4466.581, 3936.618, 2551.772, 1529.796, 1225.804, 1185.416, 1170.846, 
    1186.658, 1149.756, 1173.267, 1364.58, 2012.139, 2864.934, 3708.189, 
    4220.437, 4108.575, 3883.59, 3378.89, 2934.686, 2709.543, 2824.293, 
    3108.43, 3076.333, 3295.794, 3656.051, 3385.662, 3217.673, 3000.589, 
    2639.363, 2225.868, 2004.855, 1872.814, 1614.911, 1220.716, 921.0709, 
    856.4285, 921.3516, 950.4296, 616.0353, 308.2891, 110.1128, 48.46398, 
    55.95203, 45.66961, 26.53019, 25.74332, 58.75687, 44.34055, 7.046542, 
    9.698866, 7.823508, 0.1154567, 0, 0,
  873.5029, 932.446, 802.8636, 679.261, 728.6178, 853.7338, 757.9206, 
    581.5193, 393.3805, 206.899, 67.25694, 23.86274, 177.6185, 981.5392, 
    1598.842, 1796.156, 1947.744, 1703.935, 1375.229, 1515.294, 1642.378, 
    1676.018, 1487.45, 1227.913, 1159.733, 1323.913, 1554.071, 1138.957, 
    556.8956, 169.3183, 218.1516, 265.9337, 235.5797, 302.2885, 690.3524, 
    1159.933, 1460.098, 1501.492, 2359.936, 3452.56, 4296.354, 4520.364, 
    4153.528, 3140.282, 1694.784, 1188.321, 1116.658, 1141.684, 1149.989, 
    1137.289, 1126.685, 1111.867, 1065.968, 976.756, 1235.389, 1905.175, 
    2724.575, 3200.128, 3303.74, 2937.104, 2721.535, 2951.062, 3359.012, 
    3876.756, 3978.864, 3924.08, 3884.962, 3585.292, 3361.129, 3095.249, 
    2504.762, 2074.735, 1898.636, 1876.1, 1742.129, 1328.015, 1136.963, 
    851.3479, 765.448, 628.5696, 611.1027, 228.0393, 106.5588, 40.51612, 
    28.73609, 26.4498, 39.7077, 42.63209, 21.35075, 11.05065, 3.122396, 
    2.336835, 0.5792097, 0.1638553, 0, 0,
  546.0862, 803.7518, 720.4936, 680.9647, 811.3162, 854.0582, 728.9124, 
    554.4362, 350.1646, 161.0941, 51.3675, 48.73245, 369.3617, 1295.04, 
    1821.616, 1891.482, 1897.59, 1783.333, 1780.204, 1693.617, 841.7841, 
    444.8978, 635.6622, 896.0977, 1128.595, 1378.011, 996.2464, 523.0845, 
    123.556, 142.2115, 182.9801, 192.1028, 208.9994, 239.5104, 673.2095, 
    1674.933, 2271.34, 2666.304, 2851.325, 3098.809, 3555.89, 3740.312, 
    3572.558, 2706.249, 1709.02, 1359.368, 1286.218, 1109.896, 1039.783, 
    1053.64, 1038.432, 1022.949, 1007.573, 974.9078, 853.291, 834.8326, 
    1136.756, 1648.817, 2111.175, 2467.282, 2775.722, 3019.613, 3544.646, 
    4111.462, 4240.049, 4245.177, 4150.613, 3692.481, 3492.051, 3113.697, 
    2519.094, 1983.502, 1739.186, 1723.87, 1627.539, 1467.329, 1415.479, 
    1188.471, 862.6572, 819.2594, 613.4723, 440.3748, 103.548, 44.31029, 
    44.08937, 32.32762, 27.8348, 27.06621, 14.8008, 2.686884, 3.042891, 
    2.475014, 0.1258945, 0, 0, 0,
  287.7358, 699.6454, 753.7252, 715.9815, 790.1022, 770.7126, 621.1946, 
    429.5545, 302.6275, 146.0066, 109.7574, 238.4723, 702.8896, 1500.438, 
    1914.869, 1864.13, 1797.373, 1384.315, 1103.181, 50.18019, -29, 
    -28.77262, 25.38564, 296.886, 687.7216, 647.961, 349.3248, 83.32568, 
    112.7014, 157.216, 171.5177, 178.561, 204.0525, 312.3961, 523.767, 
    829.8365, 1039.718, 1047.279, 1355.524, 1172.16, 1411.563, 2336.885, 
    3058.305, 3226.443, 3063.086, 2861.304, 2247.198, 1404.461, 1073.007, 
    987.9013, 956.4599, 926.052, 903.3677, 896.808, 893.4102, 892.0126, 
    796.2086, 820.1337, 984.0677, 1229.673, 1469.496, 1966.5, 2469.902, 
    3181.495, 3622.321, 3652.744, 3231.653, 2652.689, 2285.655, 2040.421, 
    1670.866, 1479.306, 1414.353, 1424.594, 1447.813, 1503.411, 1473.374, 
    1250.532, 1041.187, 973.3618, 1039.013, 789.7152, 424.5931, 71.7645, 
    43.34607, 37.34945, 45.60085, 23.38318, 6.514248, 1.005424, 1.192295, 
    0.07372784, 0, 0, 0, 0,
  280.0255, 717.2288, 800.9051, 767.515, 678.3198, 625.6271, 422.783, 
    283.5512, 241.4006, 186.5598, 174.9805, 521.5108, 1183.758, 1658.958, 
    2034.699, 1761.583, 1296.187, 204.5876, -27.33, -29, -29, -28.70372, 
    31.97342, 167.3994, 247.8943, 170.875, 60.56211, 102.6041, 146.6671, 
    170.812, 176.8664, 183.8537, 244.3707, 366.5971, 502.9418, 470.5995, 
    290.3222, 581.1486, 1270.705, 1402.007, 1254.245, 1784.784, 2600.036, 
    2944.01, 3219.255, 3399.147, 3218.488, 2378.177, 1818.334, 1375.318, 
    1074.772, 1071.595, 984.6507, 961.2864, 971.7458, 1197.327, 1193.799, 
    1028.109, 963.4049, 965.5383, 1135.214, 1159.892, 1419.062, 1704.113, 
    1884.114, 1810.738, 1669.92, 1423.683, 1450.932, 1501.812, 1357.503, 
    1354.311, 1357.144, 1350.14, 1337.69, 1373.946, 1390.578, 1208.278, 
    1047.752, 1206.215, 1150.309, 1096.129, 627.1903, 92.17794, 38.86603, 
    55.03728, 97.46461, 80.68608, 19.16875, 1.530113, 0.02449018, 0, 0, 0, 0, 0,
  278.7002, 848.4108, 836.0483, 703.4719, 592.2507, 425.2289, 267.3521, 
    212.9088, 260.6262, 199.7883, 384.8431, 1051.43, 1458.136, 1718.665, 
    1860.108, 1682.248, 920.7298, -29, -29, -29, -29, -26.10924, 98.29451, 
    120.4517, 76.57224, 60.59356, 87.99368, 121.3795, 137.9679, 144.398, 
    164.9114, 216.217, 274.5612, 275.6122, 318.0442, 259.2065, 230.8655, 
    623.9655, 1918.901, 2278.465, 2228.787, 2412.379, 2568.84, 2575.392, 
    2590.898, 2936.103, 3116.961, 3308.007, 3364.986, 2819.327, 2346.359, 
    2102.324, 1968.311, 1727.268, 1581.183, 1342.206, 1030.278, 1016.645, 
    1021.907, 1084.763, 1044.676, 1257.469, 1468.743, 1774.683, 1740.715, 
    1517.49, 1302.269, 1243.797, 1198.531, 1266.439, 1397.631, 1400.947, 
    1359.057, 1343.482, 1246.818, 1367.203, 1329.797, 1222.678, 1103.928, 
    1230.625, 1299.724, 1154.313, 827.8479, 142.0308, 30.594, 63.95813, 
    176.8368, 209.5096, 94.29587, 2.645784, 0, 0, 0, 0, 0, 0,
  372.7461, 1182.848, 984.7722, 758.8289, 559.1176, 423.6849, 319.4374, 
    300.4261, 340.6555, 502.4338, 1127.504, 1562.021, 1634.167, 1688.647, 
    1848.811, 1538.005, 454.8116, -28.99981, -29, -29, -27.34004, 37.3294, 
    157.3012, 172.0072, 120.2076, 77.74836, 81.51273, 100.2689, 110.1352, 
    113.6465, 112.3892, 174.2308, 265.0841, 238.038, 208.7626, 195.9964, 
    185.5608, 428.3402, 1028.99, 1427.11, 1409.885, 1349.094, 1442.432, 
    1663.696, 1924.178, 2039.838, 2233.458, 2097.392, 2286.286, 2274.246, 
    2335.328, 2740.635, 3043.788, 3113.309, 2620.314, 1823.444, 907.4882, 
    560.1979, 721.8196, 618.8461, 714.8278, 968.9215, 1536.432, 1776.954, 
    1845.922, 1518.606, 1331.444, 1091.121, 1037.558, 1111.581, 1316.298, 
    1388.658, 1346.563, 1293.286, 1239.811, 1305.997, 1406.889, 1326.371, 
    1211.889, 1292.238, 1407.659, 1205.926, 807.7815, 109.0812, 17.7631, 
    51.74597, 188.0972, 276.9687, 185.2122, 45.17762, 0, 0, 0, 0, 0, 0,
  23.64984, 599.7591, 511.6504, 444.8416, 378.2097, 360.2961, 380.9373, 
    438.2814, 595.3414, 1348.148, 2057.229, 2197.964, 1472.968, 1671.91, 
    1237.43, 761.7867, 28.29826, -28.70648, -28.99438, -29, -24.99033, 
    18.25178, 63.3651, 174.8866, 123.8744, 57.97906, 65.55949, 76.69518, 
    97.68421, 102.3149, 131.3378, 195.444, 256.4067, 243.5822, 187.5729, 
    165.1665, 342.9257, 405.3759, 560.9412, 516.8105, 509.3314, 621.6459, 
    699.2636, 746.7856, 760.3452, 922.6527, 823.6852, 1078.508, 1096.203, 
    1233.275, 1588.237, 2370.672, 2694.676, 2629.588, 2156.679, 1783.274, 
    1690.359, 1606.746, 1283.696, 1141.156, 1217.001, 1620.093, 1467.414, 
    1503.383, 1485.695, 1331.391, 1196.225, 1032.619, 951.8022, 972.683, 
    1066.139, 1124.131, 1171.412, 1188.777, 1279.054, 1209.068, 1229.401, 
    1345.554, 1244.472, 1249.917, 1464.447, 1206.628, 878.3694, 171.7012, 
    12.43563, 7.429965, 32.89956, 78.383, 51.98663, 29.90217, 24.32074, 0, 0, 
    0, 0, 0,
  1.67216, 340.6524, 385.0545, 416.1772, 390.3365, 441.3774, 650.9087, 
    704.9575, 1160.624, 1782.02, 2326.5, 2033.687, 1439.484, 1619.828, 
    746.22, 75.66013, 201.0358, 17.39066, -28.43431, -29, -27.93392, 
    -29.96976, 155.6212, 198.6232, 113.8873, 86.04948, 76.57941, 72.31518, 
    72.27863, 74.17043, 85.37265, 140.0728, 171.7061, 157.3423, 148.0897, 
    287.3974, 366.4878, 442.8387, 367.5465, 295.4169, 339.7092, 412.319, 
    477.4836, 479.2714, 430.4697, 594.4115, 1253.493, 1810.096, 2104.204, 
    1634.684, 1001.775, 974.5079, 900.9539, 634.2441, 554.7181, 615.168, 
    911.0193, 996.5089, 1222.358, 1436.428, 1665.35, 1462.017, 1208.923, 
    960.894, 1190.559, 1318.656, 1208.269, 1155.516, 1205.878, 1180.793, 
    1165.779, 1183.944, 1099.437, 1158.785, 1276.583, 1278.646, 1152.482, 
    1210.833, 1241.654, 1143.037, 1397.42, 1334.603, 1178.972, 665.2888, 
    53.88091, 2.508959, 0.1916037, 1.167866, 4.74597, 36.34115, 73.30758, 
    20.18326, 0, 0, 0, 0.04834903 ;

 land_mask =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01177494, 
    0.2004458, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01095872, 0, 0.003575196, 0, 
    0.04133711, 0.4170527, 0.86152, 0.830821, 0.6877613,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1264342, 0.5097121, 0.8753754, 
    0.7817355, 0.2817629, 0.5366528, 0.9293424, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1668709, 0.9869201, 1, 1, 1, 
    0.9988317, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.06910358, 0.8185359, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.08511406, 0.7756319, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.5162452, 0.9977401, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.3129568, 0.9959389, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.02861756, 0.6951866, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1453591, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1453354, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.6664422, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0.02644386, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.175007, 0.9126859, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1,
  0.6233622, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2911646, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1,
  0.6379205, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.7788954, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1,
  0.6378774, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.005386431, 0.309769, 0.4789902, 
    0.1082563, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.7179049, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0.6374285, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01172521, 1, 1, 0.7862632, 
    0.2317922, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.6998634, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0.06200648, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2357621, 1, 1, 1, 0.9253088, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.8606739, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.5966171, 1, 1, 1, 0.9915225, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.519107, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1,
  0.3754489, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.5966566, 1, 1, 1, 0.9932248, 
    0.07400899, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.2909555, 1, 0.9996659, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0.9468521, 0.2389454, 0, 0, 0, 0, 0, 0, 0, 0, 0.1795021, 1, 1, 1, 1, 
    0.5510066, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1121078, 
    0.2244427, 0.2677908, 0.8841233, 0.9811913, 0.7802478, 0.9785666, 
    0.8345276, 0.9690673, 0.8673143, 1, 1, 1, 1,
  1, 0.9377849, 0.1510155, 0, 0, 0, 0, 0, 0, 0, 0.004869109, 0.7091162, 1, 1, 
    1, 0.7690508, 0.04686088, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.08630638, 0.05072459, 0.00715183, 0.05010708, 0.0435742, 
    0.04084156, 0.4005074, 1, 1, 1, 1,
  1, 1, 0.5535783, 0, 0, 0, 0, 0, 0, 0, 0.0003298247, 0.4347998, 1, 1, 1, 1, 
    0.1105905, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.1101263, 0.8236522, 1, 1, 1,
  1, 1, 0.9985871, 0.7174072, 0.04896508, 0, 0, 0, 0, 0, 0.0117381, 
    0.9759874, 1, 1, 1, 1, 0.5814301, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.5950869, 0.9525636, 
    0.9839157, 1,
  1, 1, 1, 1, 0.9804606, 0.1933275, 0, 0, 0, 0, 0.01173972, 1, 1, 1, 1, 1, 
    0.6657338, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.0211766, 0.02256984, 0.21058, 0.6582654,
  1, 1, 1, 1, 1, 0.8694932, 0.1387404, 0, 0, 0, 0.01174129, 1, 1, 1, 1, 1, 
    0.9328697, 0.1643069, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.3509133,
  1, 1, 1, 1, 1, 1, 0.8173901, 0, 0, 0, 4.984859e-05, 0.3204487, 0.9584024, 
    1, 1, 1, 1, 0.3567966, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 0.8408963, 0, 0, 0, 0, 0, 0.2506884, 0.7998602, 1, 1, 1, 
    0.7708181, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 0.8408804, 0, 0, 0, 0, 0, 0, 0.002590244, 0.3868952, 1, 
    1, 0.9516376, 0.2383268, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 0.8408653, 0, 0, 0, 0, 0, 0, 0, 0.00495693, 0.7948567, 1, 
    0.7986782, 0.05182758, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 0.8408509, 0, 0, 0, 0, 0, 0, 0, 0, 0.2693094, 0.9602194, 
    0.7707613, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 0.8408375, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.6405759, 
    0.6084861, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 0.8408248, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01842676, 
    0.01816703, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.004960603, 0, 0, 0, 0.4832949, 0.5081044,
  1, 1, 1, 1, 1, 0.822592, 0.252383, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1190309, 
    0.4765593, 0.5912097, 0, 0, 0, 0.1877966, 0.5820142,
  1, 1, 1, 1, 1, 0.6266645, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.07368479, 0, 
    0.06970806, 0.1497295, 0.2323898, 0.3694812, 0.09263787, 0.1388984, 
    0.02827013, 0,
  1, 1, 1, 1, 1, 0.6266469, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01073292, 0.03063297, 0.5991629, 
    0.6986423, 0.8001084, 0.4512461, 0.2554947, 0.185261, 0.05334708, 0, 
    0.08976555, 0.01147698, 0,
  1, 1, 1, 1, 1, 0.6266309, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.04137734, 0.2410906, 0.3296587, 0.6321196, 
    0.8407705, 0.5324757, 0.1355897, 0.1754358, 0.02694144, 0.0008469501, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 0.3423578, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.005920551, 0.2284444, 0.6276525, 0.7197345, 0.8359697, 1, 
    1, 0.8431623, 0.505213, 0.04540349, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 0.01733314, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.284229, 0.6896634, 1, 0.8693293, 0.349668, 0.3810897, 
    0.6086794, 0.240112, 0.01585283, 0.1599976, 0, 0, 0, 0, 0, 0, 0, 
    1.805722e-05, 0, 0.03666643, 0.119504, 0, 0,
  1, 1, 1, 1, 1, 0.03475345, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.1117143, 0.4876121, 0.4447544, 0.2373162, 0.01928726, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.7862673, 0.3681437, 0.1774964, 0.787069, 
    0.4654977, 0, 0,
  1, 1, 1, 1, 1, 0.6265825, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.3158722, 0.9526677, 0.9008846, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.8407551, 0.3746317, 0.4537332, 0.9686775, 0.3652169, 0, 0,
  1, 1, 1, 1, 1, 0.8866345, 0.1598364, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.03936394, 0.6387691, 0.9943234, 1, 0.9008874, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.01252412, 0.4860564, 0.5318119, 0.2620075, 0, 0, 0.1320914, 
    0.8908585, 0.3907566, 1, 0.8389638, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 0.4656247, 0.0110646, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.6010675, 1, 1, 1, 0.9167563, 0.07269689, 0.2391122, 0.2968679, 0, 
    0.2234619, 0.3493941, 0.8015904, 0.8455765, 0.9577049, 1, 1, 0.4179517, 
    0, 0, 0.4412683, 1, 0.6472766, 1, 0.3203639, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 0.6503397, 0.01531898, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.2558588, 0.9597831, 1, 1, 0.972702, 0.9489372, 0.4348444, 0.1722408, 
    0.04735889, 0, 0.7706258, 1, 1, 1, 1, 1, 1, 0.5972056, 0, 0, 0.1294438, 
    0.8859251, 1, 0.8678412, 0.2493258, 0.1075096, 0.1135316, 0.3466776,
  1, 1, 1, 1, 1, 1, 1, 1, 0.287686, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1325035, 0, 
    0.8317441, 1, 1, 0.9539555, 0.2448101, 0.2613218, 0, 0, 0.1152575, 
    0.2170084, 0.900425, 1, 1, 1, 1, 1, 1, 0.8761324, 0.1775864, 0, 0, 
    0.8103314, 0.4596019, 0.6510904, 0.7820377, 0.592761, 0.06109875, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 0.920251, 0.1775966, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.3923621, 0.987651, 1, 1, 0.3509198, 0.2281306, 0, 0, 0, 0, 0.7061847, 
    1, 1, 1, 1, 1, 1, 1, 1, 0.7719379, 0, 0, 0.6054041, 0, 0, 0.02613228, 
    0.1559717, 0.01388168, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 0.7677791, 0.09293438, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.1779837, 0.3241267, 0.9822798, 1, 1, 0.9843383, 0.2598756, 0.01625016, 
    0, 0, 0, 0, 0.866449, 1, 1, 1, 1, 1, 1, 1, 1, 0.8224034, 0.07974907, 0, 
    0.2945428, 0.6333175, 0.5063159, 0.446091, 0.3369552, 0.4868954, 0.174956,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9503866, 0.2001637, 0.005799863, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.1038464, 0.6664168, 1, 1, 0.8380957, 0.2760953, 0.4406356, 
    0.1536544, 0, 0, 0, 0, 0.8664498, 0.9701261, 0.9560779, 1, 1, 1, 1, 1, 1, 
    1, 0.9252388, 0.3537527, 0.03041064, 0.3419223, 0.4810721, 0.4459109, 
    0.1816519, 0.1972405, 0.5183649,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.6181571, 0.04856747, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.6580371, 1, 0.8227324, 0.4224875, 0.510656, 0.9363688, 0.6996492, 0, 0, 
    0, 0, 0, 0.1081687, 0.109901, 0.5228179, 1, 1, 1, 1, 1, 1, 1, 0.3901491, 
    0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8356921, 0.1330075, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.005403113, 
    0.4351665, 0.9745526, 0.7136913, 0.2152697, 0.3135631, 0.9907392, 1, 
    0.2640299, 0, 0, 0, 0, 0, 0, 0, 0.03659684, 0.3494267, 0.8000365, 
    0.9991509, 1, 1, 1, 0.8337656, 0.1029233, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8476309, 0.1004762, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002844633, 
    0.6518675, 1, 0.7256781, 0.03523427, 0, 0.6580248, 1, 1, 0.2640252, 0, 0, 
    0, 0, 0.3051819, 0, 0, 0, 0, 0, 0.8034117, 1, 1, 1, 0.9529892, 0.2843654, 
    0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.7001464, 0.03844476, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.1336879, 0.05886054, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.2070477, 0.4348271, 0.2998562, 0.06389595, 0, 0.1970171, 0.9302663, 1, 
    0.8744631, 0.138245, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1508173, 0.772752, 
    0.9572471, 1, 1, 0.8470377, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.3652858, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 0.7193018, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.5087034, 0.9593135, 0.7576354, 0.1099733, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.318427, 0.9950952, 1, 0.9854341, 0.3656026, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.7283692, 0.04570163, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.06553631, 0.005726846, 0, 1, 0.448386, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.2178526, 0.8641504, 0.4405744, 0.03868152, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.7589623, 0.9413608, 0.3499206, 
    0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.5236878, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.2793671, 0.9727733, 0.3410493, 0.004538658, 0.9128425, 0.1045216, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2580416, 0.9425887, 0.64642, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1441312, 0.3183418, 0, 
    0, 0, 0, 0.1504084, 0.08207643, 0, 0.1264589, 0.6360483,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8886915, 0.171717, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.4181546, 1, 1, 0.2572959, 0.09995186, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.2655529, 0.9644211, 0.5325517, 0, 0, 0, 0, 0.09022734, 
    0.2022693, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.5111119, 0.0366355, 0.2737309, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.7781987, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0143113, 
    0.8599525, 1, 1, 0.8562455, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.1380162, 0.923599, 0.1353773, 0, 0, 0, 0.03968213, 0.2221394, 
    0.7275295, 0.3227897, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1441023, 
    0.2176893, 0, 0, 0, 0, 0.1160006, 0.885816, 0.6751633, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8664993, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.4873159, 
    1, 1, 1, 0.68866, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.1955505, 0.939324, 0.3395239, 0, 0, 0.1328799, 0.7831334, 1, 1, 
    0.7539828, 0.4905147, 0.03082606, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.04012534, 
    0.5083878, 0, 0, 0, 0, 0, 0.1388984, 0.256223, 0.6417912,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9953002, 0.5326272, 0.519923, 0.4552467, 
    0.5700993, 0.8583444, 0.7375726, 0.923451, 0.9061459, 0.1658801, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1702366, 
    0.9217622, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1872573, 0, 
    0, 0, 0, 0.3864902, 1, 0.6463704, 0, 0.1308702, 0.7559305, 1, 1, 1, 1, 1, 
    0.8225404, 0.1237965, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.084927, 0.5631165, 
    0.1094015, 0, 0, 0.08819825, 0.6943044, 0.07551906, 0.006831904,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.4421961, 0, 0, 0, 0, 0, 0, 0.01769246, 
    0.1738239, 0, 0, 0.1787293, 0.04062913, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.3148586, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0808153, 0.9058402, 0.6547354, 0.2428028, 
    0.7843866, 1, 1, 1, 1, 1, 1, 1, 0.6807549, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.2588764, 0.1009072, 0, 0, 0.2429036, 0.7849156, 0.4656103, 0.169591,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9108992, 0.188346, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.7856974, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.3914096, 1, 1, 0.9854771, 1, 1, 1, 1, 1, 1, 1, 1, 0.6807355, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.7825689, 0.6956174, 0.09677283, 
    0.1274765,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 0.7852127, 0.4266168, 0.8433919, 0.4879982, 
    0.2553098, 0.4059382, 0.1131723, 0.02167348, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2218162, 0.963348, 1, 1, 
    1, 1, 1, 0.688597, 0.09377675, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.01462167, 0.002184577, 0, 0, 0.8908938, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 0.3777061, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.003051978, 
    0.07014503, 0.1355046, 0.1359438, 0.006367458, 0.6373758,
  1, 1, 1, 1, 1, 1, 1, 1, 0.8328858, 0.2307329, 0.8818867, 1, 1, 1, 1, 1, 
    0.691934, 0.4109589, 0.2119478, 0.1284744, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.5544662, 1, 1, 1, 1, 1, 1, 1, 
    0.946013, 0.1113746, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.3114816, 0.7581814, 
    0.5352249, 0.1977297, 0.9311432, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.1334493, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.181796, 0.5997484, 0, 0, 
    0.3158956, 0.500448,
  1, 1, 1, 1, 1, 1, 1, 1, 0.1062542, 0.1823296, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.9209124, 0.0554863, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.7544572, 1, 1, 1, 1, 1, 1, 1, 1, 0.9121619, 0.5140178, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.8938125, 1, 0.7836286, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 0.9445137, 0.6255063, 0.02327494, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.316875, 0.3196791, 0.2422916, 0.0662774, 0.6194771, 0,
  1, 1, 1, 1, 1, 1, 0.8702384, 0.2501028, 0.005983606, 0.5771939, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 0.8631834, 0.8403694, 0.5729032, 0.2040605, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.00724657, 0.7643476, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0.9984289, 0.3873025, 0, 0, 0, 0, 0, 0, 0, 0, 0.2322503, 
    0.9433986, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9763494, 0.1368165, 
    0.0004370618, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1078297, 0.7730162, 
    1, 0.6829644, 0.4463389, 0.2076392, 0.1887735,
  1, 1, 1, 1, 1, 0.8587388, 0.1308349, 0, 0, 0.4788192, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 0.9391835, 0.775203, 0.1979599, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.239585, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9413478, 
    0.3537645, 0.05398361, 0, 0, 0, 0, 0, 0, 0.8853288, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0.9915676, 0.4714071, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.2355691, 1, 0.7928132, 0.1206847, 0, 0, 0,
  1, 1, 1, 1, 1, 0.4860172, 0, 0, 0, 0.7716876, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0.9360449, 0.2212868, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.1080709, 0.2082748, 0.2002707, 0.8915246, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 0.6313275, 0, 0, 0, 0, 0.0001691831, 0.5004879, 0.9755507, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 0.6524076, 0, 0, 0.2558733, 0.5018113, 0.2678142, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.136077, 0.8694932, 0.7911853, 0.08738397, 
    0, 0, 0,
  1, 1, 1, 1, 1, 0.01735635, 0, 0, 0.1874817, 0.9048839, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 0.5105418, 0.01035661, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.1085859, 0.8962955, 1, 0.9106531, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 0.8520856, 0.3672015, 0.313609, 0.2533256, 0.03519395, 0.3614787, 
    0.9965006, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9207106, 0.068037, 0, 
    0.3333627, 0.9408049, 0.8420026, 0.07602482, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.6269207, 1, 0.3631722, 0, 0, 0,
  1, 1, 1, 1, 0.7065716, 0.007449343, 0, 0, 0.8899581, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9990095, 0.6469289, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.302171, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 0.2509532, 0.7259984, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.4962145, 0.009399206, 0, 0.163563, 0.8311784, 0.2532057, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.6269538, 1, 0.7403622, 0, 0, 0,
  1, 1, 1, 0.9591063, 0.2903444, 0, 0, 0.3821371, 0.9899979, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8423643, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.1113189, 0.9288797, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 0.9148951, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.7166897, 0.193198, 0.378679, 0.7709084, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.2623808, 0.6417641, 0.1763478, 0, 0, 0,
  1, 1, 1, 0.4600145, 0, 0, 0.06470905, 0.7741343, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9729096, 0.4085401, 0, 0, 0, 0, 0, 0, 0, 
    0.09763272, 0.8372439, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.8914483, 0.9574527, 0.9569234, 0.6728632, 0.2309492, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 0.9083645, 0.1139706, 0, 0.006719753, 0.6425024, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.6623873, 0.3399824, 0, 0, 0, 0, 0, 
    0.01343901, 0.1122996, 0.2740395, 0.8126243, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9409829, 0.4917598, 0.01190909, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 0.5350372, 0, 0, 0.3691856, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.9817434, 0.7555508, 0.5806262, 0.721405, 0.9975661, 0.7792664, 
    0.03027645, 0, 0.05746033, 0.4528793, 0.6003847, 0.7402431, 0.8724493, 
    0.9833708, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0.9409539, 0.3217609, 0.0036727, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  1, 1, 0.5350789, 0, 0, 0.8339525, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.5068051, 4.62555e-05, 0, 0.01343513, 0.4826073, 0.6908599, 0.1210046, 
    0.6430895, 0.8287125, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9063402, 0.1092877, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 0.5351219, 0, 0, 0.9826248, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.6957842, 0.4102102, 0, 0, 0, 0.04356555, 0.1127979, 0.72868, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 0.9970281, 0.3331997, 0, 0, 0, 0.3913397, 0, 0, 
    0, 0, 0,
  1, 0.952481, 0.2011694, 0, 0, 0.9826218, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.8811629, 0.2063091, 0.1352319, 0.007285898, 0.3884326, 0.8899049, 
    0.8934386, 0.7892479, 0.9770009, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.9107391, 0.1889964, 0, 0.1838041, 0.8709035, 0.1881444, 0, 0, 0, 0,
  0.9999014, 0.380338, 0, 0, 0.4566294, 0.9974383, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 0.6904973, 0.03093301, 0.01432722, 0.6824431, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8582283, 0.03906883, 0.08034394, 
    0.7920045, 0.5992478, 0, 0, 0, 0,
  0.6594298, 0, 0, 0.3033189, 0.9943448, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.8270786, 0.08996841, 0.002212425, 0.4717253, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.7097963, 0.03884534, 0.4686598, 
    0.7735896, 0.07057529, 0, 0, 0,
  0.6233622, 0, 0.156587, 0.9117836, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.4757935, 0, 0.1331947, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 0.4924225, 0.007284605, 0.6021019, 0.1786143, 0, 0, 0,
  0.02644386, 0, 0.4743553, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9506161, 
    0.08966529, 0.03939142, 0.6957731, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8284553, 0.06092081, 0, 0, 0, 0, 0,
  0, 0.07934966, 0.98106, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.5513756, 0, 
    0.5253358, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 0.3725595, 0, 0, 0, 0, 0,
  0, 0.4350433, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9976279, 0.3553158, 
    0.6696817, 0.9791158, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 0.8894136, 0.02892898, 0, 0, 0, 0,
  0.01680065, 0.7740205, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9978701, 
    0.8976342, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 0.5902183, 0, 0, 0, 0,
  0.5105151, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8744972, 
    0.1220256, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9973416, 
    0.2167705, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9901414, 0.2867822, 
    0.3897793, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.816124, 
    0.1255585, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9809267, 0.9553849, 
    0.3948242, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.2193899, 0.1200667, 0, 
    0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.4875835, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.1584725, 0, 0, 0, 0, 0, 0,
  0.5802633, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.6097519, 0, 0, 
    0, 0, 0, 0,
  0.08221136, 0.7452577, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9897885, 
    0.9358599, 0.9987948, 0.7364435, 0, 0, 0, 0, 0,
  0, 0.7250001, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9684403, 0.774133, 
    0.3314505, 0.8281783, 0.9904674, 0.221187, 0, 0, 0, 0 ;

 zsurf =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.007482118, 
    4.885016, 6.027729, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.712759, 58.8956, 
    114.3027, 105.147, 66.36284,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.754428, 58.17822, 103.8941, 
    76.19964, 51.16923, 83.5846, 145.4227, 210.3575, 222.043, 166.9021, 
    138.0394,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12.60223, 150.9446, 238.0754, 281.3481, 
    288.7326, 300.3335, 276.3248, 277.1753, 296.433, 282.2253, 207.1847, 
    170.1954,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.971491, 107.903, 253.5528, 311.8893, 
    314.664, 349.46, 376.1395, 363.9048, 328.7521, 316.8185, 308.9201, 
    249.6144, 213.1554,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1077713, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.728832, 54.67075, 280.7457, 
    309.0462, 322.4052, 368.6298, 412.7725, 423.5071, 379.2067, 346.22, 
    351.7698, 329.3646, 274.3772,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.078801, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17.70223, 257.5212, 295.4054, 
    313.6127, 373.5954, 422.1055, 435.1128, 393.682, 374.0881, 409.6835, 
    409.2048, 354.9377,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26.2593, 246.0138, 296.1431, 348.5571, 
    410.7598, 429.6357, 435.3861, 395.7879, 402.5177, 442.4218, 430.7854, 
    398.5805,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 113.7163, 268.1346, 336.5029, 392.1589, 
    444.2632, 443.9155, 420.9473, 421.8472, 452.1077, 471.5658, 444.4251, 
    418.9319,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.859579, 200.0244, 305.7336, 330.6553, 
    391.9315, 444.2378, 439.8025, 441.541, 463.3921, 503.8092, 497.416, 
    462.6526, 441.0611,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14.25746, 228.6333, 312.2241, 361.2495, 
    416.0756, 482.3185, 484.5522, 484.6867, 507.3547, 509.7314, 483.8749, 
    461.7263, 442.7195,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.007934935, 91.5881, 260.8788, 351.2304, 
    404.0062, 456.2148, 509.2211, 528.7908, 527.3947, 511.4882, 494.72, 
    462.9256, 467.0975, 450.041,
  7.299402, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8.026843, 190.214, 291.695, 351.6114, 
    434.4432, 470.4533, 537.1084, 567.7097, 561.1059, 537.2833, 494.2285, 
    457.0371, 454.9888, 443.677,
  46.47058, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32.85493, 192.2326, 276.3241, 346.8046, 
    419.9743, 473.221, 539.5166, 587.4988, 579.1885, 551.3723, 502.3163, 
    438.6668, 426.6781, 416.2831,
  56.36044, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2935236, 29.53243, 141.496, 253.5633, 
    345.4431, 426.5362, 485.1349, 548.7592, 600.852, 588.0337, 535.9756, 
    460.5315, 394.231, 382.3351, 380.9086,
  39.45049, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32.83228, 53.73461, 1.585332, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3.041326, 10.00888, 
    106.9153, 227.8007, 348.7626, 445.4996, 478.5939, 575.4977, 600.4197, 
    570.2203, 506.0541, 415.3415, 330.4285, 332.2667, 343.1945,
  13.59347, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26.08635, 195.4105, 256.4257, 146.537, 
    55.481, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.186994, 
    18.06586, 130.0469, 253.3653, 363.8199, 394.896, 513.6748, 590.4353, 
    558.9642, 518.7917, 454.3615, 363.8717, 303.3865, 300.713, 321.3069,
  0.9656757, 0, 0, 0, 0, 0, 0.03586638, 0, 0, 0, 49.68565, 326.9774, 
    455.3936, 576.6316, 425.3625, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.01508173, 21.43529, 144.3786, 255.7441, 319.1965, 459.2542, 
    569.7118, 604.0175, 513.782, 425.8328, 371.0454, 316.678, 281.3964, 
    295.9887, 312.7417,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 188.9793, 461.0893, 744.1964, 857.3239, 
    577.0432, 10.22077, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    28.41998, 89.48728, 170.1808, 341.458, 487.3284, 552.6357, 471.7288, 
    351.3307, 336.5912, 295.8323, 257.3056, 256.7657, 275.5327, 266.8901,
  14.46666, 0, 0, 0, 0, 0, 0, 0, 0, 0, 98.10371, 430.0524, 658.2639, 
    869.6558, 593.5727, 27.91763, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 28.79319, 27.47902, 102.3828, 250.1567, 353.9292, 297.6356, 
    194.349, 196.082, 204.2073, 194.9052, 184.4335, 186.8029, 202.2491, 
    201.6232,
  63.77672, 3.367655, 0, 0, 0, 0, 0, 0, 0, 0, 20.47009, 226.3262, 481.9063, 
    847.3206, 850.9589, 97.98926, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 5.864242, 1.030459, 11.5586, 92.8717, 81.6533, 37.3248, 
    45.25832, 55.12968, 71.40536, 80.22321, 109.8221, 156.4528, 158.7244, 
    139.6773,
  92.77831, 10.55024, 0.7231424, 0, 0, 0, 0, 0, 0, 0, 0.06683189, 88.24445, 
    325.958, 897.7953, 1142.866, 334.1817, 0.2153307, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.6444512, 1.022004, 0.2444094, 0, 
    0.1744056, 0, 0, 11.61093, 95.71937, 140.5593, 109.8717, 89.47809,
  148.8612, 111.2776, 10.43683, 0.2487843, 0, 0, 0, 0, 0, 0, 0, 26.9947, 
    302.4542, 900.6857, 1410.459, 722.3347, 26.92253, 0, 0, 0, 0, 0, 0, 
    0.2948902, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.04675792, 32.30137, 73.17574, 45.04506, 113.3446,
  356.8611, 272.9169, 144.0292, 36.66886, 4.051232, 0, 0, 0, 0, 0, 
    0.00622688, 95.44665, 402.4702, 1000.551, 1468.909, 1068.681, 138.7007, 
    0, 0, 0, 0, 0, 0, 224.4563, 0.7204035, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 40.79513, 46.98636, 44.90553, 135.4555,
  607.5697, 617.0065, 415.9779, 222.5245, 82.16385, 13.76159, 0, 0, 0, 0, 
    0.7036354, 167.195, 549.0036, 865.797, 1297.997, 1084.883, 386.271, 0, 0, 
    0, 0, 0, 0, 0, 0, 38.47579, 1.349345, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.05735796, 3.489815, 17.0652, 91.46315,
  805.8144, 689.3148, 665.8074, 521.1199, 295.9792, 99.36646, 9.087084, 0, 0, 
    0.005802704, 0.3102686, 111.6922, 363.4742, 565.2116, 806.0615, 1016.094, 
    629.3563, 16.26268, 0, 0, 0, 0, 0, 0, 0, 0, 0.02296036, 0, 0, 0, 0, 
    1.214581, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002000303, 0.005462797, 
    18.32721,
  760.7727, 661.396, 709.6733, 604.6326, 464.2514, 283.1679, 79.76301, 
    0.1074248, 0, 0, 0, 17.74922, 148.9407, 173.6682, 402.7549, 729.6694, 
    723.2713, 46.89246, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1074003,
  860.9228, 736.6833, 628.5461, 564.9741, 466.655, 335.0508, 169.4657, 
    9.562907, 0, 0, 0, 0, 7.39888, 15.74615, 103.3149, 461.4926, 652.2623, 
    214.472, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, -0.0001159482, 0, 0,
  954.5076, 825.0037, 642.887, 541.5004, 467.5988, 374.7963, 167.8485, 
    1.774008, 0, 0, 0, 0, 0, 0.3348222, 19.11695, 171.6814, 741.9515, 
    374.4197, 25.98872, 0, 0, 0, 0.0003252521, 0, 0, 0, 0, 0.001458651, 
    7.516816e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  858.3884, 673.0359, 533.1504, 448.0885, 424.8119, 345.4697, 166.7318, 0, 0, 
    0, 0, 0, 0, 0, 0.567318, 193.9483, 883.2621, 655.3737, 12.50792, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.0002288724, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.005102882, 0, 0,
  765.3333, 667.6134, 488.7987, 363.019, 313.4333, 341.2213, 122.4717, 0, 0, 
    0, 0, 0, 5.00687, 0, 0, 60.76902, 616.8209, 406.96, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  892.0968, 795.8924, 625.4323, 432.2025, 321.9835, 331.9277, 130.2014, 
    0.004251794, 0, 0, 57.24534, 20.8572, 0.7291545, 0, 0, 0, 119.2905, 
    99.81622, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 13.85986, 0.004370535, 0,
  1001.771, 792.1298, 674.5222, 541.9408, 384.3335, 350.6531, 103.3347, 
    0.1868827, 0, 0, 18.48727, 0, 0, 0, 0, 0, 9.2637, 4.286283, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.02841037, 
    1.063279, 1.850597, 3.574715, 3.295839, 153.8647, 199.7177,
  1318.781, 598.8708, 526.7117, 510.9486, 354.2004, 223.6784, 15.55483, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.01238247, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10.38296, 174.51, 148.3694, 0, 0, 0, 
    148.5062, 285.8834,
  1220.16, 848.2032, 380.6071, 390.465, 259.5177, 95.94141, 0, 0, 0, 0, 0, 0, 
    0, 0.01723676, 0.0002739781, 0.009286015, 0, 0, 0, 0.006633122, 0, 0, 0, 
    0, 0.003201818, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001933358, 
    0, 0, 0, 0, 0, 0, 0, 0, 2.528343, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.01048129, 0, 35.29255, 81.26061, 161.3701, 172.8166, 125.7769, 
    60.08969, 51.96622, 164.8291,
  1338.663, 964.2402, 591.19, 291.6062, 139.8224, 33.77381, 0.002896692, 0, 
    0, 0, 0, 0, 0, 0.09759907, 0, 0, 0, 0, 0.003041361, 0, 0, 0, 0, 0, 
    0.003417519, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.214117, 10.05566, 31.4626, 
    198.6635, 257.3435, 200.3842, 110.9841, 79.73378, 263.6654, 36.78745, 
    1.378057, 31.15954, 8.130059, 1.005422,
  1026.086, 1045.23, 716.394, 366.1234, 142.9799, 30.33171, 0.4619157, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10.88786, 
    115.5257, 170.2808, 339.2503, 395.8933, 151.5352, 149.8366, 27.3561, 
    4.022614, 20.95062, 0, 0, 3.260029, 1.872875, 0.0508271, 0, 0, 0,
  974.4459, 1067.982, 927.8552, 494.0284, 130.0466, 22.65291, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.899872, 139.8198, 
    115.3161, 168.5896, 352.7554, 266.0829, 177.1721, 131.6926, 43.10759, 
    1.240668, 4.394837, 0.006916575, 0.0003986534, 0.0104446, 0.0172614, 0, 
    2.609623, 0, 0.001365404, 0.09803439, 0.2262536, 0.004817449,
  1204.486, 1237.256, 1141.603, 688.0075, 263.0531, 10.36784, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001947393, 0, 0, 0, 0.01043915, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01680503, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.04407993, 32.09272, 400.8964, 597.5397, 333.6716, 124.2354, 104.7639, 
    67.59129, 23.81756, 3.731113, 1.087241, 0, 0, 0, 0, 0, 0, 4.881635, 
    10.31701, 0, 6.561506, 40.6811, 3.38201, 0.01358287,
  1440.196, 1303.7, 1187.572, 799.9657, 447.4943, 28.87032, 0.287935, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.008367683, 0, 0.0005597501, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.006913288, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 17.87501, 27.6564, 41.68385, 40.07766, 2.412819, 0, 0.3703949, 0, 0, 
    2.694052, 0, 0.06298108, 0, 0, 0.007401017, 0.01018163, 0.5245222, 
    314.3598, 25.13958, 10.84065, 64.80965, 69.94651, 0.2126305, 0,
  1507.507, 1338.634, 1162.16, 895.2739, 556.3425, 113.5388, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.003531589, 0, 0.3608332, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.645804e-05, 0.008660849, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.399279, 1.708197, 228.0259, 260.7763, 73.72216, 0.01350134, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.04154294, 0.6853305, 0.0007041242, 0, 0, 0, 222.6289, 
    19.51247, 152.801, 98.75947, 68.60026, 0, 0,
  1593.552, 1288.948, 1293.234, 1037.663, 604.3491, 220.0716, 11.92896, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3.231213, 0.1002754, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.003929192, 0.06615317, 
    326.9998, 382.6881, 215.296, 6.51867, 0, 0, 0.0005210711, 0, 0, 0, 
    0.00945402, 0, 0.04497931, 26.08819, 57.13885, 7.390703, 0, 0, 69.87069, 
    559.0273, 111.9894, 624.2891, 262.6683, 1.642632, 0, 0,
  1658.693, 1261.843, 1404.586, 1067.003, 563.8726, 182.1493, 36.27239, 
    0.3323672, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002778716, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3.277349, 3.089526, 
    220.2578, 271.9154, 232.9942, 11.41514, 6.090748, 2.68348, 5.510962, 
    3.529593, 0, 1.621469, 5.491666, 9.77548, 7.35185, 3.514773, 53.89715, 
    161.2589, 24.12606, 0, 0.007201126, 433.8056, 1036.646, 400.0064, 
    500.544, 149.6249, 0, 0, 0,
  1645.619, 1472.14, 1404.025, 1096.18, 483.7211, 188.2313, 50.92135, 
    15.02244, 0.3012842, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9.016459, 125.5137, 
    477.9677, 315.6645, 11.36371, 6.38086, 10.82686, 9.825094, 2.584005, 
    0.8772991, 0, 14.4698, 70.73858, 64.99486, 20.69061, 17.08455, 32.61346, 
    164.0018, 34.12597, 0.002215982, 0, 41.34579, 1159.648, 903.4078, 
    550.6257, 25.76042, 12.09169, 7.678148, 124.0715,
  1967.175, 1791.275, 1808.567, 1089.094, 523.5789, 218.3327, 97.51249, 
    52.39918, 11.84871, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26.70954, 0.01252906, 
    573.1802, 456.6572, 67.73898, 16.5005, 4.31343, 5.305326, 0.0450154, 0, 
    0.8252385, 6.159415, 65.49741, 194.1909, 179.5106, 157.9093, 77.64091, 
    91.67677, 141.2131, 99.64323, 8.659935, 0, 4.571824, 614.8233, 532.0992, 
    483.2188, 457.6458, 209.052, 8.435591, 0,
  2024.533, 2181.229, 2001.106, 1283.735, 528.7686, 242.7618, 136.9167, 
    79.82225, 23.44122, 3.95113, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.004921097, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.6401625, 
    6.308005, 158.2323, 422.013, 185.8305, 17.01043, 4.866463, 8.841109, 
    0.001300426, 0, 0, 0, 11.91, 84.76138, 176.0108, 242.7657, 291.476, 
    330.5183, 200.2534, 138.5459, 34.58592, 22.24334, 0, 0, 144.1948, 0, 
    6.173299, 15.85019, 45.24471, 0.213134, 0,
  1923.579, 1771.256, 1778.076, 1070.793, 505.6136, 241.9928, 148.163, 
    76.44843, 32.30178, 17.09214, 7.496256, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01376197, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.004098975, 22.05864, 72.32189, 406.9106, 296.7709, 13.30871, 10.29677, 
    4.396094, 1.765978, 0, 0.01962267, 0.09792335, 0.3374118, 51.71622, 
    88.17578, 76.92102, 159.3824, 380.0949, 535.228, 499.3378, 330.4606, 
    165.3464, 41.27188, 2.509667, 0.02632017, 117.6165, 245.3032, 188.3384, 
    112.4978, 172.8582, 310.4585, 94.6843,
  1794.133, 1276.998, 1319.927, 847.228, 358.8172, 233.8158, 187.9514, 
    116.8452, 68.52618, 71.37233, 45.78811, 16.83432, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.009340961, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2.670939, 25.97792, 355.1271, 272.5902, 27.50756, 10.82965, 
    10.10394, 20.80869, 2.207196, 0, 0.004632319, 0.4954259, 0, 54.69146, 
    103.1393, 87.46021, 162.231, 378.5865, 622.8563, 789.714, 748.1737, 
    514.2153, 211.2245, 106.0069, 43.93421, 0, 117.153, 217.9034, 176.2699, 
    56.00568, 72.75879, 291.925,
  1122.184, 817.0998, 942.5208, 629.3625, 367.3386, 319.362, 310.6506, 
    233.7132, 219.4219, 172.6176, 170.9612, 87.88506, 52.56012, 6.837942, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.01282556, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.003567874, 9.907857, 7.509503, 341.4931, 669.8797, 266.7873, 
    11.2073, 57.75204, 56.43156, 49.87582, 0.7429065, 0.01104457, 0.2828173, 
    0, 0.04069449, 4.1862, 0.06066301, 11.07728, 86.06728, 187.3697, 
    479.2986, 762.8614, 937.4857, 601.6578, 195.3882, 27.83612, 0.1914168, 0, 
    0, 0, 0, 0, 0, 11.51637,
  846.5782, 504.4499, 654.7703, 570.2628, 501.0254, 542.6677, 483.9015, 
    424.1021, 332.9808, 314.234, 333.5416, 253.9334, 130.1149, 111.9619, 
    7.31144, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.0009155833, 0.003754308, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.204808, 504.0269, 598.7817, 428.9163, 
    11.3934, 12.47365, 231.9589, 136.3775, 6.838151, 0, 2.634708, 3.781463, 
    0.1162148, 0.6912898, 0.01993117, 0, 0.4706172, 7.387184, 44.55817, 
    244.1146, 594.9794, 933.8558, 513.5035, 77.61767, 4.361522, 0, 0, 0, 0, 
    0, 0, 0, 0,
  681.6527, 442.5084, 578.8173, 717.4026, 922.1249, 813.6738, 759.1872, 
    525.2695, 321.9953, 302.5872, 458.9889, 403.1359, 243.0368, 181.6122, 
    107.4319, 9.799197, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.0001312634, 0.006848679, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.3214408, 335.2546, 813.2599, 438.9796, 
    1.541609, 0.004860971, 141.2879, 433.2815, 256.4115, 14.89001, 0, 0, 0, 
    0.1404909, 6.80957, 0, 0, 0, 0, 0.4797853, 35.22785, 388.0224, 854.2148, 
    528.0695, 83.28231, 2.967625, 0, 0, 0, 0, 0, 0, 0, 0,
  545.9903, 500.1561, 701.9286, 1102.757, 1219.171, 1147.172, 956.5318, 
    675.6527, 331.725, 351.9229, 475.9785, 420.0756, 313.623, 228.7287, 
    180.0209, 134.015, 0.3182439, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01651771, 0, 0, 0, 0, 0, 0, 22.53872, 
    0.65847, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30.20723, 195.3939, 
    90.67072, 4.860431, 0, 5.169554, 264.6625, 416.897, 223.7468, 2.467426, 
    0, 0, 0, 0.01299047, 0.1073577, 0, 0, 0, 0, 0, 2.723956, 80.23975, 
    657.4532, 634.125, 285.9821, 125.6809, 2.169004, 0.1452292, 0, 0, 0, 0, 
    0, 0,
  575.7665, 549.1124, 1004.394, 1257.504, 1520.269, 1214.792, 1053.349, 
    760.7601, 506.7095, 417.5125, 432.6968, 399.7943, 364.9707, 304.9736, 
    209.8668, 138.7341, 27.90703, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001978899, 0.02694878, 0, 0, 0, 0, 0, 
    7.94479, 361.0423, 148.2079, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3.387879, 
    0.004412269, 0, 0, 0, 1.012016, 28.95815, 159.6374, 162.7487, 6.871452, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002113436, 123.6737, 502.31, 
    321.5427, 69.19288, 34.57666, 4.016514, 0.6476752, 0, 0, 0, 0, 0,
  771.0378, 731.9822, 1232.212, 1579.218, 1810.72, 1665.98, 1247.325, 
    891.9006, 552.7863, 534.0606, 470.0626, 487.2615, 500.9968, 399.5934, 
    301.6216, 216.2957, 101.2677, 1.366401, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7.578414, 0, 10.02934, 
    217.377, 48.73487, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2398228, 7.076045, 0, 
    0, 0, 0.5435731, 5.565549, 79.59003, 18.13072, 1.341174, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.07269884, 342.0459, 154.1556, 9.21379, 
    0.01240786, 0.0236598, 5.468072, 10.2199, 0.1744068, 0, 0, 1.12455,
  1005.523, 1089.269, 1428.493, 1729.941, 2157.611, 2366.877, 1791.208, 
    1172.936, 789.075, 679.2053, 769.5369, 774.6565, 661.5249, 538.7116, 
    499.1805, 452.9259, 318.8668, 107.7354, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.003257784, 0, 0, 14.33969, 
    269.4527, 18.4388, 2.629723, 63.20306, 3.818854, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.4436082, 0.4391197, 0, 0, 0, 11.42085, 94.30405, 98.075, 
    0.03083581, 0, 0, 0, 0.03971905, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9.149135e-05, 
    0, 0, 9.795963, 11.95197, 0.4926467, 0.0001121615, 0, 0.0542269, 
    0.1652767, 35.90819, 0, 61.54511, 395.5136,
  1443.506, 1620.422, 1765.2, 1789.817, 2168.043, 2356.399, 1999.072, 
    1344.355, 974.863, 966.6523, 1036.74, 970.4948, 807.8265, 729.062, 
    640.0353, 622.3807, 558.9814, 343.8018, 29.92353, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0003971517, 0.002529405, 0, 0, 
    121.7922, 429.6986, 193.016, 6.398975, 3.334329, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.2867806, 0, 0, 0, 0, 3.61325, 129.9913, 54.15724, 0, 0, 0, 
    0.1055335, 0.3423316, 0.3816859, 0.8894814, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3.002282, 0, 0, 0, 0, 0, 91.78906, 15.18766, 64.01128, 362.9198,
  1620.956, 2030.3, 1884.991, 2049.509, 2068.68, 2175.013, 1586.164, 
    1522.586, 1346.341, 1360.391, 1342.486, 1150.649, 1009.675, 798.4236, 
    803.64, 793.613, 751.2167, 539.5749, 185.2117, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.00889502, 0.008948714, 0, 1.305878, 
    327.1373, 460.4203, 183.9435, 19.73282, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.001868226, 3.177953, 0, 0, 0, 0, 5.91536, 94.78001, 1.925256, 0, 0, 
    0.02996243, 4.757724, 2.262005, 0.8893167, 0.6945848, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 38.47111, 40.73141, 0, 0, 0, 0, 68.93193, 198.6472, 
    337.3564, 558.7494,
  1649.085, 1708.983, 1942.575, 2064.672, 2304.163, 2042.305, 1346.739, 
    1341.973, 1536.301, 1614.115, 1351.418, 1085.79, 943.1578, 900.9448, 
    952.3292, 1066.381, 834.631, 657.6016, 280.5684, 3.45371, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001200154, 0.001476862, 0, 
    152.6915, 685.7798, 660.864, 391.5136, 81.102, 0.08322787, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.1983324, 8.214144, 0, 0, 0, 0, 7.976196, 96.0976, 
    32.68804, 0, 0, 11.5986, 136.4807, 24.27074, 1.852875, 7.053572, 
    56.97015, 4.038934, 0.03956408, 0, 0, 0, 0, 0, 9.457328e-05, 0, 0, 
    0.1137195, 89.28968, 12.82965, 0, 0.000534966, 0, 0, 46.44008, 85.76493, 
    411.291,
  1466.144, 1621.266, 1631.515, 2122.453, 2175.795, 2267.993, 1097.97, 
    824.9056, 896.3997, 932.9909, 568.8134, 122.1493, 139.7222, 230.9751, 
    585.2339, 743.4264, 595.6318, 653.7233, 457.3597, 15.86434, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.980672, 440.7948, 
    848.3855, 797.6866, 593.3608, 199.7116, 8.479733, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 11.56622, 0.1151541, 0, 0, 0, 11.44357, 154.1412, 126.2073, 
    0.02027015, 0.8643358, 204.4469, 257.3035, 118.653, 15.25982, 90.17926, 
    348.3282, 451.6818, 20.03893, 0, 0, 0, 0, 0, 0.0003784416, 0, 0, 0, 
    0.3295275, 73.48798, 1.209638, 0.001240408, 0.04867897, 35.55901, 
    205.4684, 37.47905, 55.50045,
  1265.107, 1271.335, 1965.781, 1997.247, 2257.103, 2371.452, 1157.836, 
    568.8094, 507.9307, 527.9256, 61.88685, 0, 0, 0, 0, 0, 0, 0, 25.08505, 
    2.611548, 1.012719, 54.77631, 55.46979, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 56.8435, 558.8643, 753.3204, 685.9753, 529.2399, 
    221.9993, 6.638701, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.390496, 0.1437027, 
    0, 0, 0, 5.025319, 296.0272, 133.192, 26.48146, 105.7203, 124.3082, 
    133.4471, 18.79172, 41.91351, 168.925, 502.5459, 687.1468, 145.1467, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 9.612703, 23.07717, 0.1670243, 0.3258666, 
    40.60841, 178.4189, 98.15704, 58.47993,
  935.9797, 1371.701, 1933.655, 2314.278, 2206.839, 2331.325, 1047.749, 
    519.5513, 454.4148, 405.1205, 26.92118, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 244.4359, 
    576.6982, 579.9873, 438.5885, 334.7599, 131.4858, 3.241302, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.0453538, 0.0158177, 0, 0, 0, 75.12135, 375.2448, 
    88.78672, 19.92136, 145.9868, 126.3988, 55.09162, 79.25726, 93.2966, 
    89.02313, 311.1271, 517.6355, 122.5172, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.03161435, 9.429642, 0.6056394, 0.146424, 207.0213, 126.4081, 45.91529, 
    85.9324,
  705.9424, 1077.602, 1789.276, 2157.059, 2121.644, 2145.599, 927.7297, 
    349.9645, 414.1831, 239.4039, 205.0616, 535.8789, 337.7988, 224.2843, 
    93.21812, 12.07225, 4.108486, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21.81651, 480.2482, 616.3601, 509.2854, 
    411.6318, 353.8981, 172.9756, 23.66262, 1.744636, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.001127199, 0.426254, 0.06272013, 0, 158.0811, 521.639, 
    141.0725, 99.96737, 247.5734, 203.0635, 144.6472, 146.9874, 146.9239, 
    291.5794, 505.7589, 561.468, 82.04576, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7.754673, 7.457764, 24.7692, 42.12467, 9.055123, 4.078703, 80.82257,
  560.522, 873.38, 1472.261, 1866.38, 1992.183, 1959.356, 668.1165, 250.8919, 
    291.7672, 17.91137, 626.5022, 1631.719, 1588.758, 1237.268, 972.5966, 
    822.8162, 666.3598, 231.6238, 95.20377, 24.35091, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 93.28631, 598.2587, 574.9574, 
    508.1927, 475.7988, 445.4901, 244.6739, 75.22868, 59.67073, 26.13394, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 7.006592, 9.506021, 2.820326, 1.543359, 
    144.5288, 485.7056, 157.8752, 139.0608, 306.2983, 182.6353, 140.4857, 
    150.7803, 237.6682, 550.9364, 811.1963, 598.2958, 25.34849, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 140.1268, 241.5589, 39.90154, 11.41144, 38.09826, 
    75.28021,
  520.9725, 685.0739, 1104.142, 1548.977, 1849.273, 1977.533, 530.145, 
    203.5752, 23.72789, 27.13107, 956.7662, 2034.414, 1627.404, 1195.415, 
    1080.397, 1104.885, 1093.357, 887.1946, 732.5614, 442.7809, 42.32203, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 227.5572, 
    614.1383, 604.0764, 532.1347, 527.2681, 501.3772, 266.3045, 197.5267, 
    319.5226, 439.0925, 52.55056, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01218646, 
    68.76542, 10.88835, 49.6851, 244.7333, 434.6059, 156.4234, 331.7645, 
    396.8661, 241.47, 169.5624, 150.5604, 254.91, 544.6859, 578.8292, 
    122.1243, 0.04935317, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.776042, 
    88.48724, 86.04845, 37.06418, 36.67148, 83.62952, 1.168923,
  520.364, 623.9707, 845.1304, 1182.964, 1794.826, 1631.395, 245.3956, 
    30.59338, 0.1295522, 65.68732, 1191.472, 1929.175, 1380.801, 898.722, 
    945.2995, 1004.129, 951.7753, 889.402, 807.7346, 725.3493, 650.4291, 
    576.4832, 399.0143, 189.4995, 1.069616, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 290.6859, 650.6129, 587.6777, 538.5913, 469.5362, 
    367.0397, 239.3359, 267.2038, 520.4188, 582.6263, 354.7753, 95.80848, 0, 
    0, 0, 0, 0, 0, 0, 0, 10.50261, 205.8622, 156.8265, 367.9012, 536.3768, 
    554.2907, 339.4029, 439.8899, 418.0555, 214.6228, 185.1647, 265.1077, 
    310.9288, 294.0193, 49.32493, 0, 0, 0, 0.0004447775, 0.0008141641, 
    0.0001843075, 0, 0, 0, 0, 0, 0.00153388, 0, 9.762164, 91.66759, 151.5858, 
    43.30084, 69.43888, 56.62251, 23.58093,
  527.755, 558.0959, 777.8425, 1038.259, 1442.285, 857.6389, 34.7822, 
    0.06794915, 0.1317989, 65.86896, 1226.782, 1676.783, 1155.866, 959.6856, 
    863.8164, 851.5259, 757.8932, 699.1624, 691.1156, 647.6199, 588.8004, 
    448.2683, 337.8521, 251.0181, 128.1548, 0.6675929, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1.583894, 274.4207, 587.1978, 539.9442, 498.1378, 
    401.8043, 324.701, 235.9535, 351.3758, 472.5636, 586.2536, 372.6698, 
    260.64, 20.91498, 0.5449734, 0, 0, 0, 0, 0, 0.1160287, 111.142, 209.0083, 
    276.4948, 646.7979, 765.1041, 724.9354, 477.4805, 577.1857, 463.0179, 
    431.689, 425.1302, 450.4791, 382.4208, 78.48548, 0, 0, 0, 0, 0, 
    0.003998051, 0.002220947, 0, 0, 0, 0, 0, 0, 0, 105.1281, 169.7474, 
    236.0875, 9.81155, 0.1445957, 0, 0,
  489.275, 506.2431, 635.707, 891.2947, 1140.819, 104.9125, 0.5735672, 
    0.0001255112, 2.393601, 199.3139, 1536.486, 1511.392, 1079.511, 820.4056, 
    728.9279, 624.3528, 521.0572, 428.4595, 417.1996, 391.4514, 321.5363, 
    234.6511, 206.3434, 187.8103, 161.0246, 103.9707, 3.567678, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 4.888042, 22.56903, 1.230958, 202.7648, 429.525, 
    412.595, 342.0215, 395.2505, 348.6987, 285.1621, 336.5508, 375.4762, 
    287.4457, 307.1478, 204.0902, 144.1289, 12.40784, 0, 0, 0, 0, 0.09297946, 
    48.31137, 410.1348, 219.7555, 321.0481, 912.0163, 957.0075, 782.5162, 
    689.6246, 672.2351, 803.3319, 900.5595, 921.7489, 653.4254, 113.7043, 0, 
    0, 14.97981, 163.9573, 16.21266, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34.01518, 
    399.7357, 415.947, 11.40101, 0, 0, 0,
  423.9285, 419.6786, 540.4236, 810.2414, 880.0971, 25.37736, 0, 0, 43.69834, 
    958.8488, 1720.627, 1412.165, 928.663, 770.8799, 633.066, 510.455, 
    402.9467, 319.4293, 278.5269, 235.3018, 194.7553, 149.0402, 112.7481, 
    124.9141, 133.1899, 112.3536, 20.9965, 2.64545, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2.267793, 70.71137, 122.5515, 31.54795, 87.75684, 313.0298, 326.2078, 
    392.7047, 459.9867, 517.2142, 481.4169, 442.511, 390.7699, 276.8941, 
    289.5733, 344.4179, 305.1668, 167.0574, 9.916601, 1.032431, 1.048887, 
    0.2411555, 23.19702, 397.0361, 721.8358, 320.7461, 332.2949, 979.869, 
    1030.202, 931.765, 809.9, 823.1024, 793.5685, 951.8102, 1033.525, 
    719.0648, 119.1517, 0.833892, 0, 14.80536, 271.7417, 152.8016, 
    0.00275539, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 621.5582, 558.1843, 245.3577, 
    0, 0, 0,
  389.9949, 432.4892, 525.9587, 618.4981, 485.3033, 0.03390811, 0, 1.35604, 
    605.9611, 1549.469, 1794.849, 1175.007, 871.842, 714.1773, 567.928, 
    445.1647, 359.2397, 288.548, 230.5943, 181.9214, 144.2462, 113.5117, 
    92.68795, 83.6313, 99.99515, 113.782, 90.98781, 80.63214, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 10.24857, 59.58021, 91.44401, 35.23301, 92.64501, 269.2377, 
    433.9703, 408.1391, 449.0736, 489.8803, 490.6386, 587.921, 538.6768, 
    542.0423, 504.0613, 493.4232, 387.6947, 149.3013, 21.24825, 2.08333, 
    3.27737, 3.702941, 63.49332, 591.3827, 870.5641, 260.2408, 218.9506, 
    877.173, 980.9655, 1040.86, 1143.761, 991.8488, 921.4819, 835.4803, 
    934.3461, 614.5713, 122.0434, 14.56706, 2.029026, 0, 21.34945, 37.91715, 
    4.003912, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 419.2063, 402.9444, 268.8748, 0, 
    0, 0,
  431.8418, 536.3006, 574.058, 315.8998, 41.75761, 0, 0, 59.75841, 954.189, 
    1557.024, 1298.473, 942.2996, 752.2569, 616.2059, 486.4283, 377.0709, 
    312.1561, 255.6407, 198.0654, 142.262, 116.617, 107.7247, 90.60133, 
    80.00478, 98.95425, 307.284, 343.9886, 272.9455, 6.16348, 0, 0, 0, 0, 0, 
    0, 0, 2.050448, 40.84933, 34.03916, 33.79316, 71.37947, 217.7432, 
    315.7126, 443.3457, 437.9484, 458.0936, 444.2867, 431.0873, 447.9553, 
    504.2306, 471.0587, 559.8055, 493.2112, 392.4747, 196.1293, 47.81644, 
    8.629056, 4.509862, 7.082555, 123.9592, 629.7461, 843.9626, 281.6333, 
    305.7295, 690.8347, 1054.628, 1119.722, 1335.16, 1190.468, 1065.214, 
    984.9171, 869.7607, 546.3845, 225.0289, 150.4363, 163.5934, 3.164987, 
    1.992715, 22.49724, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 167.7594, 192.5879, 
    127.9389, 0, 0, 0,
  464.4328, 710.1633, 619.1936, 47.74748, 0.006608745, 0, 1.039034, 425.7875, 
    1205.512, 1296.795, 937.6955, 818.3823, 688.7088, 615.1889, 470.3323, 
    343.0821, 270.3759, 214.7289, 163.605, 112.6529, 104.0565, 122.8048, 
    107.724, 95.03403, 378.6848, 553.5956, 557.1316, 213.1545, 0, 0, 0, 0, 0, 
    0, 0, 3.253178, 4.987194, 15.42553, 23.11442, 53.14434, 198.1807, 
    390.6396, 476.5912, 416.6757, 370.3962, 423.6606, 388.2758, 315.9665, 
    300.9809, 279.9049, 272.6179, 240.4554, 254.8682, 231.5103, 158.6761, 
    75.81209, 21.71908, 9.130775, 31.90206, 180.6022, 519.5223, 818.9929, 
    367.1069, 232.1573, 540.9075, 1020.897, 1331.289, 1515.057, 1429.161, 
    1326.372, 1300.804, 1167.494, 857.9363, 537.9557, 430.6571, 235.6319, 
    105.8424, 52.64319, 52.60298, 48.16794, 5.177803, 0.0127918, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 7.925615, 7.623189, 0, 0, 0,
  541.9563, 702.7642, 525.0195, 0.008912559, 0, 0.7958623, 220.1246, 
    1012.623, 1381.692, 1054.735, 911.1928, 865.9833, 754.9418, 683.0833, 
    507.5714, 339.2844, 241.6909, 185.5594, 133.8963, 81.90056, 93.08733, 
    116.5835, 104.0461, 220.4304, 362.2358, 272.5128, 22.4466, 0, 0, 0, 0, 0, 
    0.464163, 2.217875, 1.132218, 118.9751, 48.45937, 24.96659, 68.75862, 
    119.5871, 168.0666, 359.0999, 420.4307, 372.978, 292.5229, 326.5298, 
    261.4095, 174.0229, 145.3442, 113.1015, 90.15494, 74.61478, 49.53991, 
    51.27683, 45.57203, 19.36777, 16.3014, 20.58949, 212.4812, 371.5741, 
    567.3152, 837.6189, 773.0519, 254.7844, 402.2862, 1117.507, 1593.182, 
    1713.899, 1657.007, 1585.993, 1660.75, 1626.9, 1297.729, 1008.488, 
    628.0763, 368.5419, 180.6032, 125.0678, 198.4454, 235.6197, 149.7811, 
    32.02615, 2.138504, 0.001609906, 0, 0.0001999206, 0, 0, 0, 0, 0, 
    0.04724865, 3.110864, 0, 0, 0,
  549.2347, 686.2816, 401.375, 0, 0, 65.01826, 822.366, 1329.428, 1219.403, 
    975.2758, 969.5549, 932.9362, 803.3354, 731.2571, 572.4413, 387.7809, 
    255.709, 181.6068, 113.3861, 42.95264, 32.65179, 33.98416, 38.83173, 
    138.7656, 318.7718, 0.7992804, 0, 4.0433, 27.02569, 43.15045, 65.88136, 
    171.93, 328.6717, 326.6402, 310.495, 300.1921, 112.6526, 39.34247, 
    116.7174, 196.2544, 210.7351, 281.5956, 376.5725, 369.3636, 290.0414, 
    245.2731, 172.5113, 134.9192, 115.1656, 85.47749, 72.11951, 66.97635, 
    58.92198, 81.27972, 173.3912, 214.537, 108.2215, 198.1225, 218.5382, 
    378.2805, 263.0815, 752.1837, 870.6851, 687.0273, 413.0518, 1141.952, 
    1943.944, 2054.098, 1926.115, 1828.285, 1968.703, 1788.26, 1402.79, 
    904.152, 675.1245, 442.3218, 270.6985, 164.4036, 201.3591, 233.2095, 
    139.005, 55.39569, 31.88385, 19.8936, 0, 0, 0, 0, 0, 0, 0, 0.36459, 
    2.782869, 0, 0, 0,
  535.8906, 600.8014, 335.9744, 0, 0, 154.2405, 912.732, 1109.16, 989.4586, 
    950.7682, 958.7252, 936.9157, 774.5905, 743.4534, 586.5957, 444.2589, 
    308.8711, 197.4996, 96.48969, 12.3244, 0.1483047, 0.03790293, 0.1436228, 
    37.92851, 155.9851, 30.76747, 221.6138, 252.8131, 416.8718, 624.1976, 
    699.0229, 728.5979, 841.8627, 953.5579, 886.6041, 601.1133, 92.53477, 
    32.85394, 103.7375, 188.0701, 216.8431, 268.9015, 362.442, 393.7513, 
    334.8778, 224.5274, 158.4746, 126.387, 112.2802, 112.7532, 257.5196, 
    397.1968, 538.8138, 1240.1, 2032.906, 2200.138, 2236.536, 1966.697, 
    1706.219, 1459.807, 783.1836, 362.6883, 642.8234, 493.0027, 840.9872, 
    1130.427, 2271.913, 2496.004, 2172.94, 1901.212, 2118.338, 2085.24, 
    1574.87, 1081.068, 810.9539, 635.4389, 423.6662, 250.8699, 288.964, 
    307.7717, 284.6146, 159.4874, 139.9633, 136.567, 123.2743, 19.75318, 0, 
    0, 0, 0, 0, 0, 0.3498602, 0, 0, 0,
  617.859, 478.8044, 162.5502, 0, 0.316467, 273.1028, 967.5567, 1024.078, 
    960.9479, 962.3912, 987.4086, 923.9738, 816.1489, 736.3137, 601.2943, 
    460.8235, 324.0718, 168.9982, 49.51987, 10.05844, 0.003400783, 0, 
    0.6139406, 3.471415, 65.67765, 299.1868, 664.0464, 680.472, 861.0681, 
    1173.805, 1176.411, 882.2818, 935.2615, 1119.443, 1414.621, 875.902, 
    96.9949, 90.53958, 68.45934, 107.9565, 151.2383, 211.1697, 253.7371, 
    301.2069, 273.2981, 195.7737, 154.6178, 177.9713, 194.5825, 716.4048, 
    1805.13, 2597.123, 3127.537, 3920.587, 4658.365, 4768.674, 4483.495, 
    4462.699, 4175.957, 3900.408, 2836.106, 1404.504, 405.8325, 765.2993, 
    1341.417, 1822.338, 2584.409, 2872.491, 2385.164, 1991.338, 2122.929, 
    2156.027, 1849.882, 1308.424, 1070.509, 911.2019, 667.9567, 410.6019, 
    468.2829, 439.6035, 464.8657, 421.4958, 294.738, 311.5735, 259.9264, 
    141.5647, 14.46012, 0, 0, 0, 196.0959, 1.784637, 0, 0, 0, 0,
  589.6921, 369.2813, 29.13641, 0, 10.16494, 462.0075, 953.4734, 992.8953, 
    961.825, 980.4223, 959.9498, 878.5264, 782.0342, 714.8068, 590.7191, 
    438.146, 255.681, 89.16268, 4.204259, 2.031146, 0, 103.8879, 350.6954, 
    283.9107, 257.0193, 369.5965, 704.6323, 645.6995, 1036.557, 1464.105, 
    1060.085, 778.238, 741.6763, 1037.683, 1462.557, 1146.481, 278.6887, 
    344.5007, 247.6657, 85.39928, 122.3622, 162.2269, 193.9326, 217.9708, 
    211.0545, 208.4449, 336.8265, 831.7836, 1583.831, 2516.133, 3871.765, 
    4676.438, 4954.179, 5109.451, 5170.38, 4871.32, 4830.958, 4825.001, 
    4712.904, 4750.763, 4316.47, 2986.506, 1810.279, 1907.389, 3094.098, 
    3158.578, 3400.082, 3428.866, 3037.146, 2417.081, 2381.95, 2137.81, 
    1823.436, 1536.647, 1236.298, 1032.425, 829.5073, 612.1199, 627.1792, 
    549.0421, 514.0405, 437.2412, 523.9689, 332.4905, 376.6574, 324.6547, 
    278.9478, 18.89644, 0.006937383, 11.19048, 622.1964, 266.2146, 0, 0, 0, 0,
  418.7992, 35.6242, 0, 0.003005615, 134.9476, 670.2584, 953.2305, 938.2223, 
    913.4232, 907.8433, 847.9294, 775.7874, 707.1496, 637.6665, 506.9577, 
    328.1991, 144.9271, 21.72296, 0.001061579, 0, 193.2861, 655.1348, 
    890.2563, 1015.931, 1077.46, 1348.436, 1022.688, 766.3108, 1302.777, 
    1343.477, 1030.237, 887.298, 1036.799, 1030.548, 1415.412, 1369.234, 
    954.7562, 897.3719, 604.0056, 161.5459, 117.0032, 160.0316, 186.1864, 
    199.844, 234.4324, 490.8765, 1452.577, 2787.096, 3704.978, 4565.677, 
    5041.605, 5282.9, 5283.827, 5293.211, 5223.339, 5147.862, 5045.44, 
    5014.276, 4810.225, 4833.973, 4828.4, 4279.334, 3368.46, 3630.062, 
    4304.909, 4239.586, 3954.809, 3997.183, 3638.99, 3208.818, 2409.19, 
    1711.776, 1245.757, 1107.457, 1129.331, 956.4644, 789.5651, 568.699, 
    588.8917, 465.5713, 293.4032, 391.9729, 524.9534, 425.9501, 367.7643, 
    501.6449, 504.5149, 232.682, 5.703031, 0.4608422, 517.0116, 853.5552, 0, 
    0, 0, 0,
  208.9919, 0.07399444, 0, 86.20094, 452.0786, 852.0658, 1002.409, 962.3193, 
    888.443, 812.5153, 720.5767, 644.718, 631.5153, 512.2603, 381.4651, 
    213.2256, 41.59562, 0.2816853, 0, 124.2844, 722.3979, 1113.143, 1471.473, 
    1611.769, 2112.062, 2108.031, 1182.046, 772.6594, 1133.844, 1030.302, 
    594.0649, 781.9883, 976.3713, 996.936, 1344.194, 1913.446, 1758.966, 
    1584.213, 828.5089, 218.7474, 120.6228, 168.4115, 186.3442, 204.9695, 
    454.7095, 1957.652, 3490.757, 4445.193, 5092.852, 5200.075, 5270.465, 
    5072.342, 5013.149, 4973.931, 4979.826, 5028.506, 4968.484, 5000.479, 
    4901.846, 4918.038, 5056.896, 4726.156, 4305.746, 4395.774, 4665.846, 
    4441.66, 4191.952, 4342.861, 4170.3, 3571.407, 2256.272, 978.5087, 
    515.0765, 648.3031, 832.2507, 1023.514, 805.8867, 528.6307, 476.446, 
    414.0162, 249.9183, 179.4859, 455.012, 263.6515, 333.0435, 479.9664, 
    632.377, 499.215, 167.3804, 1.14105, 187.7418, 1096.691, 4.065651, 0, 0, 0,
  217.0772, 0.0330215, 14.08818, 507.184, 689.6525, 956.0153, 1135.08, 
    1068.822, 935.9532, 833.0918, 700.9478, 584.4554, 511.998, 405.4882, 
    298.7473, 151.3782, 10.5746, 0, 13.38639, 627.0316, 1415.375, 1796.191, 
    1776.488, 2020.439, 2216.457, 1986.079, 824.9573, 609.1418, 1088.619, 
    704.4744, 531.5552, 655.2637, 836.7814, 991.5665, 1400.434, 1907.079, 
    2138.898, 1730.733, 856.8054, 192.3337, 187.5201, 182.8071, 191.2734, 
    306.0225, 1638.453, 3471.865, 4649.002, 5009.791, 4932.093, 5040.752, 
    4961.458, 4920.357, 4891.655, 4887.036, 4862.397, 4830.989, 4769.84, 
    4764.334, 4749.213, 4840.669, 4871.838, 4824.714, 4635.75, 4551.147, 
    4447.096, 4367.069, 4249.624, 4367.218, 4152.088, 3556.254, 2167.627, 
    517.2781, 330.44, 333.8921, 615.7012, 814.1959, 880.6069, 573.7075, 
    426.0545, 368.3916, 209.4412, 130.0882, 280.0025, 206.5527, 246.2915, 
    389.107, 555.9575, 505.8926, 402.7588, 39.14849, 0.2409696, 211.2308, 
    10.10999, 0.2490215, 8.65174, 0.6303881,
  32.38083, 0, 51.82127, 560.3418, 760.4517, 1012.509, 1175.754, 1092.682, 
    990.1829, 844.8569, 664.1961, 527.9617, 436.3003, 353.342, 264.007, 
    111.6445, 0.1420982, 0, 120.9445, 1149.31, 1999.209, 1945.943, 1973.386, 
    1762.449, 1950.817, 1315.04, 577.0366, 879.3376, 1191.386, 623.9373, 
    548.0479, 722.4045, 1082.094, 1262.284, 1544.662, 2178.558, 2164.37, 
    1978.036, 1035.92, 460.3963, 275.0108, 282.9265, 595.8168, 1425.515, 
    3292.09, 4695.376, 5096.314, 4968.224, 4930.162, 4852.206, 4795.105, 
    4827.783, 4907.193, 5035.4, 4982.63, 5017.723, 4947.738, 4862.034, 
    4921.563, 4884.641, 4879.072, 4878.018, 4793.002, 4559.51, 4386.215, 
    4295.125, 4247.954, 4282.634, 4102.235, 3924.184, 2823.693, 1224.186, 
    358.0084, 332.7956, 348.9137, 678.3985, 848.0242, 821.4729, 618.2599, 
    296.2792, 78.22495, 69.06935, 236.8286, 218.569, 131.588, 226.8546, 
    405.3286, 521.6719, 575.6138, 185.445, 0.1386309, 0, 0.01035178, 0, 0, 
    0.3566946,
  0, 3.552063, 321.7133, 849.3109, 976.9869, 1078, 1041.034, 971.9257, 
    896.7177, 738.8071, 609.843, 479.6385, 370.4907, 299.6009, 196.0335, 
    43.93956, 1.847782, 58.31754, 820.1542, 1913.927, 2158.314, 2047.404, 
    1703.193, 1653.195, 1413.601, 1037.866, 736.9638, 1415.212, 1414.237, 
    810.8496, 802.1318, 1344.746, 1755.177, 1950.15, 2215.817, 2564.552, 
    2719.364, 2259.201, 1462.947, 672.4842, 476.5094, 949.2522, 1674.35, 
    3053.793, 4114.063, 4946.655, 5076.482, 5097.934, 5060.518, 5084.558, 
    5115.013, 5053.414, 5074.056, 5093.611, 5064.592, 5146.818, 5095.178, 
    5143.528, 5132.971, 5072.526, 4904.224, 4783.976, 4806.5, 4586.318, 
    4403.593, 4429.247, 4359.3, 4282.01, 4076.977, 3919.891, 3721.054, 
    2170.56, 812.0792, 348.9857, 379.0044, 509.2384, 835.6813, 1042.576, 
    981.3938, 473.188, 59.4187, 54.51209, 257.2173, 304.478, 147.0937, 
    83.89629, 318.8223, 480.2112, 706.43, 507.7156, 43.1609, 0, 0, 0, 
    0.06568222, 0,
  0, 74.23603, 787.8488, 1047.875, 1021.896, 987.5112, 943.1434, 865.201, 
    751.0483, 636.3491, 527.4158, 403.2906, 282.5342, 179.8925, 87.43723, 
    3.748239, 13.04159, 420.638, 1624.73, 2216.099, 2128.865, 1733.536, 
    1583.128, 1268.357, 1247.077, 910.689, 1149.7, 1639.568, 1381.821, 
    977.155, 1235.957, 1915.405, 2513.842, 2519.291, 2726.454, 3145.376, 
    2913.469, 2521.798, 1770.634, 1137.481, 1062.631, 1737.886, 2865.038, 
    3579.866, 4525.335, 4868.795, 5310.432, 5363.74, 5347.537, 5387.418, 
    5274.167, 5170.409, 5133.905, 5203.841, 5101.455, 5070.62, 5106.412, 
    5089.334, 5089.588, 4879.959, 4693.276, 4713.932, 4758.439, 4678.091, 
    4520.184, 4536.472, 4453.167, 4362.481, 4144.474, 3822.403, 3798.529, 
    3049.53, 1477.426, 703.8835, 612.568, 658.7606, 819.6526, 1062.141, 
    1055.71, 575.3791, 73.42055, 27.57079, 103.5562, 207.4734, 120.4412, 
    30.39635, 148.8998, 383.1422, 591.7628, 532.1869, 174.8339, 1.234607, 0, 
    0, 0, 0,
  6.758009, 487.5991, 1021.831, 1115.679, 886.489, 892.4991, 847.3696, 
    758.7397, 623.5787, 508.0063, 426.4549, 305.7114, 158.1539, 48.50787, 
    5.502139, 5.127207, 40.45427, 1082.158, 2018.84, 2095.057, 1691.412, 
    1381.58, 1191.657, 1015.282, 1019.028, 1079.314, 1296.271, 1340.825, 
    1178.45, 832.3215, 1319.656, 1844.028, 2394.739, 2776.184, 3035.285, 
    3199.43, 3069.708, 2704.726, 3048.322, 2788.972, 2680.07, 3130.915, 
    3342.005, 4203.668, 4655.496, 5272.828, 5415.704, 5200.595, 5129.409, 
    5031.954, 5205.507, 5085.389, 5081.525, 5094.905, 5042.618, 5019.026, 
    4992.753, 5047.111, 5006.662, 4865.849, 4714.873, 4635.37, 4685.44, 
    4620.996, 4597.202, 4502.657, 4462.631, 4332.861, 4098.364, 3766.416, 
    3657.072, 3297.008, 2097.184, 1253.378, 1089.461, 1061.64, 1174.932, 
    1281.606, 1266.194, 835.1642, 263.9403, 79.5519, 32.27344, 68.0872, 
    131.0868, 118.724, 164.2968, 321.6274, 409.3891, 379.2769, 350.8774, 
    57.88399, 0.000805264, 0, 0, 0,
  238.1623, 791.4998, 1109.681, 899.7229, 803.0744, 786.03, 737.5471, 
    634.7917, 498.6732, 393.5605, 324.9799, 180.8011, 45.09904, 5.052932, 
    12.10084, 59.62862, 665.7957, 1742.159, 2304.37, 1936.526, 1518.453, 
    1209.02, 957.4006, 869.3815, 823.4235, 999.6229, 1120.257, 1287.387, 
    1058.116, 943.8759, 842.4662, 1182.286, 1637.921, 2097.368, 2345.563, 
    2374.775, 1990.883, 2252.895, 3334.049, 3940.562, 4061.273, 4010.166, 
    4178.608, 4529.894, 4820.277, 4816.019, 4359.409, 3582.755, 3025.995, 
    3098.254, 3615.333, 4245.46, 4695.494, 5053.856, 5057.838, 5040.737, 
    4995.706, 4951.887, 5012.489, 4828.667, 4652.396, 4480.73, 4422.274, 
    4482.873, 4418.603, 4365.641, 4435.617, 4158.283, 3927.431, 3744.359, 
    3460.329, 3134.216, 2236.319, 1473.672, 1232.209, 1085.229, 938.4994, 
    930.7794, 780.1253, 518.0501, 171.889, 131.0825, 128.4954, 145.3723, 
    306.1799, 273.0995, 216.7841, 302.7602, 352.1556, 292.1012, 300.0482, 
    151.9467, 1.769033, 0, 0, 0,
  762.3385, 958.6488, 967.5426, 836.1221, 672.2523, 743.9036, 705.8074, 
    585.7993, 412.0986, 315.1353, 220.0953, 76.00178, 7.931051, 19.07306, 
    352.5095, 807.7217, 1467.913, 2206.177, 2116.3, 1479.32, 1129.964, 
    788.2949, 807.8799, 715.9404, 766.021, 992.697, 1301.655, 1434.707, 
    1353.936, 786.4489, 618.7448, 572.2695, 753.1136, 781.6061, 869.8459, 
    807.5753, 789.2447, 793.95, 2282.462, 3481.706, 4177.188, 4562.651, 
    4439.226, 4581.507, 3711.448, 2810.206, 2234.735, 1677.431, 1388.387, 
    1278.489, 1672.559, 2128.335, 3001.532, 3830.48, 4550.405, 4801.908, 
    4633.007, 4499.204, 4535.861, 4201.199, 3729.332, 3460.189, 3439.621, 
    3560.627, 3621.553, 3831.16, 4091.066, 3848.02, 3584.761, 3534.397, 
    3254.213, 2773.562, 2217.112, 1683.945, 1579.851, 1373.786, 1237.948, 
    1035.855, 892.402, 538.7142, 249.4172, 148.4552, 154.6931, 130.894, 
    219.8244, 191.3214, 59.69934, 129.1412, 212.872, 166.6351, 130.7894, 
    118.5202, 14.56528, 0, 0, 0,
  989.5663, 927.1322, 930.0528, 724.9628, 672.3023, 786.1067, 760.7014, 
    580.4506, 387.8854, 255.2157, 132.3959, 20.43845, 25.85789, 478.4587, 
    1034.186, 1562.984, 1919.749, 2048.771, 1455.002, 993.2492, 1055.018, 
    1015.837, 1037.239, 1008.556, 891.994, 1129.969, 1403.661, 1486.652, 
    921.8677, 453.2355, 336.5799, 424.1663, 397.4917, 279.882, 307.3911, 
    629.627, 392.5599, 732.6076, 1854.792, 3292.929, 4316.049, 4438.208, 
    4466.581, 3936.618, 2551.772, 1529.796, 1225.804, 1185.416, 1170.846, 
    1186.658, 1149.756, 1173.267, 1364.58, 2012.139, 2864.934, 3708.189, 
    4220.437, 4108.575, 3883.59, 3378.89, 2934.686, 2709.543, 2824.293, 
    3108.43, 3076.333, 3295.794, 3656.051, 3385.662, 3217.673, 3000.589, 
    2639.363, 2225.868, 2004.855, 1872.814, 1614.911, 1220.716, 921.0709, 
    856.4285, 921.3516, 950.4296, 616.0353, 308.2891, 110.1128, 48.46398, 
    55.95203, 45.66961, 26.53019, 25.74332, 58.75687, 44.34055, 7.046542, 
    9.698866, 7.823508, 0.1154567, 0, 0,
  873.5029, 932.446, 802.8636, 679.261, 728.6178, 853.7338, 757.9206, 
    581.5193, 393.3805, 206.899, 67.25694, 23.86274, 177.6185, 981.5392, 
    1598.842, 1796.156, 1947.744, 1703.935, 1375.229, 1515.294, 1642.378, 
    1676.018, 1487.45, 1227.913, 1159.733, 1323.913, 1554.071, 1138.957, 
    556.8956, 169.3183, 218.1516, 265.9337, 235.5797, 302.2885, 690.3524, 
    1159.933, 1460.098, 1501.492, 2359.936, 3452.56, 4296.354, 4520.364, 
    4153.528, 3140.282, 1694.784, 1188.321, 1116.658, 1141.684, 1149.989, 
    1137.289, 1126.685, 1111.867, 1065.968, 976.756, 1235.389, 1905.175, 
    2724.575, 3200.128, 3303.74, 2937.104, 2721.535, 2951.062, 3359.012, 
    3876.756, 3978.864, 3924.08, 3884.962, 3585.292, 3361.129, 3095.249, 
    2504.762, 2074.735, 1898.636, 1876.1, 1742.129, 1328.015, 1136.963, 
    851.3479, 765.448, 628.5696, 611.1027, 228.0393, 106.5588, 40.51612, 
    28.73609, 26.4498, 39.7077, 42.63209, 21.35075, 11.05065, 3.122396, 
    2.336835, 0.5792097, 0.1638553, 0, 0,
  546.0862, 803.7518, 720.4936, 680.9647, 811.3162, 854.0582, 728.9124, 
    554.4362, 350.1646, 161.0941, 51.3675, 48.73245, 369.3617, 1295.04, 
    1821.616, 1891.482, 1897.59, 1783.333, 1780.204, 1693.617, 841.7841, 
    444.8978, 635.6622, 896.0977, 1128.595, 1378.011, 996.2464, 523.0845, 
    123.556, 142.2115, 182.9801, 192.1028, 208.9994, 239.5104, 673.2095, 
    1674.933, 2271.34, 2666.304, 2851.325, 3098.809, 3555.89, 3740.312, 
    3572.558, 2706.249, 1709.02, 1359.368, 1286.218, 1109.896, 1039.783, 
    1053.64, 1038.432, 1022.949, 1007.573, 974.9078, 853.291, 834.8326, 
    1136.756, 1648.817, 2111.175, 2467.282, 2775.722, 3019.613, 3544.646, 
    4111.462, 4240.049, 4245.177, 4150.613, 3692.481, 3492.051, 3113.697, 
    2519.094, 1983.502, 1739.186, 1723.87, 1627.539, 1467.329, 1415.479, 
    1188.471, 862.6572, 819.2594, 613.4723, 440.3748, 103.548, 44.31029, 
    44.08937, 32.32762, 27.8348, 27.06621, 14.8008, 2.686884, 3.042891, 
    2.475014, 0.1258945, 0, 0, 0,
  287.7358, 699.6454, 753.7252, 715.9815, 790.1022, 770.7126, 621.1946, 
    429.5545, 302.6275, 146.0066, 109.7574, 238.4723, 702.8896, 1500.438, 
    1914.869, 1864.13, 1797.373, 1384.315, 1103.181, 50.18019, -29, 
    -28.77262, 25.38564, 296.886, 687.7216, 647.961, 349.3248, 83.32568, 
    112.7014, 157.216, 171.5177, 178.561, 204.0525, 312.3961, 523.767, 
    829.8365, 1039.718, 1047.279, 1355.524, 1172.16, 1411.563, 2336.885, 
    3058.305, 3226.443, 3063.086, 2861.304, 2247.198, 1404.461, 1073.007, 
    987.9013, 956.4599, 926.052, 903.3677, 896.808, 893.4102, 892.0126, 
    796.2086, 820.1337, 984.0677, 1229.673, 1469.496, 1966.5, 2469.902, 
    3181.495, 3622.321, 3652.744, 3231.653, 2652.689, 2285.655, 2040.421, 
    1670.866, 1479.306, 1414.353, 1424.594, 1447.813, 1503.411, 1473.374, 
    1250.532, 1041.187, 973.3618, 1039.013, 789.7152, 424.5931, 71.7645, 
    43.34607, 37.34945, 45.60085, 23.38318, 6.514248, 1.005424, 1.192295, 
    0.07372784, 0, 0, 0, 0,
  280.0255, 717.2288, 800.9051, 767.515, 678.3198, 625.6271, 422.783, 
    283.5512, 241.4006, 186.5598, 174.9805, 521.5108, 1183.758, 1658.958, 
    2034.699, 1761.583, 1296.187, 204.5876, -27.33, -29, -29, -28.70372, 
    31.97342, 167.3994, 247.8943, 170.875, 60.56211, 102.6041, 146.6671, 
    170.812, 176.8664, 183.8537, 244.3707, 366.5971, 502.9418, 470.5995, 
    290.3222, 581.1486, 1270.705, 1402.007, 1254.245, 1784.784, 2600.036, 
    2944.01, 3219.255, 3399.147, 3218.488, 2378.177, 1818.334, 1375.318, 
    1074.772, 1071.595, 984.6507, 961.2864, 971.7458, 1197.327, 1193.799, 
    1028.109, 963.4049, 965.5383, 1135.214, 1159.892, 1419.062, 1704.113, 
    1884.114, 1810.738, 1669.92, 1423.683, 1450.932, 1501.812, 1357.503, 
    1354.311, 1357.144, 1350.14, 1337.69, 1373.946, 1390.578, 1208.278, 
    1047.752, 1206.215, 1150.309, 1096.129, 627.1903, 92.17794, 38.86603, 
    55.03728, 97.46461, 80.68608, 19.16875, 1.530113, 0.02449018, 0, 0, 0, 0, 0,
  278.7002, 848.4108, 836.0483, 703.4719, 592.2507, 425.2289, 267.3521, 
    212.9088, 260.6262, 199.7883, 384.8431, 1051.43, 1458.136, 1718.665, 
    1860.108, 1682.248, 920.7298, -29, -29, -29, -29, -26.10924, 98.29451, 
    120.4517, 76.57224, 60.59356, 87.99368, 121.3795, 137.9679, 144.398, 
    164.9114, 216.217, 274.5612, 275.6122, 318.0442, 259.2065, 230.8655, 
    623.9655, 1918.901, 2278.465, 2228.787, 2412.379, 2568.84, 2575.392, 
    2590.898, 2936.103, 3116.961, 3308.007, 3364.986, 2819.327, 2346.359, 
    2102.324, 1968.311, 1727.268, 1581.183, 1342.206, 1030.278, 1016.645, 
    1021.907, 1084.763, 1044.676, 1257.469, 1468.743, 1774.683, 1740.715, 
    1517.49, 1302.269, 1243.797, 1198.531, 1266.439, 1397.631, 1400.947, 
    1359.057, 1343.482, 1246.818, 1367.203, 1329.797, 1222.678, 1103.928, 
    1230.625, 1299.724, 1154.313, 827.8479, 142.0308, 30.594, 63.95813, 
    176.8368, 209.5096, 94.29587, 2.645784, 0, 0, 0, 0, 0, 0,
  372.7461, 1182.848, 984.7722, 758.8289, 559.1176, 423.6849, 319.4374, 
    300.4261, 340.6555, 502.4338, 1127.504, 1562.021, 1634.167, 1688.647, 
    1848.811, 1538.005, 454.8116, -28.99981, -29, -29, -27.34004, 37.3294, 
    157.3012, 172.0072, 120.2076, 77.74836, 81.51273, 100.2689, 110.1352, 
    113.6465, 112.3892, 174.2308, 265.0841, 238.038, 208.7626, 195.9964, 
    185.5608, 428.3402, 1028.99, 1427.11, 1409.885, 1349.094, 1442.432, 
    1663.696, 1924.178, 2039.838, 2233.458, 2097.392, 2286.286, 2274.246, 
    2335.328, 2740.635, 3043.788, 3113.309, 2620.314, 1823.444, 907.4882, 
    560.1979, 721.8196, 618.8461, 714.8278, 968.9215, 1536.432, 1776.954, 
    1845.922, 1518.606, 1331.444, 1091.121, 1037.558, 1111.581, 1316.298, 
    1388.658, 1346.563, 1293.286, 1239.811, 1305.997, 1406.889, 1326.371, 
    1211.889, 1292.238, 1407.659, 1205.926, 807.7815, 109.0812, 17.7631, 
    51.74597, 188.0972, 276.9687, 185.2122, 45.17762, 0, 0, 0, 0, 0, 0,
  23.64984, 599.7591, 511.6504, 444.8416, 378.2097, 360.2961, 380.9373, 
    438.2814, 595.3414, 1348.148, 2057.229, 2197.964, 1472.968, 1671.91, 
    1237.43, 761.7867, 28.29826, -28.70648, -28.99438, -29, -24.99033, 
    18.25178, 63.3651, 174.8866, 123.8744, 57.97906, 65.55949, 76.69518, 
    97.68421, 102.3149, 131.3378, 195.444, 256.4067, 243.5822, 187.5729, 
    165.1665, 342.9257, 405.3759, 560.9412, 516.8105, 509.3314, 621.6459, 
    699.2636, 746.7856, 760.3452, 922.6527, 823.6852, 1078.508, 1096.203, 
    1233.275, 1588.237, 2370.672, 2694.676, 2629.588, 2156.679, 1783.274, 
    1690.359, 1606.746, 1283.696, 1141.156, 1217.001, 1620.093, 1467.414, 
    1503.383, 1485.695, 1331.391, 1196.225, 1032.619, 951.8022, 972.683, 
    1066.139, 1124.131, 1171.412, 1188.777, 1279.054, 1209.068, 1229.401, 
    1345.554, 1244.472, 1249.917, 1464.447, 1206.628, 878.3694, 171.7012, 
    12.43563, 7.429965, 32.89956, 78.383, 51.98663, 29.90217, 24.32074, 0, 0, 
    0, 0, 0,
  1.67216, 340.6524, 385.0545, 416.1772, 390.3365, 441.3774, 650.9087, 
    704.9575, 1160.624, 1782.02, 2326.5, 2033.687, 1439.484, 1619.828, 
    746.22, 75.66013, 201.0358, 17.39066, -28.43431, -29, -27.93392, 
    -29.96976, 155.6212, 198.6232, 113.8873, 86.04948, 76.57941, 72.31518, 
    72.27863, 74.17043, 85.37265, 140.0728, 171.7061, 157.3423, 148.0897, 
    287.3974, 366.4878, 442.8387, 367.5465, 295.4169, 339.7092, 412.319, 
    477.4836, 479.2714, 430.4697, 594.4115, 1253.493, 1810.096, 2104.204, 
    1634.684, 1001.775, 974.5079, 900.9539, 634.2441, 554.7181, 615.168, 
    911.0193, 996.5089, 1222.358, 1436.428, 1665.35, 1462.017, 1208.923, 
    960.894, 1190.559, 1318.656, 1208.269, 1155.516, 1205.878, 1180.793, 
    1165.779, 1183.944, 1099.437, 1158.785, 1276.583, 1278.646, 1152.482, 
    1210.833, 1241.654, 1143.037, 1397.42, 1334.603, 1178.972, 665.2888, 
    53.88091, 2.508959, 0.1916037, 1.167866, 4.74597, 36.34115, 73.30758, 
    20.18326, 0, 0, 0, 0.04834903 ;
}
