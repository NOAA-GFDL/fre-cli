netcdf frenctools_timavg_atmos.197901-198312.LWP {
dimensions:
	time = UNLIMITED ; // (1 currently)
	lat = 180 ;
	lon = 288 ;
	bnds = 2 ;
variables:
	float LWP(time, lat, lon) ;
		LWP:_FillValue = 1.e+20f ;
		LWP:missing_value = 1.e+20f ;
		LWP:units = "kg m-2" ;
		LWP:long_name = "Liquid Water Path" ;
		LWP:cell_measures = "area: area" ;
		LWP:standard_name = "atmosphere_mass_content_of_cloud_liquid_water" ;
		LWP:interp_method = "conserve_order2" ;
		LWP:cell_methods = "time: mean" ;
		LWP:time_avg_info = "average_T1,average_T2,average_DT" ;
	double bnds(bnds) ;
		bnds:long_name = "vertex number" ;
	double lat(lat) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_N" ;
		lat:axis = "Y" ;
		lat:bounds = "lat_bnds" ;
	double lat_bnds(lat, bnds) ;
		lat_bnds:long_name = "latitude bounds" ;
		lat_bnds:units = "degrees_N" ;
		lat_bnds:axis = "Y" ;
	double lon(lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_E" ;
		lon:axis = "X" ;
		lon:bounds = "lon_bnds" ;
	double lon_bnds(lon, bnds) ;
		lon_bnds:long_name = "longitude bounds" ;
		lon_bnds:units = "degrees_E" ;
		lon_bnds:axis = "X" ;
	double time(time) ;
		time:units = "days since 1979-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "JULIAN" ;
		time:calendar = "julian" ;
		time:bounds = "time_bnds" ;
	double time_bnds(time, bnds) ;
		time_bnds:units = "days since 1979-01-01 00:00:00" ;
		time_bnds:long_name = "time axis boundaries" ;
	double average_T1(time) ;
		average_T1:long_name = "Start time for average period" ;
		average_T1:units = "days since 1979-01-01 00:00:00" ;
	double average_T2(time) ;
		average_T2:long_name = "End time for average period" ;
		average_T2:units = "days since 1979-01-01 00:00:00" ;
	double average_DT(time) ;
		average_DT:long_name = "Length of average period" ;
		average_DT:units = "days" ;

// global attributes:
		:title = "c96L33_am5f1a0r0_amip" ;
		:associated_files = "area: 19830101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:code_release_version = "2022.02" ;
		:git_hash = "83acb799f47dfa27b433a131e9f7c1310767cc59" ;
		:creationtime = "Sat Feb 18 02:08:21 2023" ;
		:hostname = "pp022" ;
		:history = "fregrid --standard_dimension --input_mosaic C96_mosaic.nc --input_file 19830101.atmos_month --interp_method conserve_order2 --remap_file .fregrid_remap_file_288_by_180.nc --nlon 288 --nlat 180 --scalar_field (**please see the field list in this file**) --output_file out.nc" ;
		:external_variables = "area" ;
		:comment = "FMS time averaging, version 3.0, precision=double" ;
data:

 LWP =
  0.0008464053, 0.0008469686, 0.0008475319, 0.0008480952, 0.0008486585, 
    0.0008492218, 0.0008497852, 0.0008503484, 0.0008509118, 0.0008514751, 
    0.0008520384, 0.0008526017, 0.000853165, 0.0008537283, 0.0008542916, 
    0.0008548549, 0.0008554182, 0.0008559815, 0.0008565448, 0.0008571081, 
    0.0008576714, 0.0008582347, 0.000858798, 0.0008593613, 0.0008599247, 
    0.0008604879, 0.0008610513, 0.0008616145, 0.0008621779, 0.0008627411, 
    0.0008633045, 0.0008638678, 0.0008644311, 0.0008649944, 0.0008655577, 
    0.000866121, 0.0008666843, 0.0008672476, 0.0008678109, 0.0008683742, 
    0.0008689375, 0.0008695009, 0.0008700641, 0.0008706275, 0.0008711907, 
    0.0008717541, 0.0008723174, 0.0008728807, 0.000873444, 0.0008740073, 
    0.0008745706, 0.0008751339, 0.0008756972, 0.0008762605, 0.0008768238, 
    0.0008773871, 0.0008779504, 0.0008785137, 0.000879077, 0.0008796403, 
    0.0008802036, 0.000880767, 0.0008813302, 0.0008818936, 0.0006399711, 
    0.0006408087, 0.0006416464, 0.0006424841, 0.0006433217, 0.0006441594, 
    0.000644997, 0.0006458347, 0.0006466723, 0.00064751, 0.0006483477, 
    0.0006491853, 0.000650023, 0.0006508607, 0.0006516983, 0.000652536, 
    0.0006533737, 0.0006542113, 0.000655049, 0.0006558867, 0.0006567243, 
    0.000657562, 0.0006583997, 0.0006592373, 0.0006600749, 0.0006609126, 
    0.0006617503, 0.0006625879, 0.0006634256, 0.0006642633, 0.0006651009, 
    0.0006659386, 0.0006667763, 0.0006676139, 0.0006684516, 0.0006692893, 
    0.0006701269, 0.0006709646, 0.0006718023, 0.0006726399, 0.0006734776, 
    0.0006743153, 0.0006751529, 0.0006759905, 0.0006768282, 0.0006776659, 
    0.0006785035, 0.0006793412, 0.0006801789, 0.0006810165, 0.0006818542, 
    0.0006826919, 0.0006835295, 0.0006843672, 0.0006852049, 0.0006860425, 
    0.0006868802, 0.0006877179, 0.0006885555, 0.0006893931, 0.0006902309, 
    0.0006910685, 0.0006919061, 0.0006927438, 0.0006935815, 0.0006944191, 
    0.0006952568, 0.0006960945, 0.0006969321, 0.0006977698, 0.0006986075, 
    0.0006994451, 0.0008707179, 0.0008701738, 0.0008696297, 0.0008690857, 
    0.0008685415, 0.0008679975, 0.0008674534, 0.0008669093, 0.0008663653, 
    0.0008658212, 0.0008652771, 0.0008647331, 0.000864189, 0.0008636449, 
    0.0008631009, 0.0008625567, 0.0008620127, 0.0008614686, 0.0008609245, 
    0.0008603805, 0.0008598364, 0.0008592923, 0.0008587482, 0.0008582042, 
    0.0008576601, 0.000857116, 0.0008565719, 0.0008560279, 0.0008554838, 
    0.0008549397, 0.0008543957, 0.0008538516, 0.0008533075, 0.0008527634, 
    0.0008522194, 0.0008516753, 0.0008511312, 0.0008505872, 0.0008500431, 
    0.000849499, 0.000848955, 0.0008484108, 0.0008478668, 0.0008473227, 
    0.0008467786, 0.0008462346, 0.0008456905, 0.0008451464, 0.0008446024, 
    0.0008440583, 0.0008435142, 0.0008429701, 0.0008424261, 0.000841882, 
    0.0008413379, 0.0008407938, 0.0008402498, 0.0008397057, 0.0008391616, 
    0.0008386176, 0.0008380734, 0.0008375294, 0.0008369853, 0.0008364412, 
    0.0008358972, 0.0008353531, 0.000834809, 0.000834265, 0.0008337209, 
    0.0008331768, 0.0008326327, 0.0008320886, 0.0007604815, 0.0007596246, 
    0.0007587677, 0.0007579108, 0.0007570539, 0.000756197, 0.0007553402, 
    0.0007544832, 0.0007536263, 0.0007527695, 0.0007519125, 0.0007510557, 
    0.0007501988, 0.0007493419, 0.000748485, 0.0007476281, 0.0007467712, 
    0.0007459143, 0.0007450574, 0.0007442005, 0.0007433436, 0.0007424867, 
    0.0007416298, 0.0007407729, 0.000739916, 0.0007390591, 0.0007382022, 
    0.0007373453, 0.0007364884, 0.0007356316, 0.0007347746, 0.0007339178, 
    0.0007330609, 0.0007322039, 0.0007313471, 0.0007304902, 0.0007296333, 
    0.0007287764, 0.0007279195, 0.0007270626, 0.0007262057, 0.0007253488, 
    0.0007244919, 0.000723635, 0.0007227781, 0.0007219212, 0.0007210643, 
    0.0007202074, 0.0007193505, 0.0007184937, 0.0007176367, 0.0007167798, 
    0.000715923, 0.000715066, 0.0007142092, 0.0007133523, 0.0007124954, 
    0.0007116385, 0.0007107815, 0.0007099247, 0.0007090678, 0.0007082109, 
    0.000707354, 0.0007064971, 0.0007056402, 0.0007047833, 0.0007039264, 
    0.0007030695, 0.0007022126, 0.0007013557, 0.0007004988, 0.0006996419, 
    0.0008418988, 0.0008424622, 0.0008430255, 0.0008435888, 0.0008441521, 
    0.0008447154, 0.0008452787, 0.000845842,
  0.0005935117, 0.0005964308, 0.0005993841, 0.0006023719, 0.0006053949, 
    0.0006084533, 0.0006115477, 0.0006146784, 0.0006178459, 0.0006210506, 
    0.000624293, 0.0006275736, 0.0006308928, 0.000634251, 0.0006376488, 
    0.0006410866, 0.0006445649, 0.0006480843, 0.0006518835, 0.0006655287, 
    0.0006841312, 0.0007026145, 0.0007209495, 0.0007391091, 0.0007570683, 
    0.0007748037, 0.0007922939, 0.0008095191, 0.0008243831, 0.0008372021, 
    0.0008499718, 0.0008626513, 0.0008751972, 0.0008875636, 0.0008997022, 
    0.000911562, 0.0009230893, 0.0009310981, 0.0009326913, 0.00093411, 
    0.0009355071, 0.000936883, 0.0009382382, 0.0009395731, 0.0009408881, 
    0.0009421837, 0.0009434601, 0.0009447178, 0.0009459573, 0.0009471789, 
    0.0009483829, 0.0009495698, 0.00095074, 0.0009518936, 0.0009530311, 
    0.0009541529, 0.0009552593, 0.0009563506, 0.0009574271, 0.0009584892, 
    0.0009595371, 0.0009605712, 0.0009615918, 0.0009625991, 0.0007830141, 
    0.0007820014, 0.0007809906, 0.0007799825, 0.0007789776, 0.0007779765, 
    0.0007769799, 0.0007759883, 0.0007750025, 0.0007740229, 0.0007730504, 
    0.0007720856, 0.0007711293, 0.0007701819, 0.0007692444, 0.0007683175, 
    0.0007674019, 0.0007664983, 0.0007656076, 0.0007647305, 0.0007638679, 
    0.0007630204, 0.0007621891, 0.0007613747, 0.000760578, 0.0007598001, 
    0.0007592207, 0.0007660254, 0.00077667, 0.0007873228, 0.0007979605, 
    0.0008085607, 0.0008191019, 0.0008295631, 0.0008399246, 0.0008501671, 
    0.0008531811, 0.0008491246, 0.000845145, 0.0008412751, 0.0008375495, 
    0.0008340043, 0.0008306779, 0.0008276099, 0.0008248422, 0.0008248918, 
    0.0008298726, 0.0008349849, 0.0008401101, 0.0008452472, 0.0008503954, 
    0.0008555535, 0.0008607209, 0.0008658966, 0.0008710797, 0.0008762694, 
    0.0008814649, 0.0008866653, 0.0008918699, 0.0008970779, 0.0009022885, 
    0.000907501, 0.0009127147, 0.0009179288, 0.0009231427, 0.0009283555, 
    0.0009335668, 0.0009387758, 0.0009439819, 0.0009491844, 0.0009543828, 
    0.0009595765, 0.0009079254, 0.0009202997, 0.0009325591, 0.0009446987, 
    0.0009567129, 0.0009685964, 0.0009803436, 0.0009919488, 0.001003406, 
    0.00101471, 0.001025855, 0.001036834, 0.001047641, 0.001058271, 
    0.001068716, 0.00107897, 0.001089026, 0.001098879, 0.00110852, 
    0.001117943, 0.001127141, 0.001136107, 0.001144833, 0.001153311, 
    0.001161535, 0.001169497, 0.001176414, 0.001149954, 0.001102752, 
    0.001050926, 0.0009949337, 0.0009352159, 0.000872197, 0.0008062858, 
    0.0007378756, 0.0006673446, 0.0006478619, 0.0006798829, 0.0007112487, 
    0.0007418395, 0.0007715375, 0.000800227, 0.0008277943, 0.0008541273, 
    0.0008791158, 0.0008922874, 0.0008853488, 0.0008778291, 0.0008702141, 
    0.0008625073, 0.0008547119, 0.0008468313, 0.0008388687, 0.0008308271, 
    0.0008227098, 0.0008145198, 0.00080626, 0.0007979335, 0.0007895433, 
    0.0007810919, 0.0007725825, 0.0007640176, 0.0007554001, 0.0007467325, 
    0.0007380176, 0.0007292578, 0.0007204557, 0.0007116138, 0.0007027346, 
    0.0006938204, 0.0006848736, 0.0006758965, 0.0009540125, 0.0009522258, 
    0.0009504207, 0.0009485969, 0.0009467541, 0.0009448918, 0.0009430098, 
    0.0009411075, 0.0009391846, 0.0009372407, 0.0009352753, 0.0009332881, 
    0.0009312786, 0.0009292464, 0.0009271909, 0.0009251119, 0.0009230088, 
    0.0009208812, 0.0009187285, 0.0009165503, 0.0009143462, 0.0009121154, 
    0.0009098577, 0.0009075725, 0.0009052592, 0.0009029172, 0.000900612, 
    0.0009009008, 0.0009023316, 0.0009034501, 0.0009042681, 0.0009047968, 
    0.0009050475, 0.0009050309, 0.0009047578, 0.0009042387, 0.0009058919, 
    0.0009094568, 0.000912352, 0.000914507, 0.0009158478, 0.0009162964, 
    0.0009157713, 0.0009141868, 0.0009114532, 0.0009078488, 0.0009042128, 
    0.000900499, 0.0008967011, 0.0008928212, 0.0008888619, 0.0008848254, 
    0.0008807137, 0.0008765293, 0.0008722742, 0.0008679503, 0.0008635599, 
    0.0008591049, 0.0008545873, 0.000850009, 0.0008453719, 0.0008406778, 
    0.0008359286, 0.000831126, 0.0008262718, 0.0008213675, 0.000816415, 
    0.0008114158, 0.0008063716, 0.0008012837, 0.0007961539, 0.0007909835, 
    0.0005713421, 0.000574002, 0.000576693, 0.0005794154, 0.0005821695, 
    0.0005849558, 0.0005877747, 0.0005906265,
  0.0005652407, 0.0005645728, 0.0005639278, 0.0005633062, 0.0005627084, 
    0.0005621349, 0.0005615863, 0.000561063, 0.0005611519, 0.0005686932, 
    0.0005780329, 0.000587085, 0.000595758, 0.0006064058, 0.0006230861, 
    0.0006399983, 0.000656881, 0.0006737118, 0.0006903165, 0.0007013443, 
    0.0007094978, 0.0007176432, 0.0007257817, 0.0007339145, 0.0007420433, 
    0.0007501696, 0.0007582954, 0.0007675958, 0.0007745961, 0.0007777499, 
    0.0007808883, 0.0007832882, 0.0007849817, 0.0007860003, 0.0007863747, 
    0.0007861355, 0.0007853124, 0.0007856719, 0.0007887359, 0.0007911242, 
    0.0007927195, 0.0007935065, 0.000794004, 0.0008042656, 0.0008178611, 
    0.0008302158, 0.0008410561, 0.0008477794, 0.0008456722, 0.0008428737, 
    0.0008400372, 0.0008371635, 0.0008342533, 0.0008313073, 0.0008283263, 
    0.0008253108, 0.0008222617, 0.0008191796, 0.0008160652, 0.0008129193, 
    0.0008097424, 0.0008065352, 0.0008032985, 0.0008000329, 0.000709517, 
    0.0007119436, 0.0007143482, 0.0007167305, 0.0007190899, 0.0007214259, 
    0.0007237383, 0.0007260264, 0.0007282899, 0.0007305283, 0.0007327411, 
    0.0007349278, 0.0007370881, 0.0007392213, 0.0007413271, 0.0007434048, 
    0.0007462511, 0.0007583924, 0.0007713739, 0.000782196, 0.0007910586, 
    0.0007994896, 0.0008104808, 0.0008217535, 0.0008331785, 0.0008447414, 
    0.000856322, 0.0008639341, 0.0008695367, 0.0008752599, 0.0008811072, 
    0.0008870816, 0.0008931864, 0.0008994251, 0.000905801, 0.0009105048, 
    0.0009048613, 0.0008960417, 0.000888193, 0.0008803257, 0.0008724483, 
    0.0008645687, 0.0008566949, 0.0008488346, 0.0008409951, 0.0008317804, 
    0.0008200108, 0.0008084141, 0.0007970952, 0.0007860903, 0.0007758887, 
    0.0007770586, 0.0007858297, 0.0007990806, 0.0008175448, 0.0008379202, 
    0.0008495018, 0.000860358, 0.0008713502, 0.0008824763, 0.0008937345, 
    0.0009051228, 0.0009166391, 0.0009282817, 0.0009400485, 0.0009519377, 
    0.0009639473, 0.0009760756, 0.0009883206, 0.00100068, 0.001013153, 
    0.001025737, 7.191663e-05, 0.0001725393, 0.0002720277, 0.000370362, 
    0.0004675223, 0.0005634884, 0.0006582401, 0.0007517571, 0.0008440187, 
    0.0009350044, 0.001024693, 0.001113065, 0.001200097, 0.00128577, 
    0.001370061, 0.00145295, 0.001556354, 0.001907864, 0.002267859, 
    0.002552141, 0.002769272, 0.002869814, 0.002797071, 0.002710855, 
    0.002618187, 0.002519338, 0.002415112, 0.002324664, 0.002240648, 
    0.002153556, 0.002063332, 0.001969923, 0.001873278, 0.001773343, 
    0.001670066, 0.001494822, 0.001405652, 0.001474305, 0.001500557, 
    0.001525169, 0.001548177, 0.001569618, 0.001589527, 0.001607941, 
    0.001624894, 0.001646566, 0.001678092, 0.001707733, 0.001735202, 
    0.001760465, 0.001781024, 0.00174375, 0.001674663, 0.001594718, 
    0.001502885, 0.001416853, 0.001387342, 0.001362209, 0.001336649, 
    0.001310667, 0.001284269, 0.001257462, 0.001230252, 0.001202644, 
    0.001174644, 0.00114626, 0.001117495, 0.001088357, 0.001058852, 
    0.001028984, 0.0009987593, 0.0009681844, 0.001004882, 0.0009886702, 
    0.0009727151, 0.0009570217, 0.0009415938, 0.000926436, 0.0009115525, 
    0.0008969477, 0.000882626, 0.0008685918, 0.0008548496, 0.0008414039, 
    0.0008282592, 0.0008154201, 0.0008028912, 0.000790677, 0.0007799043, 
    0.0007866093, 0.0008054079, 0.0008319451, 0.0008648641, 0.0008954498, 
    0.0009104729, 0.0009243184, 0.0009377067, 0.0009506285, 0.0009630416, 
    0.0009735313, 0.0009829171, 0.0009919811, 0.001000702, 0.001009058, 
    0.001017028, 0.001024589, 0.001031719, 0.001044034, 0.001054366, 
    0.001050339, 0.001046355, 0.001041412, 0.001035549, 0.001028808, 
    0.001021225, 0.001012841, 0.001003692, 0.0009936484, 0.000982206, 
    0.0009693257, 0.0009549686, 0.0009390996, 0.000921588, 0.0008994209, 
    0.0008742117, 0.0008475657, 0.0008194166, 0.0007935002, 0.0007806236, 
    0.000768809, 0.0007569934, 0.0007451768, 0.0007333595, 0.0007215416, 
    0.0007097232, 0.0006979044, 0.0006860855, 0.0006742664, 0.0006624475, 
    0.0006506287, 0.0006388102, 0.0006269922, 0.0006151748, 0.0006033581, 
    0.0005713507, 0.0005705167, 0.0005697018, 0.0005689066, 0.0005681315, 
    0.0005673768, 0.0005666431, 0.000565931,
  0.0005971921, 0.0005965328, 0.0005958689, 0.0005952003, 0.0006061077, 
    0.0006428891, 0.0006815103, 0.0006983414, 0.0007055616, 0.000708074, 
    0.0007093151, 0.0007107437, 0.0007123667, 0.0007141917, 0.000716226, 
    0.0007184771, 0.0007209526, 0.0007221487, 0.0007200317, 0.0007288835, 
    0.0007451973, 0.0007600521, 0.0007730866, 0.0007823199, 0.0007903286, 
    0.0007975965, 0.0008041738, 0.000809277, 0.0008115509, 0.0008115461, 
    0.00080991, 0.0008070949, 0.0008030265, 0.0007975218, 0.0007895874, 
    0.00077928, 0.0007665658, 0.0007597876, 0.000761128, 0.0007617528, 
    0.0007620311, 0.0007618566, 0.0007612411, 0.0007601966, 0.0007587348, 
    0.0007568671, 0.0007546049, 0.0007535693, 0.0007567821, 0.0007478959, 
    0.0007096871, 0.0006678398, 0.0006508621, 0.0006465212, 0.0006421756, 
    0.0006378255, 0.0006334707, 0.0006291114, 0.0006247477, 0.0006203796, 
    0.0006160072, 0.0006116306, 0.0006072496, 0.0006028646, 0.0006253003, 
    0.0006298897, 0.0006344469, 0.0006389715, 0.0006434632, 0.0006479218, 
    0.0006523469, 0.0006567381, 0.0006610951, 0.0006654176, 0.0006697052, 
    0.0006739576, 0.0006903739, 0.0007295973, 0.0007638924, 0.0007834752, 
    0.0007959916, 0.0008000178, 0.0008016148, 0.0008030281, 0.0008042532, 
    0.0008052853, 0.0008061198, 0.0008067521, 0.0008071773, 0.0008053334, 
    0.0007963371, 0.0007862223, 0.00077598, 0.0007654194, 0.0007551736, 
    0.0007482241, 0.000741529, 0.0007345643, 0.0007273681, 0.0007213031, 
    0.0007185962, 0.0007140489, 0.0007086279, 0.0007030756, 0.0006973975, 
    0.0006914639, 0.0006846559, 0.0006778188, 0.0006711468, 0.0006874749, 
    0.0007313244, 0.0007496424, 0.0007590171, 0.0007682868, 0.0007774504, 
    0.0007865073, 0.0007954565, 0.0008042975, 0.0008130294, 0.0008243996, 
    0.0008469872, 0.0008062881, 0.0006008397, 0.0004050635, 0.0003673699, 
    0.0004007418, 0.0004346547, 0.000469103, 0.0005040814, 0.0005395841, 
    0.0005756058, 0.0006121409, 0.0006491841, 0.0006867299, 0.0007247728, 
    0.0007633076, 0.0002077, 0.0004747724, 0.0007391731, 0.001000872, 
    0.00125984, 0.001516045, 0.001769459, 0.00202005, 0.002267789, 
    0.002512644, 0.002754585, 0.00299358, 0.003623529, 0.004930741, 
    0.005976269, 0.006479072, 0.006746552, 0.006771077, 0.00672756, 
    0.006678434, 0.006623543, 0.006562732, 0.006495839, 0.006422706, 
    0.006343169, 0.006125172, 0.005511801, 0.004975589, 0.004522883, 
    0.004080678, 0.003665518, 0.0033502, 0.003049325, 0.002748513, 
    0.002448383, 0.00219959, 0.002093144, 0.002084839, 0.002117625, 
    0.002163464, 0.002223195, 0.002317469, 0.002557264, 0.002844552, 
    0.003158804, 0.003299701, 0.003213664, 0.003168174, 0.003136202, 
    0.003104743, 0.00307378, 0.003043293, 0.003013266, 0.002983682, 
    0.002954523, 0.002912867, 0.002824141, 0.002740883, 0.0026838, 
    0.002592769, 0.00251482, 0.002453057, 0.002390679, 0.002327689, 
    0.002264097, 0.002199907, 0.002135126, 0.00206976, 0.002003815, 
    0.001937297, 0.001870212, 0.001802567, 0.001810338, 0.001740607, 
    0.001671615, 0.001603372, 0.001535886, 0.001469166, 0.00140322, 
    0.001338056, 0.001273684, 0.001210112, 0.001147349, 0.001085404, 
    0.0009869896, 0.0008423678, 0.0007526975, 0.0007394674, 0.000751883, 
    0.0007608192, 0.0007682486, 0.0007765192, 0.0007856567, 0.0007956873, 
    0.0008066377, 0.0008185348, 0.0008314062, 0.0008722778, 0.0009924493, 
    0.00107037, 0.001108455, 0.001141442, 0.001169246, 0.001191869, 
    0.001211966, 0.001229941, 0.001245908, 0.001255953, 0.001253418, 
    0.001246825, 0.001237266, 0.001225267, 0.001210646, 0.001190571, 
    0.001149663, 0.001100371, 0.001045293, 0.001005411, 0.0009856841, 
    0.0009643571, 0.0009429543, 0.0009212832, 0.0008993522, 0.0008771695, 
    0.0008547433, 0.0008320818, 0.0008091929, 0.0007832427, 0.0007469876, 
    0.0007197889, 0.0007234168, 0.000732809, 0.0007301383, 0.0007207681, 
    0.000711504, 0.0007023447, 0.0006932892, 0.0006843361, 0.0006754845, 
    0.0006667331, 0.0006580807, 0.0006495264, 0.0006410689, 0.000632707, 
    0.000602302, 0.0006016792, 0.0006010519, 0.00060042, 0.0005997836, 
    0.0005991426, 0.000598497, 0.0005978469,
  0.0008215947, 0.0008073332, 0.0007160921, 0.0006600239, 0.0006757788, 
    0.0006776749, 0.0006797507, 0.0006826097, 0.00068627, 0.0006907496, 
    0.000696067, 0.0007033403, 0.0007455549, 0.0007865616, 0.0007803448, 
    0.0007746168, 0.000771512, 0.0007719651, 0.0007777563, 0.0007856713, 
    0.0007941315, 0.0008025919, 0.0008113952, 0.0008269335, 0.0008473535, 
    0.0008664801, 0.000884323, 0.0009008947, 0.0009098242, 0.0009105193, 
    0.0009085483, 0.0009038035, 0.000896187, 0.0008897493, 0.000885829, 
    0.0008819519, 0.0008780749, 0.0008734586, 0.000866537, 0.0008584341, 
    0.0008488515, 0.0008377525, 0.0008248028, 0.0008056118, 0.0007895163, 
    0.0007819444, 0.0007748746, 0.0007680514, 0.000761469, 0.0007551219, 
    0.0007490046, 0.0007424345, 0.0007163187, 0.0007220382, 0.0007460904, 
    0.0007467425, 0.0007452904, 0.0007438458, 0.0007424084, 0.0007409784, 
    0.0007395555, 0.0007381396, 0.0007367305, 0.0007353283, 0.000702236, 
    0.0007051631, 0.0007081267, 0.0007111271, 0.0007141646, 0.0007172396, 
    0.0007203524, 0.0007235034, 0.0007266928, 0.0007308453, 0.0007484577, 
    0.0007769989, 0.000804405, 0.0008102331, 0.0008153312, 0.0008203754, 
    0.0008253644, 0.0008302968, 0.0008351709, 0.0008400751, 0.0008466339, 
    0.0008505741, 0.0008463074, 0.0008388326, 0.0008284382, 0.0008171371, 
    0.0008087005, 0.0008011701, 0.0007939382, 0.0007867062, 0.000778996, 
    0.0007649718, 0.0007470445, 0.0007299288, 0.000713611, 0.0006980759, 
    0.0006860766, 0.0006777755, 0.000670828, 0.0006653192, 0.0006613279, 
    0.0006594213, 0.0006594704, 0.0006596578, 0.0006598452, 0.0006623194, 
    0.0006734057, 0.00070708, 0.0007500001, 0.0007952762, 0.0008339724, 
    0.000677889, 0.0005285956, 0.000528238, 0.0005371438, 0.0005506253, 
    0.0005685755, 0.0005908884, 0.0006174595, 0.0006445978, 0.0005666579, 
    0.0003831354, 0.0003569539, 0.000467671, 0.0005850336, 0.0007038631, 
    0.0008241475, 0.0009458748, 0.001069033, 0.001193609, 0.001319593, 
    0.001446971, 0.0006448536, 0.001019432, 0.001393654, 0.001767518, 
    0.00214102, 0.002514157, 0.002886925, 0.003259321, 0.003631342, 
    0.004194912, 0.007140378, 0.009984914, 0.0108731, 0.01093919, 0.01097821, 
    0.01101288, 0.01104308, 0.01106871, 0.01108964, 0.01106944, 0.009995311, 
    0.00876059, 0.008188468, 0.007629127, 0.007053604, 0.006572935, 
    0.006380109, 0.006174755, 0.005958537, 0.005742319, 0.00551362, 
    0.005277503, 0.00512685, 0.00502985, 0.004984098, 0.004987106, 
    0.004972721, 0.00492844, 0.004906388, 0.004906757, 0.00492974, 
    0.004978301, 0.004957482, 0.004919793, 0.004882103, 0.004846214, 
    0.004815625, 0.004762733, 0.004707931, 0.004662055, 0.004624731, 
    0.004586495, 0.004563839, 0.004545578, 0.004526595, 0.004507071, 
    0.004487026, 0.004466478, 0.004445446, 0.004422823, 0.004361136, 
    0.00442871, 0.004540156, 0.004466446, 0.004376607, 0.004286455, 
    0.004195994, 0.004105225, 0.004014151, 0.003922775, 0.003831098, 
    0.003739124, 0.002406857, 0.002294528, 0.00218275, 0.002071527, 
    0.001960864, 0.001850765, 0.001741234, 0.001632277, 0.001523897, 
    0.001423677, 0.001427787, 0.001403489, 0.001283178, 0.001246579, 
    0.001213012, 0.001180055, 0.001147729, 0.001116054, 0.001085051, 
    0.001053214, 0.0009789161, 0.0009523655, 0.00109021, 0.001231703, 
    0.001369786, 0.001483003, 0.001529896, 0.001544324, 0.001549459, 
    0.001554593, 0.001559855, 0.001528068, 0.001447734, 0.001354651, 
    0.001249465, 0.001132819, 0.001099165, 0.00114862, 0.001187593, 
    0.001215657, 0.001232368, 0.001219989, 0.001198093, 0.001178388, 
    0.001158683, 0.001138596, 0.001115326, 0.001085918, 0.001048584, 
    0.001003397, 0.0009530592, 0.0009623277, 0.0009772675, 0.0009633397, 
    0.0009487682, 0.0009345379, 0.0009206386, 0.0009070602, 0.0008937928, 
    0.0008812777, 0.0008821802, 0.0008262311, 0.0007547056, 0.0007408398, 
    0.000731503, 0.000722215, 0.0007129756, 0.0007037841, 0.0006946404, 
    0.0006855439, 0.0006764942, 0.0006674909, 0.0008843731, 0.0008761554, 
    0.0008680418, 0.000860033, 0.00085213, 0.0008443337, 0.0008366451, 
    0.0008290652,
  0.0009231612, 0.0008744201, 0.0008287061, 0.000807372, 0.0007866591, 
    0.0007665801, 0.0007471482, 0.0007283765, 0.0006955127, 0.0006467514, 
    0.0006709582, 0.0007114994, 0.0007343669, 0.0007482994, 0.0007640715, 
    0.0007817391, 0.0007958937, 0.0007992784, 0.0007999723, 0.000803022, 
    0.0008092245, 0.0008208417, 0.0008469046, 0.0008701911, 0.000888339, 
    0.0009060744, 0.0009233532, 0.0009413772, 0.0009603202, 0.0009712331, 
    0.0009756659, 0.0009789044, 0.0009810183, 0.0009787241, 0.0009705717, 
    0.0009527865, 0.0009320637, 0.0009099876, 0.0008875891, 0.0008719387, 
    0.0008622205, 0.0008514019, 0.0008413109, 0.0008319258, 0.0008210214, 
    0.0008076779, 0.0008028467, 0.0008392723, 0.0008534071, 0.0008548178, 
    0.0008563917, 0.0008581256, 0.0008600159, 0.0008620595, 0.0008716868, 
    0.0008677295, 0.0008442826, 0.0008392354, 0.0008341484, 0.0008290217, 
    0.0008238558, 0.0008186508, 0.000813407, 0.0008081247, 0.0007894966, 
    0.0007908178, 0.0007921995, 0.000793642, 0.0007951458, 0.0007967111, 
    0.0007983385, 0.0008000282, 0.0008148855, 0.0008352463, 0.0008424617, 
    0.0008472492, 0.0008520188, 0.0008567699, 0.0008615019, 0.0008662141, 
    0.0008695317, 0.0008699403, 0.0008747812, 0.0008778133, 0.0008763108, 
    0.0008729572, 0.0008691272, 0.0008648041, 0.0008603083, 0.0008579004, 
    0.0008565499, 0.000852353, 0.000845815, 0.0008352042, 0.0008105496, 
    0.0007877511, 0.0007690429, 0.0007509767, 0.000733594, 0.000710964, 
    0.0006935404, 0.0006888087, 0.0006847124, 0.0006817725, 0.0006799289, 
    0.0006788309, 0.000680431, 0.0006958326, 0.0007189334, 0.0007470654, 
    0.0007768305, 0.0007987265, 0.0007935334, 0.0007800959, 0.0007726743, 
    0.0007710902, 0.0007312358, 0.0006232786, 0.0005130275, 0.0001663895, 
    0.0002267216, 0.0004406308, 0.0006745523, 0.0009281025, 0.001200902, 
    0.001492572, 0.001801931, 0.002202737, 0.002794546, 0.003040556, 
    0.003288203, 0.003537474, 0.00378836, 0.004040849, 0.00429493, 
    0.00455059, 0.004985541, 0.0050976, 0.005216791, 0.005343161, 
    0.005476757, 0.005617626, 0.005765817, 0.005921377, 0.005751631, 
    0.006993296, 0.007937824, 0.00827382, 0.008614684, 0.008960477, 
    0.009311267, 0.009667119, 0.01012156, 0.01043838, 0.009190186, 
    0.007777534, 0.007189416, 0.006968846, 0.006732603, 0.006480212, 
    0.006254785, 0.006186235, 0.006226688, 0.006305771, 0.006404203, 
    0.006496931, 0.00654692, 0.006578842, 0.006583085, 0.006593281, 
    0.006609548, 0.006622695, 0.006532433, 0.006354307, 0.006184276, 
    0.006019029, 0.005858541, 0.005687483, 0.005531556, 0.005501015, 
    0.00550813, 0.005534859, 0.005577587, 0.005572101, 0.005474311, 
    0.005356274, 0.005243536, 0.005135965, 0.005039091, 0.004975281, 
    0.004951199, 0.004980405, 0.004940258, 0.004868015, 0.004797311, 
    0.004728123, 0.00466043, 0.00459421, 0.004582142, 0.004493081, 
    0.004284229, 0.004155776, 0.004027828, 0.003900382, 0.003773435, 
    0.003646985, 0.003521028, 0.003395562, 0.003391001, 0.003257698, 
    0.003124019, 0.002989959, 0.002855517, 0.002720691, 0.002585477, 
    0.002449874, 0.002105928, 0.00184453, 0.001850384, 0.001835028, 
    0.00181889, 0.001801949, 0.001784188, 0.001765587, 0.001853702, 
    0.002124931, 0.002073274, 0.001977063, 0.00191102, 0.001855291, 
    0.001792391, 0.00172211, 0.001681314, 0.001729458, 0.001812174, 
    0.001904508, 0.001991252, 0.002050027, 0.002008496, 0.001962775, 
    0.001932681, 0.001888658, 0.001830049, 0.001779605, 0.001757124, 
    0.001762343, 0.001772172, 0.001763033, 0.001735782, 0.001707207, 
    0.001680784, 0.001685961, 0.001675736, 0.001640218, 0.001580074, 
    0.00151773, 0.001457609, 0.001381993, 0.001299215, 0.001209494, 
    0.001124062, 0.001051749, 0.0009980919, 0.001188445, 0.001240902, 
    0.001221633, 0.001201983, 0.001181958, 0.001161565, 0.001140811, 
    0.001106465, 0.00111339, 0.00113364, 0.001122482, 0.001111187, 
    0.001099756, 0.001088189, 0.001076487, 0.001064651, 0.001052681, 
    0.001021842, 0.001008083, 0.000994471, 0.0009810055, 0.0009676879, 
    0.000954519, 0.0009415, 0.0009286317,
  0.000896978, 0.0008799646, 0.0008629503, 0.0008459346, 0.0008289168, 
    0.0008125302, 0.0008166017, 0.000756188, 0.0006933966, 0.0006733584, 
    0.0006562853, 0.0006403467, 0.0006255748, 0.0006183901, 0.0006453622, 
    0.0006793879, 0.0007232833, 0.000741323, 0.0007483428, 0.0007564161, 
    0.0007655933, 0.0007709393, 0.0007694193, 0.0007862809, 0.0008148713, 
    0.0008411838, 0.0008593563, 0.0008739923, 0.0008870388, 0.0009047506, 
    0.0009234551, 0.0009347048, 0.000940742, 0.0009472861, 0.0009559219, 
    0.0009543334, 0.0009478566, 0.0009409715, 0.000933697, 0.0009180277, 
    0.0008942769, 0.0008718719, 0.0008497309, 0.0008469649, 0.0008495448, 
    0.0008518404, 0.0008538586, 0.0008570987, 0.000890751, 0.0009247239, 
    0.0009187419, 0.0009120198, 0.0009050639, 0.0008977696, 0.000890143, 
    0.00088219, 0.0008591554, 0.000841686, 0.0008338524, 0.0008261809, 
    0.0008184894, 0.0008107779, 0.0008030467, 0.0007952959, 0.0007447067, 
    0.0007473787, 0.0007500406, 0.0007526921, 0.0007553332, 0.0007579638, 
    0.0007608443, 0.0007731508, 0.0007903713, 0.0008016946, 0.0008128576, 
    0.0008238573, 0.0008346909, 0.0008455451, 0.0008603783, 0.0008669033, 
    0.000869257, 0.0008720293, 0.0008744974, 0.0008765532, 0.0008781862, 
    0.0008752816, 0.0008630277, 0.0008471823, 0.0008287466, 0.0008230492, 
    0.0008216447, 0.000819622, 0.0008169466, 0.000813621, 0.000808309, 
    0.0007896197, 0.0007623963, 0.0007355314, 0.000712236, 0.0006955886, 
    0.0006863023, 0.0006784762, 0.0006741636, 0.0006774137, 0.0006821809, 
    0.000681472, 0.0006727813, 0.0006685632, 0.0006670173, 0.0006656246, 
    0.0006643797, 0.0006383893, 0.0005644041, 0.000525839, 0.0005050619, 
    0.0004491813, 0.0004750706, 0.0005281418, 0.0006076822, 0.0007030497, 
    0.0007347677, 0.0007567678, 0.0006650846, 0.001153427, 0.001669334, 
    0.002199389, 0.002743372, 0.003301067, 0.005653891, 0.01167343, 
    0.0121229, 0.01242298, 0.01272062, 0.01301582, 0.01330859, 0.01359895, 
    0.006106251, 0.006009297, 0.00591812, 0.005832752, 0.005753225, 
    0.005679568, 0.005651631, 0.006967605, 0.006958197, 0.006991637, 
    0.007030461, 0.007074762, 0.007124641, 0.007176133, 0.007098574, 
    0.007382647, 0.007643722, 0.007596015, 0.007524721, 0.007442334, 
    0.007348584, 0.007186629, 0.006979362, 0.006738169, 0.006443815, 
    0.006366411, 0.00635922, 0.006353027, 0.006347857, 0.006350928, 
    0.006353294, 0.006376228, 0.006405102, 0.006400875, 0.006337913, 
    0.006263965, 0.006197332, 0.006120859, 0.006031633, 0.005930156, 
    0.005797069, 0.005632889, 0.005442989, 0.005293253, 0.005172895, 
    0.005050936, 0.004927442, 0.004815473, 0.004689557, 0.00459001, 
    0.004503376, 0.004460911, 0.004428978, 0.004400979, 0.004376801, 
    0.004360361, 0.004432923, 0.004510758, 0.004485934, 0.004444385, 
    0.004404186, 0.004365887, 0.004329455, 0.004294857, 0.004261529, 
    0.004320304, 0.00420966, 0.004094806, 0.003980204, 0.003865852, 
    0.003751748, 0.003637893, 0.003172261, 0.003050965, 0.002929247, 
    0.002807103, 0.002684533, 0.002561533, 0.002438482, 0.002318006, 
    0.002160114, 0.002144809, 0.002129118, 0.002113033, 0.002096544, 
    0.002076891, 0.001990221, 0.002340479, 0.002755257, 0.002929624, 
    0.003086678, 0.00323809, 0.003383679, 0.003450359, 0.003239048, 
    0.003038165, 0.002821174, 0.002843229, 0.002954368, 0.003057417, 
    0.003151946, 0.003311024, 0.003584672, 0.003770097, 0.003879584, 
    0.003965961, 0.00404063, 0.004085046, 0.004096563, 0.004065012, 
    0.003990092, 0.003897409, 0.003764391, 0.003625174, 0.003490323, 
    0.003377413, 0.003278228, 0.003162294, 0.003030316, 0.002834006, 
    0.002526932, 0.002199023, 0.001847943, 0.001662687, 0.001580323, 
    0.001490627, 0.001393764, 0.001298147, 0.001361259, 0.001482061, 
    0.001531181, 0.001470134, 0.001402627, 0.001330693, 0.001254401, 
    0.001173819, 0.001149312, 0.001201608, 0.001173388, 0.001144087, 
    0.001114567, 0.001084828, 0.001054872, 0.001024701, 0.001104445, 
    0.001084088, 0.001063793, 0.001043561, 0.001023393, 0.001003288, 
    0.0009821362, 0.0009216809,
  0.0008944983, 0.0008741007, 0.0008532187, 0.0008318457, 0.0007691322, 
    0.0007565407, 0.0007599118, 0.0007514839, 0.0007428164, 0.0007339031, 
    0.0007201799, 0.0006607624, 0.0006028217, 0.0005744232, 0.0005810761, 
    0.0005918583, 0.0006039274, 0.000625937, 0.0006569887, 0.000672896, 
    0.0006766836, 0.0006855457, 0.0007023345, 0.0007189605, 0.0007389378, 
    0.0007641037, 0.0007919602, 0.0008175726, 0.0008398776, 0.0008576757, 
    0.000869672, 0.0008791205, 0.0008889769, 0.0009048532, 0.0009206365, 
    0.0009368286, 0.0009488476, 0.0009495965, 0.0009395689, 0.0009304334, 
    0.0009248048, 0.0009189021, 0.0009135958, 0.0009194068, 0.000930612, 
    0.0009353383, 0.0009255016, 0.000915185, 0.0009042242, 0.0008926349, 
    0.0008771922, 0.0008453412, 0.0008161801, 0.0008034278, 0.0007905681, 
    0.0007776025, 0.0007645327, 0.0007507383, 0.0007462854, 0.0007391307, 
    0.0007320283, 0.0007250001, 0.0007180458, 0.000711165, 0.0006951013, 
    0.0006997651, 0.000704372, 0.0007089217, 0.000713414, 0.0007179316, 
    0.0007568873, 0.0007800384, 0.000791779, 0.0008033076, 0.0008146218, 
    0.0008257186, 0.0008456788, 0.0008688181, 0.000875757, 0.0008769992, 
    0.0008776781, 0.000877781, 0.000874949, 0.0008750316, 0.0008723796, 
    0.0008665695, 0.000860491, 0.0008536621, 0.0008461089, 0.0008379886, 
    0.0008284471, 0.0008221115, 0.00081685, 0.0008080273, 0.0007967409, 
    0.0007851935, 0.0007754609, 0.0007652229, 0.0007496481, 0.0007303768, 
    0.0007222611, 0.0007261122, 0.0007273187, 0.000721766, 0.0007116002, 
    0.0006931055, 0.0006725119, 0.0006504632, 0.0006284151, 0.0005914781, 
    0.0005480125, 0.0005381179, 0.0005506109, 0.0005679752, 0.0005904211, 
    0.0004466925, 0.0003113448, 0.0003410224, 0.0005098836, 0.0008268101, 
    0.001171685, 0.001543901, 0.001753313, 0.00290455, 0.005344979, 
    0.006140809, 0.006916038, 0.007670941, 0.008405792, 0.009967686, 
    0.007381659, 0.007324641, 0.007274299, 0.007220242, 0.007162488, 
    0.007101054, 0.007882874, 0.007811261, 0.007735646, 0.00765601, 
    0.007572333, 0.007482975, 0.00695168, 0.007294535, 0.007360972, 
    0.007430963, 0.007504553, 0.007581786, 0.007633601, 0.007509967, 
    0.007477574, 0.007505003, 0.007523203, 0.00753196, 0.00751681, 
    0.007327095, 0.007077652, 0.006911983, 0.006877983, 0.006839043, 
    0.006791834, 0.006814673, 0.006890096, 0.006930145, 0.006925975, 
    0.006875943, 0.006788637, 0.00670636, 0.006674303, 0.00664396, 
    0.006598286, 0.006502802, 0.006446799, 0.006447217, 0.006422998, 
    0.006370917, 0.006264589, 0.006122272, 0.005965028, 0.005745075, 
    0.005470968, 0.005227386, 0.005043453, 0.00488191, 0.004750637, 
    0.004617108, 0.004482342, 0.00439573, 0.004364895, 0.004366922, 
    0.004347384, 0.004315683, 0.004286476, 0.004259716, 0.004250947, 
    0.004402272, 0.004619361, 0.004619049, 0.00462093, 0.004624974, 
    0.004631153, 0.004587804, 0.004187678, 0.004041917, 0.003896787, 
    0.003751509, 0.003606085, 0.003460515, 0.003092388, 0.00295228, 
    0.002812096, 0.002671836, 0.0025315, 0.002390778, 0.002131908, 
    0.002087112, 0.002107858, 0.002126099, 0.002141802, 0.002154933, 
    0.002184497, 0.002135621, 0.002183857, 0.002299463, 0.002416443, 
    0.002534845, 0.002718209, 0.003319942, 0.003911691, 0.004279289, 
    0.004381336, 0.00444897, 0.004508661, 0.004425582, 0.004206012, 
    0.004320873, 0.004698038, 0.005012002, 0.005218969, 0.005395611, 
    0.005473356, 0.005474819, 0.005454368, 0.00541726, 0.005471334, 
    0.005612578, 0.005724099, 0.005794383, 0.005771708, 0.005705618, 
    0.005636142, 0.005500097, 0.005304509, 0.005014037, 0.004638997, 
    0.004369051, 0.004194825, 0.004026035, 0.003864154, 0.003644441, 
    0.003405271, 0.003244369, 0.003165747, 0.003073246, 0.002973602, 
    0.002866964, 0.002780422, 0.00240496, 0.001794271, 0.001638618, 
    0.001477358, 0.001310566, 0.001138318, 0.001085004, 0.001343018, 
    0.001276425, 0.001208017, 0.001138582, 0.001068123, 0.0009966446, 
    0.001038603, 0.001005834, 0.0009733451, 0.0009411392, 0.0009092169, 
    0.0008777761, 0.0009244992, 0.0009144181,
  0.0008072847, 0.0007940978, 0.0007891504, 0.0008064545, 0.0007533784, 
    0.0007336136, 0.0007127852, 0.0006908645, 0.0006649123, 0.0006764206, 
    0.0006865911, 0.0006846773, 0.0006784084, 0.0006696523, 0.0006703117, 
    0.0006783389, 0.0006937491, 0.0007051126, 0.0007117275, 0.000718556, 
    0.0007291028, 0.0007624819, 0.0007953093, 0.0008267923, 0.0008522847, 
    0.0008692977, 0.0008843566, 0.000897821, 0.0009251551, 0.0009605064, 
    0.0009850485, 0.001005002, 0.001017316, 0.001018426, 0.001013242, 
    0.001000003, 0.0009939952, 0.000989279, 0.0009825836, 0.0009694247, 
    0.0009563376, 0.0009590266, 0.0009564828, 0.000947867, 0.0009375488, 
    0.0009248979, 0.0009012137, 0.0008708677, 0.0008508713, 0.0008371716, 
    0.0008242172, 0.0008119895, 0.0007854807, 0.0007558915, 0.0007468709, 
    0.0007393564, 0.0007322356, 0.0007255033, 0.0007235986, 0.0007199485, 
    0.0007164496, 0.000713021, 0.0007096624, 0.0007063736, 0.000681303, 
    0.0006869509, 0.0006926046, 0.000698264, 0.0007039292, 0.0007226026, 
    0.0007602169, 0.0007763781, 0.000792664, 0.0008090762, 0.0008262074, 
    0.0008540645, 0.0008782534, 0.0008907514, 0.0009032728, 0.00091582, 
    0.0009274134, 0.0009209174, 0.0009117306, 0.0009101576, 0.0009081787, 
    0.0009052457, 0.0008985343, 0.0008887615, 0.0008843652, 0.0008810013, 
    0.0008762608, 0.0008707981, 0.0008667598, 0.0008713316, 0.000872531, 
    0.0008720201, 0.0008619791, 0.0008454346, 0.0008267024, 0.0008084149, 
    0.0007860348, 0.0007621914, 0.000743222, 0.0007219278, 0.0006945984, 
    0.0006624935, 0.0006368381, 0.0006118732, 0.0005883074, 0.0005802027, 
    0.0005767257, 0.0005739451, 0.0005595238, 0.0005545776, 0.0006308682, 
    0.0007478934, 0.0008729294, 0.000977718, 0.0007911375, 0.0007755414, 
    0.001379805, 0.001998049, 0.002602946, 0.00319514, 0.00531881, 
    0.007140937, 0.00742384, 0.007626266, 0.007809144, 0.007972714, 
    0.005822144, 0.005254441, 0.00533726, 0.005420939, 0.005505475, 
    0.005590865, 0.006932634, 0.007048982, 0.007162392, 0.007272854, 
    0.007380357, 0.007176843, 0.00675344, 0.006829655, 0.006902276, 
    0.006971257, 0.007065773, 0.007306064, 0.007383614, 0.007448484, 
    0.007504221, 0.007550649, 0.007602432, 0.0078109, 0.007927052, 
    0.007957971, 0.007965066, 0.007951137, 0.007914322, 0.007873276, 
    0.007971865, 0.008058363, 0.008092282, 0.008134041, 0.008246671, 
    0.008801584, 0.009165365, 0.009473234, 0.009300694, 0.008866617, 
    0.008414, 0.007665024, 0.007211255, 0.007197417, 0.007115521, 
    0.007040026, 0.006909614, 0.006621189, 0.006350096, 0.006094104, 
    0.005982486, 0.005841566, 0.005696992, 0.005527956, 0.005264428, 
    0.004844775, 0.004501975, 0.004316244, 0.004133115, 0.00395645, 
    0.003852368, 0.00379566, 0.003752709, 0.003735836, 0.003719966, 
    0.00370513, 0.003942944, 0.004172648, 0.004167148, 0.004152673, 
    0.004140018, 0.004129162, 0.004230054, 0.004394126, 0.004264729, 
    0.004136094, 0.004008218, 0.003881098, 0.002716564, 0.002570202, 
    0.002423714, 0.002277101, 0.002130362, 0.002082031, 0.002147964, 
    0.002246312, 0.002337583, 0.002421694, 0.002542229, 0.002914126, 
    0.003035434, 0.003125171, 0.003213654, 0.003300876, 0.003282151, 
    0.003328932, 0.00345547, 0.003623111, 0.003841601, 0.004095436, 
    0.00445664, 0.004863481, 0.004912619, 0.004920394, 0.00502933, 
    0.005133905, 0.005266854, 0.005572166, 0.00583949, 0.00610654, 
    0.00619422, 0.006202313, 0.006205341, 0.006127905, 0.006130226, 
    0.0062223, 0.006248825, 0.006257548, 0.006313848, 0.00638211, 
    0.006429708, 0.006359951, 0.006171728, 0.005933081, 0.005692342, 
    0.005378258, 0.005192346, 0.005473615, 0.00563938, 0.005582016, 
    0.005510201, 0.0054109, 0.005377719, 0.005308296, 0.004922206, 
    0.004601105, 0.004279363, 0.003956909, 0.003179276, 0.003034021, 
    0.002919771, 0.002743043, 0.00256394, 0.002382489, 0.002115832, 
    0.001746466, 0.001616367, 0.001485087, 0.001352628, 0.001218998, 
    0.00102181, 0.0009545038, 0.0008879392, 0.0008221195, 0.0007570475, 
    0.0007642998, 0.0008339015, 0.000820553,
  0.0007167737, 0.00073603, 0.0009036562, 0.000908633, 0.000892792, 
    0.0008766352, 0.0008350598, 0.0007651377, 0.0007363226, 0.0007334651, 
    0.0007284158, 0.0007269679, 0.000742819, 0.0007672268, 0.0007869021, 
    0.0008033557, 0.0008202068, 0.0008430827, 0.0008463645, 0.00085072, 
    0.0008671134, 0.0008901873, 0.0009181147, 0.0009680852, 0.001015893, 
    0.001025099, 0.001024555, 0.001026954, 0.001034321, 0.001045128, 
    0.001059128, 0.001066064, 0.001050063, 0.001031033, 0.001016405, 
    0.001005828, 0.0009982238, 0.0009951353, 0.0009909429, 0.0009806174, 
    0.00096902, 0.0009561408, 0.0009435228, 0.000904783, 0.0008602511, 
    0.0008398335, 0.0008255937, 0.0008106161, 0.0007980912, 0.0007993003, 
    0.0007950395, 0.0007898457, 0.0007862972, 0.0007842024, 0.0007697212, 
    0.0007630357, 0.0007610607, 0.0007596301, 0.0007593149, 0.0007808576, 
    0.000782016, 0.000780493, 0.0007790014, 0.000777541, 0.0007560059, 
    0.0007573407, 0.0007587976, 0.0007603768, 0.0007653118, 0.0008022625, 
    0.0008127834, 0.0008227665, 0.0008331182, 0.0008459097, 0.0008623849, 
    0.0008679564, 0.0008725765, 0.0008774622, 0.0008799407, 0.0008902644, 
    0.0009005187, 0.0009026551, 0.0009047386, 0.0009068704, 0.0009017126, 
    0.0008945739, 0.0008950492, 0.0008966204, 0.0008976848, 0.0008999347, 
    0.0008945852, 0.0008879241, 0.000883512, 0.0008822101, 0.0008833542, 
    0.0008749357, 0.0008692002, 0.0008890264, 0.0009090729, 0.0009105997, 
    0.0008987477, 0.0008784989, 0.0008421692, 0.0007992099, 0.0007576997, 
    0.0007179098, 0.0006889908, 0.0006619731, 0.0006252052, 0.000577173, 
    0.0005483117, 0.0005608459, 0.00058687, 0.00062066, 0.0006671881, 
    0.0005539788, 0.000495918, 0.0007004265, 0.0009708395, 0.001274628, 
    0.001800227, 0.002520847, 0.003162763, 0.003694116, 0.004208549, 
    0.00478085, 0.004478062, 0.004334057, 0.004436063, 0.004533516, 
    0.004605534, 0.005301498, 0.005516497, 0.005645894, 0.005777267, 
    0.005910608, 0.005945837, 0.006116505, 0.006286905, 0.006457036, 
    0.006647305, 0.006754257, 0.006859637, 0.006992622, 0.007119274, 
    0.007267856, 0.007721227, 0.007954829, 0.008091124, 0.008222987, 
    0.008297659, 0.008363739, 0.008445416, 0.008545848, 0.008629723, 
    0.008709216, 0.008681938, 0.008588925, 0.008588009, 0.008606331, 
    0.008632938, 0.00865139, 0.008340389, 0.00797391, 0.007796893, 
    0.007860672, 0.008153198, 0.00843609, 0.008554537, 0.008191983, 
    0.007701761, 0.007380081, 0.007192895, 0.007069958, 0.007047096, 
    0.007007238, 0.006760895, 0.006507729, 0.006296392, 0.006138208, 
    0.006086542, 0.006182594, 0.006214739, 0.005938861, 0.005689269, 
    0.00544028, 0.00509699, 0.00456786, 0.004108507, 0.003899682, 
    0.003729042, 0.003565812, 0.003430659, 0.003380974, 0.00340788, 
    0.003442693, 0.003481823, 0.003553617, 0.00367928, 0.003698577, 
    0.003704246, 0.003706482, 0.003758854, 0.003978865, 0.003848248, 
    0.003720172, 0.00359279, 0.0034661, 0.003166264, 0.003022392, 
    0.002877511, 0.002731617, 0.002478003, 0.001730709, 0.001998177, 
    0.002244655, 0.002483314, 0.00297976, 0.004270845, 0.004541281, 
    0.004673368, 0.00479723, 0.004700304, 0.004269657, 0.004158625, 
    0.004279992, 0.004376774, 0.0045017, 0.004789947, 0.005125465, 
    0.005372032, 0.00555225, 0.005727076, 0.005832914, 0.005955341, 
    0.006055465, 0.006131846, 0.006242039, 0.006385144, 0.006459327, 
    0.006496041, 0.00650455, 0.006502255, 0.006538265, 0.006599906, 
    0.006706115, 0.006872876, 0.007019945, 0.006924472, 0.006722665, 
    0.00657359, 0.006497028, 0.006508959, 0.006718986, 0.006650073, 
    0.005906252, 0.005709137, 0.005509654, 0.005445311, 0.005889095, 
    0.006376924, 0.006343888, 0.006210258, 0.006022959, 0.005439161, 
    0.004827919, 0.00466563, 0.004430315, 0.004193324, 0.004122887, 
    0.003690095, 0.003190284, 0.002872114, 0.002553854, 0.002196417, 
    0.002183602, 0.002083037, 0.00192763, 0.001772482, 0.001617592, 
    0.001465338, 0.001361757, 0.001258543, 0.001155699, 0.001028436, 
    0.0007993139, 0.0007739355, 0.0007447547,
  0.0008547141, 0.0008152785, 0.0008720295, 0.0008837907, 0.0008960316, 
    0.0009214358, 0.0007865159, 0.0007552971, 0.0007434525, 0.0007503293, 
    0.0008171439, 0.0008661963, 0.0008731609, 0.000879872, 0.0008806252, 
    0.0008773659, 0.0009069309, 0.0009359546, 0.0009586629, 0.0009753905, 
    0.0009847659, 0.001005032, 0.001062752, 0.001102151, 0.001134237, 
    0.001140009, 0.001121615, 0.001087436, 0.001067677, 0.001069716, 
    0.001067172, 0.001049357, 0.00101884, 0.0009864939, 0.0009569354, 
    0.0009793235, 0.001005027, 0.0009956848, 0.0009698173, 0.0009333102, 
    0.0008905603, 0.000833114, 0.000790116, 0.0007556016, 0.0007207522, 
    0.000706411, 0.0007242166, 0.000731642, 0.0007403814, 0.0007545362, 
    0.0007932268, 0.0008106987, 0.0008223637, 0.0008356613, 0.000847318, 
    0.00085583, 0.0008651767, 0.0008735574, 0.0008822672, 0.0009023626, 
    0.0009088864, 0.0009038099, 0.0008985943, 0.0008932401, 0.000883973, 
    0.0008754163, 0.0008671139, 0.0008590666, 0.000844221, 0.0008476357, 
    0.0008547847, 0.0008625154, 0.0008773849, 0.0009181401, 0.0009268828, 
    0.0009341056, 0.0009414514, 0.0009382434, 0.0009166828, 0.0009135917, 
    0.0009133228, 0.0009159509, 0.0009346904, 0.0009477431, 0.0009462401, 
    0.0009440148, 0.0009407823, 0.0009410147, 0.0009459735, 0.0009397931, 
    0.0009311597, 0.0009217082, 0.0009042375, 0.0008844964, 0.0008636987, 
    0.0008519567, 0.000843491, 0.0008493964, 0.0008599235, 0.0008763989, 
    0.0008897745, 0.0008895796, 0.0008810211, 0.0008619963, 0.0008370246, 
    0.0008079702, 0.0007614911, 0.00068523, 0.0006073196, 0.0005763834, 
    0.000569126, 0.000583615, 0.00062758, 0.0006047296, 0.0006154404, 
    0.0006537042, 0.0006802842, 0.0007920833, 0.001087766, 0.001475036, 
    0.001812686, 0.002173946, 0.003122917, 0.004008229, 0.004463202, 
    0.004941554, 0.005126063, 0.004691198, 0.004954428, 0.005183103, 
    0.005409667, 0.005448715, 0.005102774, 0.005194278, 0.005282953, 
    0.005368808, 0.006326042, 0.006574166, 0.006820029, 0.007063622, 
    0.007098259, 0.007223035, 0.007445198, 0.007664811, 0.007879768, 
    0.008192736, 0.00844382, 0.008653469, 0.008858921, 0.008977191, 
    0.00888845, 0.009024842, 0.00919382, 0.009451129, 0.01022484, 0.01066259, 
    0.01055842, 0.01043146, 0.01007095, 0.00948812, 0.009742114, 0.00980232, 
    0.009696011, 0.009386506, 0.008513357, 0.007658685, 0.007952978, 
    0.008178812, 0.008233212, 0.008188119, 0.007994944, 0.007611807, 
    0.007272108, 0.007083576, 0.006916985, 0.006814213, 0.006747745, 
    0.00667255, 0.006602026, 0.006525883, 0.006472406, 0.006305098, 
    0.006068343, 0.005759687, 0.00538969, 0.004855662, 0.004466268, 
    0.004163817, 0.00386036, 0.003552113, 0.003489548, 0.003478425, 
    0.003455121, 0.003449038, 0.003635746, 0.003926971, 0.004022971, 
    0.004122522, 0.004222177, 0.004207828, 0.004157287, 0.004109181, 
    0.004056284, 0.003844972, 0.00353399, 0.003388779, 0.003242744, 
    0.003095887, 0.003098838, 0.003018955, 0.002937564, 0.002854663, 
    0.002488669, 0.002309376, 0.002623449, 0.002932869, 0.003424428, 
    0.005439143, 0.006033489, 0.006291258, 0.006533574, 0.005966833, 
    0.004926363, 0.004828253, 0.004842143, 0.004945705, 0.005511821, 
    0.006009546, 0.006194046, 0.006360969, 0.00652166, 0.00663879, 
    0.006683971, 0.006712936, 0.00676751, 0.006837241, 0.006895027, 
    0.006903021, 0.006884141, 0.006894739, 0.006910475, 0.006808821, 
    0.006717444, 0.006664064, 0.006873181, 0.007339453, 0.007843975, 
    0.008416644, 0.008813687, 0.009126945, 0.009322683, 0.01000535, 
    0.0105767, 0.01049265, 0.01001165, 0.008849075, 0.00702699, 0.006966998, 
    0.007150022, 0.00709584, 0.007101508, 0.006827631, 0.006154244, 
    0.005837315, 0.005597353, 0.005394393, 0.005602266, 0.005378282, 
    0.004959429, 0.004538946, 0.003919835, 0.003173669, 0.002933042, 
    0.002651393, 0.002369346, 0.002253616, 0.002124212, 0.001977192, 
    0.001830996, 0.00168562, 0.00146357, 0.001374094, 0.001283948, 
    0.00119313, 0.001156533, 0.00107378, 0.00101091, 0.0009488162,
  0.0008499662, 0.0007517641, 0.0007313549, 0.0007093755, 0.0007887197, 
    0.0009478268, 0.0009754279, 0.0009983139, 0.0009560653, 0.0008839011, 
    0.0008987023, 0.0009161858, 0.0009438872, 0.0009659713, 0.0009438188, 
    0.0009443238, 0.000947129, 0.00096111, 0.0009873027, 0.001008999, 
    0.001028899, 0.001052312, 0.001088467, 0.001123549, 0.001143505, 
    0.001147013, 0.001138188, 0.001116501, 0.00109348, 0.001074862, 
    0.001056465, 0.001029603, 0.0009883918, 0.0009459291, 0.0009330591, 
    0.0009285102, 0.0009241466, 0.0009102703, 0.0008584197, 0.0008165282, 
    0.0008000255, 0.0007846793, 0.0007533476, 0.0007148796, 0.0007067309, 
    0.0007130333, 0.0007268261, 0.0007676288, 0.0008126322, 0.0008446359, 
    0.0008781691, 0.0009084066, 0.000957396, 0.0009881589, 0.001018588, 
    0.001053225, 0.001096546, 0.001107694, 0.001118017, 0.001127593, 
    0.001123544, 0.001110117, 0.00109651, 0.001082696, 0.0009901389, 
    0.0009718137, 0.0009536612, 0.0009358245, 0.0009133439, 0.0009032221, 
    0.0008983948, 0.0008938582, 0.0009020466, 0.0009200624, 0.0009269255, 
    0.0009349069, 0.0009507822, 0.0009482329, 0.000946896, 0.0009458288, 
    0.0009247942, 0.0009008895, 0.0009097867, 0.0009206901, 0.000941426, 
    0.0009756568, 0.0009879536, 0.0009960464, 0.001002652, 0.001007212, 
    0.001003619, 0.0009893527, 0.0009748495, 0.0009553128, 0.0009303078, 
    0.0009430221, 0.0009488432, 0.0009502816, 0.0009505484, 0.0009557788, 
    0.0009347023, 0.0008915027, 0.000866931, 0.0008569944, 0.0008663181, 
    0.0008846908, 0.0008800667, 0.0008700513, 0.000861702, 0.0008453829, 
    0.0008459475, 0.0008405988, 0.0008351575, 0.0008252679, 0.0007533282, 
    0.0007518044, 0.0008017409, 0.0008488381, 0.0008533779, 0.0004690211, 
    0.0003679645, 0.0007848222, 0.001205395, 0.00237438, 0.00358942, 
    0.004195911, 0.004802284, 0.005600413, 0.007918324, 0.00826762, 
    0.008578902, 0.008610162, 0.00510957, 0.005130595, 0.005198204, 
    0.005266453, 0.006633791, 0.006987378, 0.007339893, 0.007690265, 
    0.007754554, 0.008011205, 0.008312098, 0.008611537, 0.009045206, 
    0.009274669, 0.009479834, 0.009679803, 0.009811556, 0.01001494, 
    0.01022443, 0.01043639, 0.01066272, 0.01092367, 0.01118529, 0.01137546, 
    0.01137322, 0.01090711, 0.01058597, 0.01073624, 0.01086677, 0.01109746, 
    0.01135988, 0.0115606, 0.01184549, 0.01231602, 0.01390106, 0.01385512, 
    0.0139912, 0.01332138, 0.01209015, 0.01016486, 0.008592875, 0.007577594, 
    0.006596746, 0.005851947, 0.005587565, 0.005233787, 0.005428829, 
    0.005098102, 0.004614853, 0.004396067, 0.004497864, 0.004470521, 
    0.004157827, 0.003830619, 0.003404153, 0.003228596, 0.003139186, 
    0.003074024, 0.003070764, 0.003233558, 0.003458481, 0.003641411, 
    0.003827824, 0.004316356, 0.00473763, 0.00481885, 0.004895871, 
    0.004927164, 0.004901492, 0.004807312, 0.0047115, 0.00456848, 
    0.004197764, 0.004018233, 0.003839043, 0.003659411, 0.003175289, 
    0.003070422, 0.002966712, 0.00286666, 0.003040047, 0.003379765, 
    0.003748039, 0.004117523, 0.005225632, 0.0062282, 0.006767121, 
    0.007307287, 0.007511064, 0.006795798, 0.006787769, 0.00679856, 
    0.007190526, 0.007700513, 0.007835452, 0.007909422, 0.007829463, 
    0.00758685, 0.007792909, 0.00799084, 0.008181096, 0.008312558, 
    0.008358429, 0.008383198, 0.008396914, 0.008353617, 0.008282222, 
    0.008621965, 0.008829132, 0.008835169, 0.008645792, 0.008500185, 
    0.008470574, 0.008588645, 0.008881054, 0.009205962, 0.009716212, 
    0.01011169, 0.01095362, 0.01123922, 0.01132306, 0.01069948, 0.009008897, 
    0.007755488, 0.00753484, 0.007511023, 0.008272675, 0.007972617, 
    0.007440897, 0.007088289, 0.006781018, 0.007075228, 0.006887978, 
    0.006123284, 0.005265744, 0.004372436, 0.004375961, 0.003910473, 
    0.003397324, 0.002983354, 0.002670557, 0.002178835, 0.001678567, 
    0.001197177, 0.001660681, 0.001488082, 0.001303692, 0.001118178, 
    0.001409572, 0.001336495, 0.001262784, 0.001185991, 0.001060849, 
    0.001038788, 0.0009969909, 0.0009557298,
  0.0008559796, 0.0008698052, 0.0008817408, 0.0009367511, 0.0009092678, 
    0.0009050228, 0.0009045794, 0.0009440907, 0.000964452, 0.0009692429, 
    0.0009777838, 0.001013502, 0.001049887, 0.001061488, 0.001069813, 
    0.001064781, 0.00105907, 0.001061496, 0.001068214, 0.001077193, 
    0.00110155, 0.001133663, 0.001152203, 0.001164079, 0.001169902, 
    0.001169345, 0.001168599, 0.001158428, 0.00113476, 0.001093582, 
    0.001044558, 0.001017362, 0.00100149, 0.0009807135, 0.0009519846, 
    0.0009279018, 0.0009111151, 0.0008974447, 0.0008796437, 0.0008676504, 
    0.0008709832, 0.0008722342, 0.000856596, 0.000841236, 0.0008069715, 
    0.0007611825, 0.0007711576, 0.0007912892, 0.0008389683, 0.000929166, 
    0.0009931956, 0.001053572, 0.001130653, 0.001175768, 0.001197471, 
    0.001217302, 0.00123992, 0.001243015, 0.001241101, 0.001238702, 
    0.001209194, 0.00118294, 0.001164796, 0.001146744, 0.001096164, 
    0.001077704, 0.001059082, 0.001035172, 0.001012465, 0.00100254, 
    0.0009927958, 0.000991967, 0.0009784221, 0.0009692714, 0.0009612649, 
    0.0009650425, 0.0009761392, 0.0009709751, 0.0009668014, 0.0009615251, 
    0.0009512141, 0.0009409894, 0.0009282315, 0.0009014742, 0.0009277383, 
    0.0009468789, 0.0009691006, 0.0009820602, 0.0009804727, 0.0009927452, 
    0.00100852, 0.00102798, 0.001017828, 0.0009886965, 0.0009845267, 
    0.0009993144, 0.001039134, 0.001074476, 0.001094829, 0.001097074, 
    0.001084305, 0.001049748, 0.0009931384, 0.0009853075, 0.0009971702, 
    0.0009939867, 0.0009803142, 0.0009705128, 0.0009731702, 0.0009825528, 
    0.0009851464, 0.0009898506, 0.0009954614, 0.001006947, 0.001007345, 
    0.001002844, 0.0009767105, 0.0009439944, 0.0009363879, 0.0009266419, 
    0.0008348427, 0.00076046, 0.00101803, 0.001298913, 0.001659347, 
    0.002326204, 0.002948162, 0.003534172, 0.004998889, 0.005093454, 
    0.005283689, 0.005487962, 0.006018795, 0.006969673, 0.007378745, 
    0.007797393, 0.007038936, 0.007486813, 0.007933085, 0.008561647, 
    0.009371255, 0.009764478, 0.01015151, 0.01048403, 0.01085322, 0.01109416, 
    0.01133989, 0.0115083, 0.01153661, 0.01169118, 0.01187482, 0.01231954, 
    0.0125811, 0.01267777, 0.01273844, 0.01260505, 0.01231111, 0.01244298, 
    0.01264356, 0.01405624, 0.01603386, 0.0168117, 0.01712987, 0.01681314, 
    0.01914815, 0.02311167, 0.02431144, 0.0231868, 0.01871834, 0.01484923, 
    0.01385119, 0.01304167, 0.01175776, 0.01016303, 0.008449506, 0.006982205, 
    0.005492915, 0.004586642, 0.004257523, 0.00450965, 0.004268989, 
    0.003416583, 0.002766939, 0.002434212, 0.003065709, 0.003374172, 
    0.003246038, 0.002971506, 0.002848027, 0.003652379, 0.003818605, 
    0.003902602, 0.004371281, 0.004988146, 0.005208452, 0.005402798, 
    0.00558538, 0.005838114, 0.005983004, 0.006132911, 0.006122622, 
    0.005868241, 0.005833397, 0.005806476, 0.005884121, 0.005748162, 
    0.005529738, 0.005310617, 0.005225935, 0.004861091, 0.004503256, 
    0.003994718, 0.003709083, 0.003952277, 0.004216138, 0.005829875, 
    0.006935074, 0.007271945, 0.007603493, 0.007720774, 0.008880395, 
    0.009425664, 0.009902327, 0.009610871, 0.009479913, 0.009693731, 
    0.009894454, 0.009971725, 0.009579452, 0.009500431, 0.009477062, 
    0.009809166, 0.01021792, 0.01033486, 0.01035509, 0.01025096, 0.01005099, 
    0.009840114, 0.009804744, 0.009856655, 0.0100025, 0.01022677, 0.01065593, 
    0.01104219, 0.01125467, 0.0113876, 0.01129706, 0.0107258, 0.01000991, 
    0.009871581, 0.01011315, 0.01097713, 0.01158381, 0.01160308, 0.01128093, 
    0.01089025, 0.01047949, 0.009873161, 0.009332065, 0.008943346, 
    0.008865032, 0.01255797, 0.01368921, 0.01437739, 0.01166174, 0.006052906, 
    0.006067122, 0.006631104, 0.008254532, 0.007442991, 0.006834394, 
    0.006199464, 0.005061842, 0.003948243, 0.003189458, 0.002396524, 
    0.002004065, 0.001640659, 0.001259512, 0.0008726233, 0.001158932, 
    0.001063836, 0.0009698671, 0.0009582182, 0.001033425, 0.0009893527, 
    0.0009438248, 0.000847108,
  0.0008790845, 0.0008949853, 0.001044603, 0.001207278, 0.001226308, 
    0.001230708, 0.001105564, 0.001066564, 0.001061668, 0.001071622, 
    0.001101921, 0.001118213, 0.001130051, 0.001127032, 0.001122117, 
    0.001126339, 0.001133629, 0.001140262, 0.001144402, 0.001151781, 
    0.001163877, 0.001191653, 0.001212936, 0.00121694, 0.001205909, 
    0.0011797, 0.001176397, 0.001165831, 0.001131827, 0.001081322, 
    0.001028607, 0.001013982, 0.001004378, 0.0009860334, 0.000948998, 
    0.0009266594, 0.0009266579, 0.0009325683, 0.0009471448, 0.0009576469, 
    0.0009569648, 0.0009481186, 0.0009252719, 0.0009044681, 0.0008942818, 
    0.0008819418, 0.0008482845, 0.0008644837, 0.0009147155, 0.001003862, 
    0.001192443, 0.001259974, 0.001306717, 0.001301406, 0.001261086, 
    0.00125907, 0.001253481, 0.001266578, 0.00126787, 0.00126219, 
    0.001242709, 0.001223824, 0.001220345, 0.001217313, 0.00121959, 
    0.001208761, 0.001197724, 0.00119411, 0.001182008, 0.001165296, 
    0.001147219, 0.001143173, 0.001127935, 0.0011111, 0.001079124, 
    0.001043796, 0.001023071, 0.001000448, 0.0009681858, 0.0009584217, 
    0.0009537364, 0.0009658174, 0.0009616864, 0.0009492454, 0.0009440804, 
    0.0009550587, 0.001002264, 0.001021452, 0.001029308, 0.001031675, 
    0.001051623, 0.001073148, 0.00108941, 0.001104948, 0.001113575, 
    0.00113596, 0.001154943, 0.001164529, 0.00115068, 0.001130045, 
    0.001112918, 0.001106132, 0.001101661, 0.001092873, 0.001087387, 
    0.001073344, 0.001046484, 0.001031304, 0.001036018, 0.001051356, 
    0.001091084, 0.001132327, 0.00114382, 0.001147392, 0.001140703, 
    0.00112644, 0.001095527, 0.001051, 0.0009897744, 0.0009452846, 
    0.0009051089, 0.0007439006, 0.0003904896, 0.0006571365, 0.001002705, 
    0.001688163, 0.002819935, 0.003366414, 0.003767193, 0.002146384, 
    0.002599352, 0.003261462, 0.005146864, 0.006932722, 0.007689364, 
    0.008452629, 0.008427769, 0.009055394, 0.009678655, 0.01076663, 
    0.01172373, 0.01221523, 0.01263609, 0.01249758, 0.01268207, 0.01288933, 
    0.01312126, 0.01338363, 0.01357257, 0.01374023, 0.01376817, 0.01396096, 
    0.01419399, 0.01441431, 0.01452406, 0.01477884, 0.01510458, 0.01540548, 
    0.01563481, 0.01610453, 0.01684061, 0.01778432, 0.01789299, 0.01796741, 
    0.01833916, 0.01923659, 0.02047679, 0.01975243, 0.01868755, 0.01766768, 
    0.02068896, 0.02311298, 0.02293057, 0.01993798, 0.01592445, 0.0147204, 
    0.01413064, 0.01353313, 0.01279288, 0.01182098, 0.01072543, 0.00955887, 
    0.008270202, 0.007871772, 0.007750522, 0.008002465, 0.00901756, 
    0.008419398, 0.008509354, 0.008599635, 0.008230257, 0.007856202, 
    0.007995214, 0.008087225, 0.008151709, 0.00861139, 0.009112193, 
    0.009770376, 0.01027541, 0.01065132, 0.01099235, 0.01148408, 0.01183168, 
    0.01206781, 0.01257373, 0.01271459, 0.01234899, 0.01197734, 0.01102117, 
    0.01013714, 0.009264468, 0.007927125, 0.006941531, 0.006580312, 
    0.006151704, 0.007614808, 0.008442021, 0.009084444, 0.009133575, 
    0.007940213, 0.008194831, 0.008640477, 0.01094046, 0.01184735, 
    0.01223587, 0.01225657, 0.01215282, 0.01223462, 0.01229223, 0.01234579, 
    0.01291433, 0.01309854, 0.01308635, 0.01293925, 0.01275607, 0.01260711, 
    0.0125453, 0.0129013, 0.01334566, 0.01328829, 0.01293632, 0.0126096, 
    0.01236283, 0.01238942, 0.01260131, 0.01286605, 0.01309812, 0.01292491, 
    0.01259158, 0.01212385, 0.01190721, 0.01170934, 0.01167964, 0.01175301, 
    0.01196561, 0.01205862, 0.01188174, 0.01146513, 0.01001536, 0.009801862, 
    0.01022338, 0.01131789, 0.01150957, 0.009436795, 0.008879168, 0.01047397, 
    0.01827736, 0.01878444, 0.01825431, 0.01517336, 0.01367763, 0.01275846, 
    0.01179545, 0.008323735, 0.006692323, 0.005437521, 0.003895082, 
    0.002719756, 0.001982315, 0.001237293, 0.00135227, 0.001061582, 
    0.0007763044, 0.0007439958, 0.0008750043, 0.000836977, 0.0008364525, 
    0.0008766109,
  0.001116553, 0.001181516, 0.001286187, 0.001256834, 0.001226059, 
    0.001156649, 0.001137581, 0.001126938, 0.001152955, 0.001184605, 
    0.001203945, 0.001207792, 0.001192643, 0.00119218, 0.001203537, 
    0.001267111, 0.001305151, 0.001283178, 0.001228183, 0.001218841, 
    0.001261576, 0.00127504, 0.001292495, 0.001282986, 0.001225713, 
    0.001168811, 0.001129547, 0.001094047, 0.001062408, 0.001037618, 
    0.001022671, 0.001012632, 0.001011582, 0.001018536, 0.001019563, 
    0.001021979, 0.00103153, 0.001046535, 0.001055245, 0.001061065, 
    0.001037209, 0.000993612, 0.0009733471, 0.0009564659, 0.0009350615, 
    0.0009201333, 0.0009293112, 0.000967484, 0.001074485, 0.001143289, 
    0.00122387, 0.001326941, 0.001356525, 0.00139291, 0.001346838, 
    0.001324335, 0.001313978, 0.001285532, 0.001193865, 0.001150525, 
    0.001145288, 0.001327217, 0.001336426, 0.001345776, 0.001359499, 
    0.001347354, 0.001335361, 0.001334399, 0.001320517, 0.001301965, 
    0.001269742, 0.001240897, 0.001223046, 0.001209331, 0.00118204, 
    0.001154515, 0.001123392, 0.001082087, 0.001060369, 0.001041823, 
    0.001034267, 0.001045766, 0.0010468, 0.001047981, 0.001030955, 
    0.001021104, 0.001018738, 0.001013204, 0.001018764, 0.001039261, 
    0.001071344, 0.001099893, 0.001114248, 0.001142324, 0.001178754, 
    0.001215575, 0.001231791, 0.001241301, 0.001251024, 0.001252993, 
    0.001254167, 0.001257262, 0.001249564, 0.001231921, 0.001206022, 
    0.001176543, 0.001160412, 0.001154344, 0.001160249, 0.001192725, 
    0.001224961, 0.001249909, 0.001240631, 0.001196502, 0.00117893, 
    0.001165581, 0.001151561, 0.001123174, 0.00107922, 0.0009598664, 
    0.0007649845, 0.0006969526, 0.0005902249, 0.0004063772, 0.000720535, 
    0.001098464, 0.002722106, 0.003323262, 0.003752066, 0.003524902, 
    0.003522909, 0.004185895, 0.00504382, 0.006673868, 0.007558302, 
    0.008439738, 0.009572385, 0.01046312, 0.01134954, 0.01238239, 0.01307958, 
    0.01366634, 0.01409294, 0.01417343, 0.01439482, 0.01445948, 0.01448268, 
    0.01468961, 0.01487466, 0.01485051, 0.01506361, 0.01534588, 0.01577833, 
    0.01612047, 0.01642877, 0.01673461, 0.01716381, 0.01752456, 0.01780574, 
    0.01785794, 0.01802623, 0.01841456, 0.01885207, 0.01941676, 0.02003795, 
    0.02072818, 0.02162262, 0.02241703, 0.02187463, 0.02182285, 0.02294649, 
    0.02579695, 0.02609213, 0.02391874, 0.02328334, 0.02284596, 0.02280566, 
    0.0261631, 0.02826427, 0.02782984, 0.02298358, 0.0196939, 0.0198968, 
    0.0199194, 0.02161328, 0.02360537, 0.02251365, 0.01946842, 0.01564499, 
    0.01486658, 0.0140103, 0.01336696, 0.01420408, 0.01449745, 0.01487846, 
    0.01582178, 0.01635524, 0.01677104, 0.01715714, 0.01756838, 0.01788718, 
    0.01856097, 0.0189762, 0.0189719, 0.01907593, 0.01905993, 0.01830042, 
    0.01753421, 0.01451937, 0.01340105, 0.01228296, 0.009372049, 0.008312964, 
    0.00777573, 0.006309491, 0.005837661, 0.006438271, 0.007504833, 
    0.01008481, 0.01121021, 0.01223183, 0.01074896, 0.01110034, 0.01217933, 
    0.01448664, 0.01497364, 0.01481273, 0.01343095, 0.01250332, 0.01314376, 
    0.01359305, 0.01384633, 0.01376641, 0.01412895, 0.01386662, 0.01391968, 
    0.01474376, 0.01511726, 0.0154243, 0.01558317, 0.01610384, 0.01631013, 
    0.01594065, 0.01481747, 0.01406629, 0.01382772, 0.01362256, 0.01355955, 
    0.01366206, 0.01358159, 0.01343751, 0.01328406, 0.01304999, 0.01284629, 
    0.0127775, 0.0127725, 0.01292106, 0.0130793, 0.01305762, 0.01302643, 
    0.0132815, 0.01348189, 0.01344351, 0.01219296, 0.01199737, 0.01264818, 
    0.01309866, 0.01279891, 0.01305611, 0.01337893, 0.01549282, 0.01462082, 
    0.01343132, 0.01153732, 0.01024611, 0.009041631, 0.007832026, 
    0.006743997, 0.005696241, 0.004643342, 0.002759551, 0.002161574, 
    0.001569652, 0.001374557, 0.00129781, 0.001182444, 0.001106257, 
    0.001137732,
  0.001721645, 0.001413508, 0.001377413, 0.001326324, 0.001056554, 
    0.0009610981, 0.0009722775, 0.001123555, 0.001213955, 0.001265326, 
    0.001164155, 0.001245642, 0.001339659, 0.001364455, 0.00129268, 
    0.001314469, 0.001306643, 0.001169526, 0.001168108, 0.001243317, 
    0.001379441, 0.001485165, 0.001521096, 0.001467103, 0.001331093, 
    0.001167677, 0.001066127, 0.001035266, 0.001029448, 0.001019641, 
    0.001031288, 0.001050359, 0.001071145, 0.001089543, 0.001100546, 
    0.001109862, 0.001116731, 0.001117843, 0.00112457, 0.001146363, 
    0.001149292, 0.00113225, 0.001072971, 0.001054221, 0.001065369, 
    0.001080801, 0.001164888, 0.001228136, 0.00129594, 0.001313319, 
    0.001359543, 0.001371905, 0.001379872, 0.001516543, 0.001679638, 
    0.002021112, 0.002100362, 0.002127694, 0.001619243, 0.001450071, 
    0.001310598, 0.001547451, 0.001549584, 0.0015439, 0.001490403, 
    0.00147248, 0.001453563, 0.001401198, 0.00137468, 0.00134824, 
    0.001307283, 0.001288911, 0.001272976, 0.001291232, 0.001278222, 
    0.001256258, 0.001197378, 0.001166507, 0.001145785, 0.00113181, 
    0.001130558, 0.001130845, 0.001158001, 0.001152458, 0.00113139, 
    0.001106906, 0.001085009, 0.001067639, 0.001054264, 0.001060763, 
    0.001125179, 0.001172589, 0.001210947, 0.001249788, 0.001288779, 
    0.001312205, 0.001331947, 0.001346768, 0.001361066, 0.001369374, 
    0.001364353, 0.001350224, 0.001332865, 0.001320043, 0.001309752, 
    0.001300758, 0.00129076, 0.001286847, 0.001289674, 0.001302711, 
    0.001341039, 0.001320029, 0.001285449, 0.001250734, 0.001230644, 
    0.001199976, 0.001165319, 0.001147623, 0.001066305, 0.001006288, 
    0.0009178513, 0.0009134508, 0.0009264678, 0.0008068304, 0.0005298535, 
    0.000931376, 0.001318671, 0.001628403, 0.002539485, 0.003523337, 
    0.006598975, 0.007974953, 0.009201253, 0.00629953, 0.006805865, 
    0.007495991, 0.01101538, 0.0119665, 0.01289819, 0.01322228, 0.01388597, 
    0.01452943, 0.01498821, 0.01531809, 0.01564417, 0.0155996, 0.01569864, 
    0.01587672, 0.01627985, 0.01660309, 0.01688984, 0.01722531, 0.01762609, 
    0.01798677, 0.01836986, 0.01869786, 0.01897603, 0.01917732, 0.01924703, 
    0.01941964, 0.01966725, 0.01988179, 0.02017667, 0.02065725, 0.02119531, 
    0.02196697, 0.02328497, 0.02444434, 0.02520729, 0.02567064, 0.02661815, 
    0.02742743, 0.02886469, 0.03040965, 0.03056857, 0.02884406, 0.02825677, 
    0.0298716, 0.03277626, 0.02919394, 0.02611569, 0.02648504, 0.02895361, 
    0.0278256, 0.02643822, 0.0253638, 0.02214537, 0.02084174, 0.02082932, 
    0.0216356, 0.02098972, 0.02102695, 0.02141095, 0.0213829, 0.02155479, 
    0.02197929, 0.0226864, 0.02286469, 0.02301219, 0.02304325, 0.02305354, 
    0.02303423, 0.02293178, 0.02269575, 0.02243908, 0.02146228, 0.02060568, 
    0.01977439, 0.01698362, 0.01625783, 0.01561185, 0.01616459, 0.01547912, 
    0.01474242, 0.01338656, 0.01353753, 0.01412221, 0.01672363, 0.01619138, 
    0.01543141, 0.01730253, 0.01834662, 0.01840668, 0.01999778, 0.0210792, 
    0.02100311, 0.02057208, 0.01645767, 0.01460076, 0.01529447, 0.01955873, 
    0.02034165, 0.02101712, 0.02171093, 0.01601925, 0.01289505, 0.01413697, 
    0.01663062, 0.01643872, 0.01628718, 0.01715224, 0.01796867, 0.01757465, 
    0.01666919, 0.01564718, 0.01514065, 0.01485641, 0.0148754, 0.01496683, 
    0.01484744, 0.0147167, 0.01458636, 0.01447724, 0.01441664, 0.01433313, 
    0.01432787, 0.01434983, 0.01433982, 0.014029, 0.01397589, 0.01412928, 
    0.01477972, 0.01479171, 0.01468881, 0.01453917, 0.01500877, 0.0152805, 
    0.01554637, 0.01600509, 0.01595691, 0.01561651, 0.01395532, 0.01328927, 
    0.01277737, 0.01225069, 0.01093007, 0.009689236, 0.008533913, 
    0.007127277, 0.005719243, 0.003505507, 0.002901491, 0.002292129, 
    0.00200964, 0.001957031, 0.001958816, 0.002399925, 0.002057662,
  0.002417803, 0.001758274, 0.001520382, 0.001771749, 0.001983506, 
    0.001876456, 0.001381995, 0.00134536, 0.001463124, 0.001605003, 
    0.001696072, 0.001802181, 0.001829981, 0.001688606, 0.001755803, 
    0.001451801, 0.001350824, 0.001508397, 0.001852926, 0.002181288, 
    0.002363023, 0.002352623, 0.002141467, 0.001840682, 0.001594381, 
    0.00132156, 0.00118941, 0.001216189, 0.001182874, 0.001091002, 
    0.001169206, 0.001334136, 0.001331003, 0.001264016, 0.001177605, 
    0.001134617, 0.001091374, 0.001093678, 0.001132351, 0.001168989, 
    0.00120139, 0.001149928, 0.001149219, 0.0011649, 0.001226761, 
    0.001304257, 0.001431201, 0.001584405, 0.001649146, 0.001610595, 
    0.001359378, 0.001371407, 0.001507797, 0.00175074, 0.002015792, 
    0.002764663, 0.003596299, 0.003666621, 0.002802831, 0.00191187, 
    0.001555959, 0.001514346, 0.001513753, 0.001463465, 0.001542812, 
    0.001531846, 0.001518301, 0.001480582, 0.001448566, 0.001405199, 
    0.001370462, 0.001356499, 0.00137449, 0.001377956, 0.001357946, 
    0.001305849, 0.001267184, 0.001246027, 0.001252259, 0.001249675, 
    0.001241561, 0.001247929, 0.001271272, 0.001269559, 0.001209563, 
    0.001150416, 0.001132498, 0.001134045, 0.001106667, 0.001107749, 
    0.001146111, 0.001226749, 0.001284539, 0.001324907, 0.001352222, 
    0.001366945, 0.001381952, 0.001390424, 0.00139923, 0.001412445, 
    0.001418993, 0.001419516, 0.001422129, 0.00142251, 0.001412432, 
    0.001395751, 0.001366071, 0.001334791, 0.001322906, 0.001361423, 
    0.001348437, 0.001294634, 0.001241706, 0.001266748, 0.001236777, 
    0.001176923, 0.001093168, 0.001048763, 0.001019925, 0.001180243, 
    0.001214159, 0.001164661, 0.0009153609, 0.0009403228, 0.001173185, 
    0.001526613, 0.001771658, 0.001787322, 0.002512284, 0.003615769, 
    0.006209889, 0.008027151, 0.009593952, 0.01188314, 0.01334769, 
    0.01413692, 0.01064613, 0.01141125, 0.01289626, 0.01598708, 0.01687139, 
    0.01705021, 0.01662092, 0.01684286, 0.01737709, 0.01780829, 0.01802887, 
    0.01816023, 0.01841843, 0.01869805, 0.01907908, 0.01944164, 0.01977558, 
    0.0201122, 0.02048054, 0.02079448, 0.02107588, 0.02129685, 0.02152463, 
    0.02175412, 0.0220028, 0.0222551, 0.02255823, 0.02289904, 0.02315174, 
    0.02349596, 0.02398469, 0.02456393, 0.02524822, 0.02616864, 0.02658299, 
    0.02668552, 0.02771988, 0.02991933, 0.0314234, 0.0318163, 0.03240944, 
    0.03361097, 0.03468924, 0.03472659, 0.03442381, 0.03552414, 0.03520811, 
    0.03372834, 0.03256307, 0.03608278, 0.03691777, 0.03484324, 0.03198192, 
    0.0308372, 0.02951323, 0.02977225, 0.02984557, 0.0295566, 0.02889973, 
    0.02864742, 0.0278983, 0.02701809, 0.02663582, 0.02608319, 0.02558575, 
    0.02532461, 0.02516296, 0.0248791, 0.02453083, 0.02331922, 0.02282834, 
    0.02258433, 0.02241156, 0.02236948, 0.02251799, 0.02394284, 0.02388858, 
    0.02354332, 0.02354188, 0.02444094, 0.02805904, 0.03245135, 0.03364899, 
    0.02879564, 0.02411062, 0.02350582, 0.02408631, 0.02480749, 0.02514051, 
    0.02608124, 0.02710788, 0.02749817, 0.02573393, 0.02465165, 0.02499351, 
    0.02524271, 0.03000187, 0.03250623, 0.03074062, 0.02389304, 0.0217635, 
    0.02194259, 0.02027017, 0.01636804, 0.01618192, 0.01857826, 0.01965288, 
    0.01861787, 0.01798715, 0.0168868, 0.01634336, 0.01652612, 0.01649096, 
    0.01636211, 0.01625543, 0.01617618, 0.01613732, 0.01621607, 0.01621645, 
    0.01615546, 0.01609295, 0.01605596, 0.0159927, 0.0159793, 0.01595436, 
    0.01591986, 0.01579914, 0.01579477, 0.01586158, 0.0159489, 0.01590467, 
    0.01609991, 0.01671063, 0.01735478, 0.01725398, 0.0170595, 0.0163204, 
    0.01561951, 0.01447413, 0.01324934, 0.01198266, 0.009960115, 0.008212185, 
    0.006633304, 0.003122209, 0.003055546, 0.003934701, 0.007067197, 
    0.006854956, 0.005575064, 0.003958275, 0.003149339,
  0.004398178, 0.004308423, 0.005113937, 0.005226979, 0.004612932, 
    0.003959151, 0.003484639, 0.003386427, 0.004436084, 0.004518376, 
    0.004442599, 0.00495003, 0.00526281, 0.005419597, 0.005270286, 
    0.004792825, 0.004421249, 0.003988937, 0.003814303, 0.004130327, 
    0.004562837, 0.004371749, 0.0039203, 0.003182758, 0.002390682, 
    0.002000905, 0.001686248, 0.001429338, 0.001455869, 0.001638761, 
    0.001959288, 0.002156454, 0.001973639, 0.00154286, 0.001308057, 
    0.001136632, 0.00108282, 0.001049728, 0.001086489, 0.001191107, 
    0.001214206, 0.001187531, 0.001187, 0.001231083, 0.001276698, 
    0.001396838, 0.001549135, 0.001732265, 0.001925128, 0.002046651, 
    0.002077293, 0.002046576, 0.002055571, 0.001714844, 0.001657961, 
    0.002006525, 0.003984288, 0.004240484, 0.003770373, 0.002233195, 
    0.001789459, 0.001558437, 0.001468286, 0.001312375, 0.001584205, 
    0.001543092, 0.001531044, 0.001538209, 0.001500887, 0.001442931, 
    0.001409743, 0.001396363, 0.001466104, 0.001472588, 0.00145771, 
    0.001411022, 0.001397692, 0.001388197, 0.001379397, 0.001365504, 
    0.001339877, 0.001323861, 0.0013112, 0.001311644, 0.001292961, 
    0.001245895, 0.001185134, 0.001193779, 0.001203022, 0.001232728, 
    0.001267582, 0.001312026, 0.001350014, 0.001386027, 0.001412905, 
    0.001432475, 0.001432088, 0.001423824, 0.001415967, 0.001421429, 
    0.001450708, 0.001492035, 0.001531178, 0.001548903, 0.001534113, 
    0.001491955, 0.001452556, 0.001400285, 0.001370368, 0.0013435, 
    0.001302226, 0.001249839, 0.001244177, 0.001240074, 0.001149491, 
    0.00107235, 0.001027659, 0.001000131, 0.001051648, 0.001180019, 
    0.001270738, 0.001251196, 0.001186953, 0.001211036, 0.001315524, 
    0.001209308, 0.00147685, 0.001899876, 0.001810738, 0.002559826, 
    0.003376668, 0.005399637, 0.007735927, 0.0143829, 0.01782939, 0.01866922, 
    0.01079916, 0.0116498, 0.01464081, 0.01953161, 0.02075453, 0.01975152, 
    0.01913049, 0.01929823, 0.02015513, 0.02044291, 0.02047125, 0.02027157, 
    0.0204987, 0.02089374, 0.02130771, 0.02168045, 0.02201716, 0.02240781, 
    0.02283158, 0.02326109, 0.0235839, 0.02383879, 0.0240063, 0.02440417, 
    0.02484129, 0.02536381, 0.02570993, 0.02588426, 0.02594118, 0.02620484, 
    0.02645038, 0.02657227, 0.02682025, 0.02728261, 0.02769621, 0.02800919, 
    0.02817906, 0.02830775, 0.02891425, 0.02991678, 0.03019075, 0.02997342, 
    0.03060511, 0.03202534, 0.03224374, 0.03185317, 0.03168845, 0.03164826, 
    0.03214049, 0.03370491, 0.03312569, 0.03135039, 0.03100734, 0.03126445, 
    0.03068666, 0.03078145, 0.03067013, 0.02993477, 0.0294103, 0.02917386, 
    0.0286511, 0.02811116, 0.02770298, 0.02733936, 0.02706004, 0.02695703, 
    0.02687723, 0.02667627, 0.0266023, 0.02648343, 0.02685308, 0.02735204, 
    0.03165439, 0.03190928, 0.03130044, 0.02972779, 0.0293586, 0.0287183, 
    0.028456, 0.02854946, 0.02894002, 0.0291327, 0.03009058, 0.03214407, 
    0.03171682, 0.03036861, 0.02926684, 0.02850891, 0.02703112, 0.02647595, 
    0.02601364, 0.02572295, 0.02535976, 0.02518117, 0.02454891, 0.02282313, 
    0.0212022, 0.01963061, 0.01932778, 0.01990039, 0.02174569, 0.02745678, 
    0.02943743, 0.02410152, 0.02011281, 0.02157452, 0.02185565, 0.02061763, 
    0.01915215, 0.01804413, 0.01761013, 0.01783929, 0.01815535, 0.01824817, 
    0.01833187, 0.01830982, 0.01822472, 0.01818432, 0.01810605, 0.01798122, 
    0.01791865, 0.01788145, 0.01792211, 0.01788782, 0.01778177, 0.01754596, 
    0.01739995, 0.01726916, 0.0171021, 0.01706082, 0.01714928, 0.01749174, 
    0.01772275, 0.01816034, 0.018459, 0.01860704, 0.01869318, 0.01851256, 
    0.01837254, 0.017373, 0.01606389, 0.01307122, 0.0105621, 0.009052051, 
    0.008211194, 0.008545873, 0.01084547, 0.01459443, 0.01454343, 0.01119978, 
    0.008144137, 0.006047094,
  0.009100329, 0.008520901, 0.01359689, 0.01460812, 0.01235479, 0.008710956, 
    0.008180961, 0.00929861, 0.009499241, 0.008690834, 0.007753916, 
    0.008442702, 0.01094901, 0.01331892, 0.0126459, 0.01007051, 0.01060301, 
    0.01069041, 0.01012196, 0.009888779, 0.009126402, 0.007925607, 
    0.006748541, 0.005811404, 0.004882419, 0.003868736, 0.0035243, 
    0.004074375, 0.004587229, 0.004319855, 0.004117374, 0.003270986, 
    0.002662544, 0.001806666, 0.001515733, 0.001450126, 0.001295995, 
    0.001225342, 0.001234697, 0.001188174, 0.001166942, 0.001214935, 
    0.001215919, 0.001161178, 0.001152235, 0.001268451, 0.001488564, 
    0.001675297, 0.001921565, 0.002194722, 0.002519226, 0.003009042, 
    0.003270296, 0.003126146, 0.001762113, 0.001839371, 0.002903, 0.00406872, 
    0.004501408, 0.003600866, 0.003250128, 0.002984086, 0.002472189, 
    0.0018228, 0.001846484, 0.001652542, 0.001629506, 0.001668959, 
    0.001590447, 0.001496414, 0.0014409, 0.001417818, 0.001428061, 
    0.001427201, 0.001447823, 0.001466404, 0.001480219, 0.001475491, 
    0.001467013, 0.001416239, 0.001404837, 0.001419603, 0.001431814, 
    0.001407313, 0.00135681, 0.001290317, 0.001276663, 0.001261665, 
    0.001284317, 0.001335558, 0.001438202, 0.001490029, 0.00148715, 
    0.001505608, 0.001525953, 0.001540625, 0.001498761, 0.001493993, 
    0.001493587, 0.001523583, 0.001568681, 0.001609547, 0.001645752, 
    0.001667898, 0.001678544, 0.001652906, 0.001588457, 0.00154173, 
    0.001537951, 0.001506333, 0.001438349, 0.001429943, 0.001453947, 
    0.001386936, 0.001354309, 0.001311499, 0.001328435, 0.001383048, 
    0.00152829, 0.001650978, 0.001726605, 0.001770538, 0.001833041, 
    0.001589333, 0.001823118, 0.002524169, 0.004445503, 0.005568419, 
    0.005277664, 0.004562756, 0.005340681, 0.008597227, 0.01064011, 
    0.01224252, 0.01297617, 0.01412849, 0.014658, 0.01618364, 0.01969442, 
    0.02276604, 0.02358929, 0.02167103, 0.02159333, 0.02217214, 0.02285731, 
    0.02304639, 0.02275193, 0.02292083, 0.02333373, 0.02385269, 0.02417202, 
    0.02437179, 0.02468564, 0.02503899, 0.02561579, 0.0260582, 0.02635791, 
    0.02655309, 0.02689385, 0.02732125, 0.02785129, 0.02823293, 0.02853005, 
    0.02871191, 0.02893971, 0.02919837, 0.02940894, 0.0295425, 0.02971753, 
    0.03010275, 0.0304644, 0.03080481, 0.03112692, 0.03139804, 0.03164336, 
    0.03176283, 0.03210051, 0.03227922, 0.03222983, 0.0321945, 0.03249945, 
    0.032756, 0.03321956, 0.03329245, 0.03322172, 0.03299969, 0.03260304, 
    0.0322712, 0.03217556, 0.03177935, 0.03125447, 0.03109189, 0.03088165, 
    0.03076298, 0.03063871, 0.03038145, 0.03006354, 0.02985578, 0.02966233, 
    0.02955123, 0.02966971, 0.02994342, 0.03007477, 0.03054136, 0.03084423, 
    0.03109525, 0.03151148, 0.03202381, 0.03354261, 0.03377207, 0.03358038, 
    0.03292146, 0.03266753, 0.0326682, 0.03273698, 0.03252126, 0.03244563, 
    0.03271087, 0.03189976, 0.03162689, 0.03074578, 0.02960693, 0.02953827, 
    0.02971977, 0.02936683, 0.02926073, 0.02847072, 0.02756312, 0.0272548, 
    0.02690742, 0.02569723, 0.02321345, 0.02030683, 0.01934952, 0.02054977, 
    0.02090107, 0.02048428, 0.02285977, 0.02568826, 0.02425469, 0.02223559, 
    0.02362485, 0.02379234, 0.02190861, 0.02029826, 0.01970167, 0.0195474, 
    0.02006911, 0.02036144, 0.02052573, 0.0206232, 0.02048383, 0.02026576, 
    0.02008441, 0.02011671, 0.02007348, 0.01999348, 0.01990903, 0.01985862, 
    0.01982519, 0.01974132, 0.01958234, 0.01935538, 0.01928896, 0.01915285, 
    0.0189701, 0.01893831, 0.0188935, 0.01891949, 0.01909081, 0.019617, 
    0.01991578, 0.02068841, 0.02120054, 0.0212126, 0.02117689, 0.0204534, 
    0.01893976, 0.01726686, 0.01623876, 0.01495247, 0.01508196, 0.01650676, 
    0.01785585, 0.01785131, 0.01591592, 0.01438717, 0.01162958,
  0.01704672, 0.01582384, 0.01473479, 0.01401379, 0.0129546, 0.01251961, 
    0.01276979, 0.01321664, 0.01322089, 0.01102807, 0.01035659, 0.01044652, 
    0.01200516, 0.01404245, 0.01407968, 0.01255273, 0.01285886, 0.01430967, 
    0.01497417, 0.01565911, 0.01458641, 0.01355149, 0.01254849, 0.01117019, 
    0.009854652, 0.00863444, 0.008771504, 0.01093793, 0.01451174, 0.0171564, 
    0.0128201, 0.006766732, 0.004643837, 0.003621981, 0.002976614, 
    0.002467385, 0.002113166, 0.002125981, 0.001599582, 0.001581688, 
    0.00141044, 0.001210662, 0.001253396, 0.00124693, 0.001296695, 
    0.001401823, 0.001479175, 0.001563241, 0.001860175, 0.002370029, 
    0.003290094, 0.004087062, 0.005138325, 0.005420402, 0.004617678, 
    0.003444934, 0.003415806, 0.004549127, 0.005477785, 0.009254038, 
    0.01098959, 0.009259311, 0.004814223, 0.0034388, 0.002802524, 
    0.002399981, 0.002094621, 0.001968414, 0.001841422, 0.00171069, 
    0.001581736, 0.001490057, 0.001438878, 0.001454488, 0.001499958, 
    0.001557849, 0.001680165, 0.001700258, 0.001631423, 0.001563001, 
    0.001515259, 0.00155941, 0.001592764, 0.001555149, 0.001498751, 
    0.001458568, 0.001364912, 0.001562891, 0.001697969, 0.001755126, 
    0.0018768, 0.001799825, 0.001711499, 0.001707161, 0.001818676, 
    0.001806564, 0.00173823, 0.001680209, 0.001667881, 0.001784249, 
    0.001841209, 0.001797619, 0.001822587, 0.001799574, 0.00170556, 
    0.001645234, 0.001654134, 0.001637325, 0.001639255, 0.001586942, 
    0.001565715, 0.001712064, 0.001781165, 0.001778376, 0.001891092, 
    0.002079024, 0.002217801, 0.002445073, 0.002815916, 0.003144495, 
    0.00331471, 0.003395531, 0.003377733, 0.003701513, 0.00357499, 
    0.005616192, 0.009986222, 0.01446907, 0.01572, 0.01224897, 0.01290915, 
    0.01488437, 0.01637006, 0.01627682, 0.01563759, 0.01730197, 0.02463863, 
    0.02624577, 0.0264145, 0.0261547, 0.0259505, 0.02489242, 0.02483861, 
    0.02569245, 0.0260479, 0.02590062, 0.02575341, 0.02605269, 0.02684555, 
    0.02724245, 0.02726906, 0.02751063, 0.02793987, 0.02834643, 0.02870044, 
    0.02905803, 0.02942493, 0.02986689, 0.03038574, 0.03079944, 0.03126866, 
    0.03177278, 0.03200738, 0.03216838, 0.03252774, 0.03278894, 0.03295604, 
    0.03314595, 0.03338411, 0.03368632, 0.03406315, 0.03446738, 0.03481623, 
    0.03504209, 0.03508908, 0.03511139, 0.03530358, 0.03551438, 0.03570057, 
    0.03574442, 0.03559684, 0.03555827, 0.03547588, 0.03520061, 0.03489316, 
    0.03461502, 0.03420788, 0.03395312, 0.03365011, 0.03339045, 0.03337378, 
    0.03347648, 0.03351171, 0.03357949, 0.03360173, 0.03357887, 0.03344883, 
    0.03330584, 0.03306692, 0.03284641, 0.03282067, 0.03306016, 0.03327212, 
    0.03389751, 0.03429623, 0.03455603, 0.03478998, 0.03493682, 0.03418799, 
    0.03405252, 0.03380341, 0.03350984, 0.0331615, 0.03282934, 0.0326814, 
    0.03247841, 0.03241637, 0.03274488, 0.03298515, 0.03285128, 0.03263643, 
    0.03226241, 0.03189014, 0.03219702, 0.03248149, 0.03386197, 0.0342976, 
    0.033967, 0.03281288, 0.03150821, 0.02885315, 0.026349, 0.02293514, 
    0.02034315, 0.02334785, 0.0309553, 0.0286906, 0.02665764, 0.02487977, 
    0.02379579, 0.02419739, 0.02429149, 0.0236556, 0.02172381, 0.0211004, 
    0.021664, 0.02230716, 0.02268447, 0.02287122, 0.02288743, 0.02280814, 
    0.02259638, 0.02218716, 0.02204432, 0.02199242, 0.02208122, 0.02202533, 
    0.0218736, 0.02187737, 0.02185527, 0.02174888, 0.02162584, 0.02155462, 
    0.02153116, 0.02136838, 0.02120375, 0.02116597, 0.02102829, 0.02058083, 
    0.0205482, 0.02065078, 0.02097177, 0.02132641, 0.02188429, 0.02212027, 
    0.02296977, 0.02304616, 0.02305393, 0.02293352, 0.02235331, 0.02082636, 
    0.02050772, 0.02031256, 0.02020365, 0.02008603, 0.01965245, 0.01883185, 
    0.01783001,
  0.02158652, 0.02112942, 0.02076766, 0.02093717, 0.02072678, 0.0203742, 
    0.02018641, 0.01952082, 0.01916181, 0.01848803, 0.01830864, 0.0184637, 
    0.01841864, 0.01941817, 0.01936545, 0.0198949, 0.02081148, 0.0201758, 
    0.01999004, 0.02065898, 0.02078436, 0.02011767, 0.01894153, 0.01673457, 
    0.01454174, 0.01429368, 0.01655193, 0.01886255, 0.02140623, 0.0233671, 
    0.01888321, 0.01334679, 0.01024241, 0.007234108, 0.005907793, 
    0.006529467, 0.007220151, 0.006856086, 0.004706662, 0.002720512, 
    0.002037875, 0.002012472, 0.00191927, 0.001877272, 0.001775768, 
    0.001808468, 0.001801293, 0.001788274, 0.002268057, 0.002952025, 
    0.003536453, 0.004543921, 0.00627323, 0.009316626, 0.01027338, 
    0.007696514, 0.006885932, 0.006649194, 0.007380696, 0.009787989, 
    0.01081708, 0.009301495, 0.005984996, 0.004706946, 0.00368647, 
    0.003346028, 0.003158081, 0.002898086, 0.00288542, 0.002700804, 
    0.002296068, 0.001951809, 0.001737181, 0.00178575, 0.001798947, 
    0.001791412, 0.001943141, 0.002127378, 0.002126222, 0.00195612, 
    0.001676121, 0.001648843, 0.001778598, 0.00192466, 0.001881479, 
    0.001793657, 0.002318833, 0.002823448, 0.002659754, 0.002855862, 
    0.002935685, 0.003174143, 0.003153873, 0.002870697, 0.00304288, 
    0.002823343, 0.002345251, 0.002281612, 0.002319703, 0.002335067, 
    0.002348963, 0.002066858, 0.002292301, 0.002089967, 0.002033389, 
    0.001952741, 0.001822529, 0.001926287, 0.00196486, 0.001907439, 
    0.00203093, 0.002239418, 0.002426241, 0.002805484, 0.003193519, 
    0.003455104, 0.003816644, 0.004736159, 0.005991231, 0.006802457, 
    0.007256037, 0.007823344, 0.008375852, 0.009179664, 0.01056875, 
    0.01258509, 0.01482336, 0.0204487, 0.02181237, 0.0213428, 0.02222879, 
    0.02357847, 0.02500319, 0.02581843, 0.02648723, 0.02804584, 0.03137213, 
    0.03237081, 0.03087487, 0.02987167, 0.02934201, 0.02908798, 0.02913555, 
    0.02953855, 0.02981791, 0.02979131, 0.02990822, 0.03007295, 0.03044063, 
    0.03108512, 0.03156143, 0.03187837, 0.03233957, 0.03262604, 0.03285912, 
    0.03310445, 0.03344912, 0.03391185, 0.03426726, 0.03455146, 0.03477934, 
    0.03506576, 0.0352481, 0.0355153, 0.03583993, 0.0361348, 0.03638614, 
    0.03657211, 0.03677835, 0.03705826, 0.03737474, 0.03784761, 0.0382175, 
    0.03849623, 0.03856456, 0.0386273, 0.0388736, 0.0392097, 0.03943544, 
    0.03947225, 0.03940885, 0.03924349, 0.03892444, 0.03857003, 0.03799502, 
    0.03744929, 0.03710571, 0.03687743, 0.03681866, 0.03672367, 0.03674514, 
    0.03680572, 0.03687712, 0.03698212, 0.03723069, 0.03745338, 0.03750504, 
    0.03738608, 0.03718781, 0.03669676, 0.036604, 0.03654063, 0.03667402, 
    0.03682929, 0.03701352, 0.03723317, 0.03732865, 0.03739106, 0.03739729, 
    0.03720635, 0.03675129, 0.03637193, 0.0360449, 0.03582916, 0.03586024, 
    0.03612386, 0.03610555, 0.03637213, 0.03650811, 0.03655453, 0.03650141, 
    0.03645195, 0.03637525, 0.03643687, 0.03687723, 0.03741177, 0.03886518, 
    0.03964744, 0.03959062, 0.03894797, 0.03758214, 0.03367203, 0.02968609, 
    0.0308057, 0.03860651, 0.04353018, 0.03979633, 0.03122364, 0.02648096, 
    0.02515572, 0.0272907, 0.02659093, 0.02428849, 0.02299551, 0.02272493, 
    0.02372256, 0.02443653, 0.0249004, 0.02517952, 0.02514603, 0.0249776, 
    0.02471899, 0.02449141, 0.0243363, 0.02427394, 0.02424367, 0.02417065, 
    0.0240765, 0.02411743, 0.02420306, 0.02416304, 0.02412626, 0.02401358, 
    0.02382343, 0.02354065, 0.0233239, 0.02316868, 0.02298612, 0.02275834, 
    0.02256011, 0.02253233, 0.02273794, 0.02285845, 0.02288217, 0.02298024, 
    0.0232465, 0.0234867, 0.02360935, 0.02370322, 0.02343771, 0.02321171, 
    0.02290916, 0.02251778, 0.02229048, 0.02214009, 0.02202401, 0.02190822, 
    0.02186943,
  0.02275468, 0.02291653, 0.02294606, 0.02291797, 0.0229541, 0.02298411, 
    0.02319518, 0.02325083, 0.0233217, 0.02294351, 0.02269694, 0.02274576, 
    0.02306839, 0.02347953, 0.02297758, 0.02272344, 0.02255169, 0.02203631, 
    0.02190703, 0.02170551, 0.02185106, 0.02245686, 0.02217847, 0.02198286, 
    0.02127945, 0.02279422, 0.02464733, 0.02468149, 0.02391777, 0.02249625, 
    0.02088207, 0.01862012, 0.01685973, 0.01451465, 0.01549693, 0.02243349, 
    0.02122975, 0.01532549, 0.0114221, 0.007394964, 0.004925088, 0.003982954, 
    0.0040178, 0.003506174, 0.003892129, 0.004127693, 0.003564123, 
    0.003438456, 0.003592812, 0.004217834, 0.004499763, 0.005083567, 
    0.006464504, 0.01197985, 0.01426647, 0.01250445, 0.01108352, 0.01070914, 
    0.01049156, 0.0104227, 0.009784148, 0.009283567, 0.007598829, 
    0.006961418, 0.009307809, 0.008969269, 0.0086241, 0.008028169, 
    0.006967073, 0.006057765, 0.004665843, 0.003854823, 0.003273543, 
    0.003099338, 0.002905646, 0.002750613, 0.003302905, 0.00421877, 
    0.003842462, 0.002700527, 0.002213409, 0.002046972, 0.002497282, 
    0.002764126, 0.00293372, 0.003994021, 0.005654367, 0.00705604, 
    0.006113566, 0.005788269, 0.006923703, 0.00762708, 0.007649832, 
    0.007755369, 0.007519965, 0.006662814, 0.005379632, 0.004893005, 
    0.005171153, 0.005516147, 0.006062517, 0.006229423, 0.005168078, 
    0.004155916, 0.004030162, 0.003303543, 0.002862925, 0.003192305, 
    0.003214923, 0.003251225, 0.003543634, 0.004026875, 0.004816526, 
    0.006217945, 0.007116603, 0.007836801, 0.008522086, 0.009758891, 
    0.01190143, 0.01401279, 0.0155468, 0.0164955, 0.01774885, 0.01912466, 
    0.02032072, 0.0196605, 0.0205902, 0.02245707, 0.02401687, 0.02594412, 
    0.02729296, 0.02839461, 0.02962347, 0.0306268, 0.03165676, 0.03275617, 
    0.03375345, 0.03432761, 0.03416196, 0.03389052, 0.03343825, 0.03342239, 
    0.03375868, 0.03419519, 0.03470486, 0.03521675, 0.0354231, 0.0354941, 
    0.03586541, 0.03651204, 0.03689208, 0.03725148, 0.03743598, 0.03750766, 
    0.03766581, 0.03784364, 0.03808225, 0.03826254, 0.03847524, 0.03869257, 
    0.03884105, 0.03887795, 0.03891766, 0.03881309, 0.03891233, 0.03937362, 
    0.03972473, 0.03995635, 0.04004807, 0.04023871, 0.0406336, 0.04116438, 
    0.04169086, 0.0420999, 0.04246472, 0.04259864, 0.04259818, 0.04268837, 
    0.04289703, 0.04302497, 0.04295747, 0.04271776, 0.04226464, 0.04158495, 
    0.0408961, 0.04049968, 0.04027925, 0.04009466, 0.04000783, 0.03999023, 
    0.04021841, 0.04048332, 0.04060948, 0.04085787, 0.04107138, 0.04144685, 
    0.04155269, 0.04140769, 0.0412746, 0.04113008, 0.04107944, 0.04112053, 
    0.04126661, 0.04144014, 0.04159865, 0.0418148, 0.04216486, 0.04228979, 
    0.04245763, 0.04228116, 0.04190911, 0.04149976, 0.04107647, 0.04077264, 
    0.04057815, 0.04054718, 0.04024203, 0.04009325, 0.04039286, 0.04097034, 
    0.04119106, 0.04122456, 0.04124399, 0.04110047, 0.0413685, 0.04218593, 
    0.04341989, 0.04420124, 0.04525281, 0.04636003, 0.04864153, 0.04899324, 
    0.04280157, 0.04117412, 0.04478398, 0.03454597, 0.02621605, 0.02851322, 
    0.02859368, 0.02742295, 0.02608227, 0.02422001, 0.02351818, 0.02408926, 
    0.02492619, 0.02549321, 0.02606784, 0.02680774, 0.02754019, 0.02775599, 
    0.02766357, 0.0276292, 0.02741065, 0.02700002, 0.0267143, 0.02677709, 
    0.02704163, 0.02699155, 0.02700256, 0.02706377, 0.02702036, 0.0268751, 
    0.02661733, 0.0263453, 0.02606467, 0.02573766, 0.02547673, 0.02512436, 
    0.02487257, 0.02464923, 0.02454145, 0.02455457, 0.0245835, 0.02441495, 
    0.02416451, 0.02411665, 0.02412842, 0.02403564, 0.02373736, 0.0235314, 
    0.02323726, 0.02304208, 0.02306733, 0.02296398, 0.02287743, 0.0227816, 
    0.02271505, 0.02269745,
  0.02387859, 0.02382624, 0.02397162, 0.02389706, 0.02373393, 0.02352794, 
    0.02324174, 0.02305694, 0.02290985, 0.02290661, 0.02314818, 0.02352956, 
    0.02365579, 0.0234897, 0.02345756, 0.02333793, 0.02326968, 0.02327608, 
    0.02334975, 0.0234489, 0.02354726, 0.02384689, 0.02419454, 0.02447586, 
    0.02447193, 0.02484801, 0.0256831, 0.02615253, 0.02620431, 0.02600107, 
    0.02561039, 0.02615786, 0.02608047, 0.02237128, 0.0211452, 0.02405377, 
    0.02388556, 0.02244086, 0.01880492, 0.01469757, 0.01211285, 0.01077013, 
    0.01163378, 0.01110262, 0.009833529, 0.009558233, 0.009170984, 
    0.009132682, 0.009323054, 0.00934867, 0.009152327, 0.008909766, 
    0.008032642, 0.00939852, 0.01102367, 0.01233, 0.0145417, 0.01490099, 
    0.01474826, 0.01482121, 0.01549464, 0.01556648, 0.01587779, 0.01559061, 
    0.01278729, 0.01227187, 0.01156915, 0.01106797, 0.0105418, 0.009515391, 
    0.007706819, 0.007242564, 0.008260825, 0.007904949, 0.00739111, 
    0.007234997, 0.009314484, 0.009341858, 0.006563017, 0.004830703, 
    0.003654108, 0.003948086, 0.004914449, 0.006146853, 0.01154959, 
    0.01633393, 0.01206633, 0.007536747, 0.007266983, 0.01076336, 0.01529859, 
    0.01663236, 0.01467555, 0.01513542, 0.01649756, 0.01673386, 0.01413447, 
    0.01101396, 0.01090358, 0.01358119, 0.02114948, 0.02694139, 0.01920601, 
    0.01127138, 0.008621251, 0.008701597, 0.008854854, 0.008442116, 
    0.0075371, 0.007117746, 0.007577156, 0.009856638, 0.01145352, 0.01297017, 
    0.01405557, 0.01520183, 0.01699365, 0.01913753, 0.02102498, 0.02264641, 
    0.02428207, 0.02548722, 0.02680025, 0.02783836, 0.02849931, 0.02887858, 
    0.02962987, 0.02988019, 0.02994891, 0.03050123, 0.03077592, 0.03182961, 
    0.03320097, 0.03437055, 0.03527645, 0.03624547, 0.03726393, 0.03783145, 
    0.03817374, 0.03823319, 0.03794169, 0.03808952, 0.03874293, 0.03927761, 
    0.03980999, 0.0402861, 0.04060768, 0.04101941, 0.04152592, 0.04189071, 
    0.04210889, 0.04225579, 0.04220938, 0.04212701, 0.04214032, 0.04219435, 
    0.04238741, 0.04252926, 0.04268001, 0.0427813, 0.04291755, 0.04302983, 
    0.04334764, 0.0435344, 0.04341845, 0.04353544, 0.04365977, 0.04389545, 
    0.04409453, 0.04450307, 0.04509054, 0.04550561, 0.04610689, 0.04671618, 
    0.04685908, 0.04678923, 0.04662363, 0.04643991, 0.04632454, 0.04632405, 
    0.046312, 0.04616835, 0.04582935, 0.04534334, 0.04494552, 0.04467396, 
    0.044605, 0.04443663, 0.04433456, 0.04455749, 0.04478895, 0.04494883, 
    0.04515335, 0.04532028, 0.04543938, 0.04561813, 0.04585688, 0.04601916, 
    0.04615923, 0.04617488, 0.04622192, 0.0463756, 0.04707035, 0.04736881, 
    0.0474725, 0.04767037, 0.04784796, 0.04792831, 0.0479684, 0.04780838, 
    0.04741298, 0.04704349, 0.04643919, 0.0461388, 0.04586709, 0.04560539, 
    0.04519096, 0.04502203, 0.0452714, 0.04548658, 0.04618849, 0.04639725, 
    0.04621498, 0.0459068, 0.045433, 0.04527493, 0.04550327, 0.04638546, 
    0.04784979, 0.05064502, 0.05279703, 0.05360264, 0.05218739, 0.04930366, 
    0.06133253, 0.05838382, 0.03312972, 0.02886951, 0.02924831, 0.02962655, 
    0.02706174, 0.02415, 0.02301866, 0.02404788, 0.02560244, 0.02669765, 
    0.02789699, 0.02906662, 0.02999532, 0.03050725, 0.03081574, 0.03088391, 
    0.03063921, 0.03019956, 0.0295917, 0.02934606, 0.02937087, 0.02962215, 
    0.02980869, 0.02992809, 0.02978883, 0.02951575, 0.02920617, 0.02891059, 
    0.02848786, 0.02811552, 0.02782566, 0.02752646, 0.02728834, 0.02702921, 
    0.02686805, 0.02674728, 0.02664024, 0.0263679, 0.02583576, 0.0256357, 
    0.02560128, 0.02546009, 0.02512608, 0.02491895, 0.02483171, 0.02462849, 
    0.02434756, 0.02421814, 0.02425341, 0.0241759, 0.02409133, 0.02397775,
  0.02540516, 0.0253404, 0.02534527, 0.02509245, 0.02457957, 0.02429855, 
    0.0239642, 0.02368894, 0.02345101, 0.02337785, 0.02340749, 0.0237628, 
    0.02408874, 0.02416251, 0.02421799, 0.02428312, 0.02441361, 0.02459853, 
    0.0248622, 0.02508665, 0.02530929, 0.02562232, 0.02582533, 0.0258638, 
    0.02575446, 0.02585275, 0.02618013, 0.02648836, 0.02717801, 0.02801473, 
    0.02851452, 0.02900815, 0.03047085, 0.03222195, 0.03115308, 0.03049228, 
    0.03136629, 0.03014128, 0.02761288, 0.02336124, 0.01751986, 0.0172783, 
    0.02572192, 0.03181164, 0.02699309, 0.02311064, 0.01993178, 0.01904934, 
    0.01865847, 0.01836568, 0.01797795, 0.01791694, 0.01749565, 0.01749254, 
    0.01754643, 0.01812649, 0.01902781, 0.01936396, 0.01926854, 0.0193413, 
    0.01967942, 0.02001535, 0.0210894, 0.0212309, 0.02111208, 0.02083638, 
    0.02052696, 0.01990825, 0.01883951, 0.01736533, 0.01533278, 0.01460893, 
    0.01556984, 0.01550637, 0.01516662, 0.01476681, 0.01381168, 0.01398678, 
    0.01270423, 0.01058135, 0.008701781, 0.00966705, 0.01581228, 0.01587749, 
    0.01936464, 0.025114, 0.01857455, 0.0141804, 0.01267339, 0.01592669, 
    0.02229514, 0.02848536, 0.0262765, 0.02434013, 0.02441606, 0.02575066, 
    0.0237505, 0.02162653, 0.02119916, 0.02411523, 0.02748825, 0.03001131, 
    0.02602062, 0.02308333, 0.02215905, 0.02519396, 0.02157971, 0.01659795, 
    0.01424053, 0.0156422, 0.01690474, 0.01805023, 0.01771805, 0.01951773, 
    0.02246664, 0.0235376, 0.02557217, 0.02678183, 0.02739614, 0.02748981, 
    0.02811751, 0.02881647, 0.02950138, 0.02999721, 0.0306153, 0.03141242, 
    0.0321709, 0.03298458, 0.03401878, 0.0349367, 0.03579094, 0.03671444, 
    0.03816513, 0.03938277, 0.04051805, 0.04147181, 0.04238794, 0.0429473, 
    0.04318219, 0.04331934, 0.04324882, 0.04345191, 0.04384699, 0.04445818, 
    0.04506821, 0.0456293, 0.04595279, 0.04628054, 0.04650513, 0.04672294, 
    0.04681281, 0.04689835, 0.04689485, 0.04702025, 0.04709131, 0.04707351, 
    0.04703639, 0.04713644, 0.04736067, 0.04745319, 0.04729952, 0.04723161, 
    0.04717271, 0.04723991, 0.04761359, 0.04794127, 0.04823159, 0.048544, 
    0.04886064, 0.04914401, 0.04944354, 0.04985377, 0.05027255, 0.05069816, 
    0.05099564, 0.05121465, 0.05111641, 0.05070881, 0.05050351, 0.05036645, 
    0.05032397, 0.05026957, 0.05015918, 0.05000679, 0.0500176, 0.05005755, 
    0.05015559, 0.0502746, 0.05012131, 0.05022985, 0.05062416, 0.05091085, 
    0.05110838, 0.05125046, 0.05132223, 0.05144333, 0.05166285, 0.05181509, 
    0.05183036, 0.05169447, 0.05146615, 0.0514281, 0.05176866, 0.0519547, 
    0.05205442, 0.05219254, 0.05253971, 0.05258799, 0.05222629, 0.05206809, 
    0.05205002, 0.05166779, 0.05108884, 0.05088511, 0.0509408, 0.05075757, 
    0.05068621, 0.05069336, 0.05079392, 0.0508125, 0.05077095, 0.05100417, 
    0.05106872, 0.05083298, 0.05024502, 0.04989465, 0.04971255, 0.04988147, 
    0.05058265, 0.05222962, 0.05667794, 0.05934421, 0.06001068, 0.05689058, 
    0.06267077, 0.07235359, 0.06264021, 0.04686175, 0.02917542, 0.02660421, 
    0.02591396, 0.02670359, 0.02673561, 0.02638015, 0.02663511, 0.02824714, 
    0.03037646, 0.03200578, 0.03305751, 0.03381689, 0.03434338, 0.03442495, 
    0.03409918, 0.03356828, 0.03295132, 0.03256457, 0.03249719, 0.03263284, 
    0.03296462, 0.03294633, 0.03258925, 0.03215883, 0.03184995, 0.03138845, 
    0.03083003, 0.03044932, 0.03013561, 0.02980637, 0.02944133, 0.02915079, 
    0.02906273, 0.02890611, 0.0285492, 0.02817084, 0.02775743, 0.02755307, 
    0.02750405, 0.02738317, 0.02721596, 0.02698166, 0.02676796, 0.02651692, 
    0.02626612, 0.02608345, 0.0260159, 0.02589753, 0.02578864, 0.02559492,
  0.02661157, 0.02636885, 0.02625616, 0.02644861, 0.02630585, 0.0259272, 
    0.02556456, 0.02518227, 0.02486245, 0.024753, 0.02485435, 0.02517943, 
    0.02537861, 0.02556192, 0.02576286, 0.02601817, 0.02613569, 0.02631021, 
    0.02654671, 0.02649922, 0.02670619, 0.02698481, 0.02707261, 0.02706606, 
    0.0271196, 0.0272901, 0.02744, 0.02795845, 0.02856408, 0.02926463, 
    0.03013359, 0.03049657, 0.03059467, 0.03097324, 0.03163278, 0.03234109, 
    0.03349822, 0.03388016, 0.03363077, 0.03337897, 0.03114286, 0.02426338, 
    0.02876302, 0.03639114, 0.03112443, 0.02789784, 0.02658114, 0.02673004, 
    0.02562773, 0.02463689, 0.02394115, 0.02363005, 0.0235373, 0.02382327, 
    0.02386686, 0.02376748, 0.02345298, 0.02299245, 0.02287332, 0.02290039, 
    0.02293129, 0.02317915, 0.02376548, 0.02422815, 0.0250597, 0.02551123, 
    0.02621276, 0.02647377, 0.02651395, 0.02620235, 0.02550461, 0.02435193, 
    0.02322806, 0.02246442, 0.02178376, 0.02227117, 0.02231009, 0.02289155, 
    0.02219241, 0.02047387, 0.01924734, 0.01660188, 0.01708635, 0.02026712, 
    0.02064048, 0.02402172, 0.02399559, 0.02192397, 0.02077822, 0.021274, 
    0.02251117, 0.02980508, 0.03183659, 0.03131123, 0.0311116, 0.03260417, 
    0.03445501, 0.0350471, 0.0333014, 0.03580736, 0.0374884, 0.03745671, 
    0.03821972, 0.03693802, 0.03683025, 0.03810652, 0.03476718, 0.03577445, 
    0.0375951, 0.03766236, 0.03710888, 0.03677298, 0.03769056, 0.03733607, 
    0.03722687, 0.03624135, 0.03626996, 0.0350881, 0.03440641, 0.03350054, 
    0.03403607, 0.03496018, 0.03598542, 0.03720587, 0.03811894, 0.0388229, 
    0.03941056, 0.03999124, 0.04068378, 0.04152657, 0.04215736, 0.04302333, 
    0.04417636, 0.04534218, 0.04643548, 0.04734096, 0.04811682, 0.04864151, 
    0.04885805, 0.04918422, 0.04953385, 0.05008694, 0.05080637, 0.05197627, 
    0.05274191, 0.05346596, 0.0536674, 0.05376843, 0.05352474, 0.05338793, 
    0.05317575, 0.05308778, 0.05298145, 0.05305073, 0.05291136, 0.0528575, 
    0.0526947, 0.05263204, 0.05266162, 0.05291089, 0.05283788, 0.05263324, 
    0.05244281, 0.05256536, 0.05278116, 0.05302028, 0.05326086, 0.05347852, 
    0.05367208, 0.05382026, 0.05392791, 0.05416363, 0.05447978, 0.05492286, 
    0.05562681, 0.05570986, 0.05551624, 0.0552404, 0.05493687, 0.0545831, 
    0.05448014, 0.05465535, 0.05484207, 0.05501157, 0.0552075, 0.05537745, 
    0.05584686, 0.05648701, 0.05694685, 0.05736879, 0.05745769, 0.05716386, 
    0.05704284, 0.05715429, 0.05724664, 0.05713746, 0.05706625, 0.05715469, 
    0.05689485, 0.05638349, 0.0558619, 0.05537274, 0.05521924, 0.05526762, 
    0.05522996, 0.05527252, 0.05553444, 0.0555566, 0.05524145, 0.05501342, 
    0.05467001, 0.05446078, 0.05424713, 0.05409795, 0.05407112, 0.05394936, 
    0.05396427, 0.05423044, 0.05446135, 0.05467093, 0.0548796, 0.05512691, 
    0.05521866, 0.05516157, 0.05516132, 0.05500526, 0.05481598, 0.05449628, 
    0.05462551, 0.05481296, 0.05628188, 0.05999019, 0.06367159, 0.06489383, 
    0.06496567, 0.06889486, 0.07792825, 0.07492945, 0.04753998, 0.03371962, 
    0.02785003, 0.02663079, 0.02744526, 0.03047673, 0.03197113, 0.03220204, 
    0.03297586, 0.0345811, 0.03641517, 0.03766133, 0.03827805, 0.03835458, 
    0.03801613, 0.03759494, 0.03701942, 0.03648471, 0.03628969, 0.03627635, 
    0.0361627, 0.03604331, 0.03571225, 0.03511059, 0.03457523, 0.03397587, 
    0.03349078, 0.03331383, 0.0330285, 0.03247651, 0.03205983, 0.03167481, 
    0.03137641, 0.03108748, 0.03060981, 0.03010946, 0.02988637, 0.02986084, 
    0.02995934, 0.02994775, 0.029678, 0.02936232, 0.02883577, 0.02850973, 
    0.02823888, 0.02790319, 0.02762436, 0.02752929, 0.0273755, 0.02696359,
  0.0282136, 0.02780632, 0.02762229, 0.02749768, 0.0272418, 0.0270511, 
    0.02693482, 0.0268093, 0.02652387, 0.02636122, 0.02635907, 0.02658187, 
    0.02683088, 0.02700156, 0.02717367, 0.0274665, 0.02772539, 0.02778169, 
    0.02764319, 0.02769501, 0.02791851, 0.02827165, 0.02845683, 0.02860052, 
    0.02887086, 0.0291471, 0.02931942, 0.02946518, 0.02977505, 0.03042693, 
    0.03144998, 0.03242496, 0.03283837, 0.03268775, 0.03291954, 0.03341903, 
    0.03435963, 0.03533552, 0.03646927, 0.03733768, 0.03944233, 0.03999969, 
    0.03979677, 0.03808955, 0.03523117, 0.03476478, 0.03285393, 0.03146069, 
    0.03041469, 0.02991831, 0.02958938, 0.02929027, 0.02896256, 0.0287291, 
    0.02850811, 0.02793209, 0.02750758, 0.02698706, 0.0267715, 0.02670044, 
    0.02666908, 0.02674115, 0.02676706, 0.02699888, 0.02755947, 0.0278146, 
    0.02798562, 0.02815158, 0.02839642, 0.02887601, 0.02918425, 0.02952396, 
    0.0295528, 0.0293987, 0.02902156, 0.0284147, 0.02819159, 0.02821846, 
    0.0282862, 0.02846857, 0.02929701, 0.03014799, 0.03082041, 0.03020674, 
    0.02958498, 0.0304456, 0.03003628, 0.03011905, 0.03100259, 0.03218412, 
    0.03368725, 0.03500056, 0.03464242, 0.03416006, 0.03518699, 0.03616364, 
    0.03715301, 0.03867538, 0.03983494, 0.04127595, 0.0422006, 0.0430281, 
    0.04487474, 0.04661885, 0.04776249, 0.04915718, 0.0508181, 0.05129344, 
    0.05117454, 0.05046671, 0.05101147, 0.05052134, 0.0499375, 0.04933666, 
    0.0490966, 0.04828966, 0.04675463, 0.04552139, 0.04422993, 0.0438, 
    0.04384176, 0.0441086, 0.04458851, 0.04522333, 0.04586758, 0.04628596, 
    0.04669324, 0.04710632, 0.04767473, 0.04821146, 0.04883178, 0.04952024, 
    0.05035898, 0.05128893, 0.05225306, 0.05308125, 0.05362639, 0.054294, 
    0.05498012, 0.05561702, 0.05634868, 0.0575383, 0.05857147, 0.06005984, 
    0.06079252, 0.06128361, 0.06148818, 0.06154497, 0.06105441, 0.06052876, 
    0.0603388, 0.06025317, 0.06030758, 0.06014396, 0.05988215, 0.05953711, 
    0.05920334, 0.0589897, 0.05895039, 0.05894561, 0.05897135, 0.05897791, 
    0.05900888, 0.05894902, 0.05902168, 0.05905557, 0.05875687, 0.05858248, 
    0.05849917, 0.05848943, 0.05846529, 0.05858393, 0.05870779, 0.0587548, 
    0.05893852, 0.05919763, 0.05946166, 0.0595315, 0.05942135, 0.05911386, 
    0.05899213, 0.05925443, 0.0597579, 0.06017888, 0.06048282, 0.06074068, 
    0.06096024, 0.06115621, 0.06153327, 0.06170112, 0.06168634, 0.06149989, 
    0.06125574, 0.06120741, 0.06127618, 0.0609119, 0.06041057, 0.06021943, 
    0.05976736, 0.05909619, 0.05837765, 0.05762149, 0.0572643, 0.0572171, 
    0.05706204, 0.05701314, 0.05713756, 0.05717674, 0.0568962, 0.05688617, 
    0.0569346, 0.05682712, 0.056752, 0.05686115, 0.05691181, 0.05694506, 
    0.05698198, 0.05719689, 0.0573597, 0.0575566, 0.05771933, 0.0580166, 
    0.0584185, 0.05874874, 0.0591998, 0.05941488, 0.05928766, 0.05918839, 
    0.05906539, 0.05919643, 0.05887094, 0.05986441, 0.06227725, 0.06557075, 
    0.06867506, 0.06788009, 0.06901586, 0.07091996, 0.06191879, 0.04875877, 
    0.04229396, 0.04338678, 0.03443348, 0.03045706, 0.0327531, 0.03630191, 
    0.03763905, 0.0388302, 0.04021199, 0.04150326, 0.04203889, 0.0421801, 
    0.04193787, 0.04152758, 0.04101151, 0.04056082, 0.04017621, 0.03988594, 
    0.03961489, 0.03943725, 0.03920224, 0.03875528, 0.03809093, 0.03739308, 
    0.03682872, 0.03644532, 0.0359687, 0.0355526, 0.03515725, 0.03466772, 
    0.03420613, 0.0337084, 0.03321181, 0.03266083, 0.03230567, 0.03211625, 
    0.03193385, 0.03172856, 0.03146138, 0.03115473, 0.03087347, 0.03045649, 
    0.02998253, 0.0295517, 0.02922929, 0.02919924, 0.02901921, 0.02860826,
  0.03004768, 0.02977649, 0.02948399, 0.0291842, 0.02888671, 0.02869569, 
    0.02863357, 0.02868224, 0.02868352, 0.02860366, 0.02862099, 0.0287213, 
    0.02883603, 0.02888243, 0.02896863, 0.02918915, 0.0295125, 0.02952248, 
    0.02962118, 0.02981724, 0.03000789, 0.03031866, 0.03069593, 0.03123947, 
    0.03163148, 0.03162295, 0.03197158, 0.0321773, 0.03244429, 0.03283654, 
    0.03319855, 0.03347022, 0.03378825, 0.03410731, 0.03426973, 0.03454455, 
    0.03522262, 0.03598194, 0.03655491, 0.03712607, 0.03769156, 0.03807658, 
    0.03807149, 0.03808618, 0.03720004, 0.0362964, 0.03554986, 0.0350913, 
    0.0348124, 0.03417179, 0.03346569, 0.03284089, 0.03266299, 0.03239711, 
    0.03212499, 0.03179606, 0.03153952, 0.03120363, 0.03091392, 0.03070395, 
    0.03054118, 0.03046945, 0.03039933, 0.03049599, 0.03074938, 0.03062063, 
    0.03025295, 0.03029118, 0.03041015, 0.03058216, 0.0307573, 0.03086473, 
    0.03083736, 0.03082324, 0.03101094, 0.03115005, 0.03148226, 0.03164685, 
    0.03183453, 0.03228259, 0.03265344, 0.03270256, 0.03287973, 0.0328338, 
    0.03299636, 0.03393757, 0.03465146, 0.0353179, 0.03613294, 0.03636622, 
    0.03687353, 0.03714569, 0.0375589, 0.0385437, 0.03942405, 0.04023542, 
    0.04105307, 0.04182578, 0.04317867, 0.04445289, 0.04546411, 0.04636465, 
    0.04767362, 0.04878615, 0.04990023, 0.05090304, 0.05162938, 0.05254064, 
    0.05339463, 0.05448731, 0.05483022, 0.05481948, 0.05492292, 0.05509447, 
    0.05472282, 0.05417257, 0.05326346, 0.05257897, 0.05232968, 0.05231324, 
    0.05236307, 0.05254881, 0.05282653, 0.05321343, 0.05374483, 0.05403639, 
    0.05418792, 0.05442095, 0.05474434, 0.0550224, 0.05552555, 0.05616898, 
    0.05705846, 0.05808109, 0.05913964, 0.05997429, 0.06051478, 0.0612509, 
    0.06209283, 0.06277958, 0.06341869, 0.06414841, 0.0647343, 0.06514908, 
    0.06523892, 0.06512432, 0.06476633, 0.06445133, 0.06427474, 0.06435881, 
    0.06457869, 0.06485542, 0.06510164, 0.06494235, 0.06492333, 0.06484827, 
    0.06498774, 0.06501214, 0.06493501, 0.06488954, 0.06483549, 0.06488307, 
    0.06476395, 0.06459511, 0.06439295, 0.06392301, 0.06355381, 0.06321755, 
    0.06293187, 0.06272335, 0.06268089, 0.06277557, 0.0628416, 0.06294351, 
    0.06321099, 0.06352504, 0.06378023, 0.06374962, 0.06353799, 0.0634557, 
    0.06355157, 0.06381805, 0.06417804, 0.06457193, 0.06460152, 0.06443907, 
    0.064281, 0.06424714, 0.06440453, 0.06488383, 0.0650409, 0.06497959, 
    0.06479173, 0.06447487, 0.06414276, 0.06365859, 0.06325006, 0.06263682, 
    0.06190101, 0.06111388, 0.0601953, 0.05941235, 0.05891697, 0.05878677, 
    0.05849482, 0.05822832, 0.05832723, 0.0584477, 0.05848588, 0.05874433, 
    0.05912542, 0.05910574, 0.05914267, 0.05947511, 0.05966026, 0.05981312, 
    0.05977206, 0.05992145, 0.06022506, 0.06042319, 0.06041244, 0.06079002, 
    0.06132586, 0.06191397, 0.0624638, 0.06292516, 0.06306072, 0.06287124, 
    0.06288373, 0.06326617, 0.06351823, 0.06317499, 0.06270726, 0.06287279, 
    0.06485251, 0.06805462, 0.06976365, 0.07016957, 0.06882269, 0.06305926, 
    0.05644709, 0.0522248, 0.04337317, 0.04029644, 0.03999258, 0.04071057, 
    0.04268883, 0.0443834, 0.04541627, 0.04601141, 0.04627912, 0.04633232, 
    0.04589136, 0.04527446, 0.04476023, 0.04440464, 0.04396849, 0.04371154, 
    0.043458, 0.04324554, 0.04287307, 0.04221876, 0.04161479, 0.04098244, 
    0.04039123, 0.03977275, 0.03930392, 0.03894189, 0.03848751, 0.03798459, 
    0.03741304, 0.03688757, 0.03641497, 0.03571691, 0.03511284, 0.03461156, 
    0.03428109, 0.03406297, 0.03376782, 0.03346798, 0.03333861, 0.03280259, 
    0.03208329, 0.03167066, 0.0312761, 0.03090419, 0.03057409, 0.0302809,
  0.0321713, 0.03188181, 0.03149214, 0.03099914, 0.03057847, 0.03046429, 
    0.03065856, 0.03098101, 0.03109451, 0.03112669, 0.03125647, 0.03133642, 
    0.03143688, 0.03168486, 0.03188398, 0.03193492, 0.03220379, 0.03251271, 
    0.03284205, 0.03285672, 0.03326717, 0.03368051, 0.03397885, 0.03400969, 
    0.03406851, 0.03419328, 0.03437713, 0.03481255, 0.03521161, 0.03545517, 
    0.03575593, 0.03595366, 0.03574612, 0.03562026, 0.03594274, 0.03647953, 
    0.03702494, 0.03739673, 0.03776152, 0.03814183, 0.03840014, 0.03871132, 
    0.03856513, 0.03855324, 0.03860791, 0.03875301, 0.03902849, 0.03909883, 
    0.03916702, 0.03873338, 0.03844684, 0.03841064, 0.03795565, 0.03724968, 
    0.03659081, 0.03611736, 0.035778, 0.0354433, 0.0351701, 0.03475654, 
    0.03443776, 0.03424858, 0.034185, 0.03422865, 0.03455925, 0.03432432, 
    0.03390817, 0.03339018, 0.0333581, 0.03359597, 0.03390022, 0.03409809, 
    0.03411854, 0.03418111, 0.03436253, 0.03453359, 0.03476714, 0.03483723, 
    0.03525316, 0.03584092, 0.0363006, 0.03645426, 0.03655045, 0.03656171, 
    0.03704603, 0.03777701, 0.03870777, 0.03930508, 0.03981319, 0.04030036, 
    0.04066227, 0.04099184, 0.04160266, 0.04191834, 0.04238575, 0.04313939, 
    0.04394875, 0.0447249, 0.0458461, 0.04701851, 0.04805891, 0.04886487, 
    0.04954926, 0.05067784, 0.05136604, 0.05220296, 0.05294529, 0.05360327, 
    0.05477272, 0.05555474, 0.05604552, 0.05679866, 0.05784554, 0.05822983, 
    0.05824046, 0.0585321, 0.05902162, 0.0593783, 0.05943376, 0.05949444, 
    0.0597329, 0.05986403, 0.06001756, 0.06030256, 0.06067786, 0.06102739, 
    0.06122276, 0.06144759, 0.06177736, 0.06217592, 0.06267332, 0.06360685, 
    0.06442913, 0.06516451, 0.06568436, 0.06617156, 0.06662417, 0.06715319, 
    0.06766331, 0.06818514, 0.06855705, 0.06870454, 0.06882339, 0.06872837, 
    0.06834464, 0.06804103, 0.06770605, 0.06718391, 0.06687615, 0.06707576, 
    0.06722982, 0.06740133, 0.06761611, 0.06792294, 0.06844827, 0.06891064, 
    0.06947111, 0.06968826, 0.06944168, 0.06939582, 0.06945658, 0.06963971, 
    0.06957401, 0.06915425, 0.06875481, 0.06835631, 0.06795081, 0.06755866, 
    0.06715335, 0.06682497, 0.06654466, 0.06676031, 0.06715079, 0.06749193, 
    0.06799857, 0.0682875, 0.0683011, 0.0679843, 0.06760515, 0.06744201, 
    0.06748352, 0.06755607, 0.06793836, 0.06800345, 0.06775267, 0.06752793, 
    0.06741859, 0.0675241, 0.0675768, 0.0678007, 0.06815112, 0.0681025, 
    0.0678262, 0.06749149, 0.06712057, 0.06667491, 0.06606104, 0.06519894, 
    0.06443939, 0.06356356, 0.06255858, 0.06177042, 0.06120466, 0.06083416, 
    0.06056806, 0.06046164, 0.06058477, 0.06082274, 0.06087963, 0.06105336, 
    0.06121204, 0.06123861, 0.06134579, 0.06156162, 0.06166949, 0.06175533, 
    0.06176925, 0.062109, 0.06265734, 0.06298451, 0.06323831, 0.06346951, 
    0.06383019, 0.06436648, 0.06518725, 0.06564632, 0.06570479, 0.06565317, 
    0.06554896, 0.06542478, 0.06528844, 0.06584544, 0.06618007, 0.06648779, 
    0.0667709, 0.06758608, 0.06898461, 0.06895547, 0.0684789, 0.06687219, 
    0.06292833, 0.05720223, 0.05395538, 0.05182242, 0.05020486, 0.04955336, 
    0.04989043, 0.05061683, 0.05111885, 0.05136164, 0.05134961, 0.05127757, 
    0.05099616, 0.05028423, 0.04962934, 0.04893072, 0.04839566, 0.04803018, 
    0.04775334, 0.04740777, 0.04718391, 0.04675449, 0.04603552, 0.04515182, 
    0.04406887, 0.04328493, 0.04286446, 0.04283305, 0.04239875, 0.04174386, 
    0.04097826, 0.04028095, 0.0397028, 0.03913802, 0.03865868, 0.03802957, 
    0.03743804, 0.03683316, 0.03636022, 0.03590521, 0.03544208, 0.03518154, 
    0.03496545, 0.03433491, 0.03372294, 0.03308908, 0.03257872, 0.03222466,
  0.03454265, 0.03423082, 0.03398146, 0.03386149, 0.0336027, 0.03350994, 
    0.03379046, 0.0338089, 0.03380091, 0.03389698, 0.03404218, 0.03411164, 
    0.03432398, 0.03471295, 0.03475368, 0.03471481, 0.03475812, 0.03504164, 
    0.03551456, 0.03585947, 0.03652541, 0.0370978, 0.03713538, 0.03703576, 
    0.0373471, 0.03750194, 0.037583, 0.03790864, 0.03831671, 0.03873501, 
    0.03911807, 0.03906832, 0.03896382, 0.03878136, 0.03885297, 0.03925269, 
    0.03961332, 0.03979517, 0.04015787, 0.04052026, 0.04080971, 0.04095051, 
    0.0411365, 0.0413892, 0.04164548, 0.0417511, 0.04214058, 0.04241736, 
    0.04275236, 0.04277344, 0.04285993, 0.04282573, 0.04263565, 0.04208964, 
    0.04160259, 0.04117727, 0.04054453, 0.03990926, 0.03915632, 0.03862633, 
    0.03818949, 0.03773519, 0.03748251, 0.03727594, 0.03701517, 0.03693707, 
    0.03690817, 0.03674878, 0.037096, 0.03769025, 0.0383774, 0.03863849, 
    0.03867099, 0.03859116, 0.03852724, 0.03847835, 0.03881837, 0.03920666, 
    0.03953161, 0.0397032, 0.03988779, 0.03975753, 0.03964875, 0.03977337, 
    0.0401613, 0.04075597, 0.04160891, 0.04243477, 0.04312058, 0.04384363, 
    0.04413361, 0.0444686, 0.04473353, 0.04489278, 0.04501662, 0.04539698, 
    0.04623022, 0.04712555, 0.04822697, 0.04944035, 0.05035366, 0.05097323, 
    0.05169793, 0.05268477, 0.05343879, 0.0542603, 0.0552507, 0.0561876, 
    0.05709744, 0.05816726, 0.05950501, 0.0604789, 0.06134077, 0.06195252, 
    0.06235715, 0.06274747, 0.06303322, 0.06339296, 0.06386378, 0.06460586, 
    0.06546132, 0.06602598, 0.06649181, 0.06681313, 0.06709539, 0.06745001, 
    0.06757743, 0.06771562, 0.06806953, 0.06851415, 0.06905662, 0.06958643, 
    0.06990662, 0.06975531, 0.07002896, 0.07044686, 0.07086833, 0.07130775, 
    0.07158072, 0.07142394, 0.0716413, 0.07187047, 0.07140064, 0.07116135, 
    0.07090231, 0.07069447, 0.0704525, 0.07025924, 0.07022265, 0.07033284, 
    0.07059861, 0.07076242, 0.07098583, 0.07150064, 0.07202663, 0.07235134, 
    0.07280208, 0.07320717, 0.07338206, 0.07323789, 0.07307339, 0.0731245, 
    0.07312777, 0.07317145, 0.07324026, 0.07296354, 0.07245678, 0.07207625, 
    0.07169686, 0.07150093, 0.07130025, 0.07132515, 0.07158486, 0.07202239, 
    0.07232621, 0.0722992, 0.07192682, 0.07160139, 0.07147074, 0.07142269, 
    0.07157279, 0.07176322, 0.07163936, 0.07125632, 0.07089955, 0.07084102, 
    0.07096385, 0.07108795, 0.07099892, 0.07108513, 0.07105417, 0.07092062, 
    0.0707265, 0.07048272, 0.06992377, 0.069401, 0.06877855, 0.06770471, 
    0.06687097, 0.06617103, 0.06531813, 0.06450507, 0.06377162, 0.06343914, 
    0.06319319, 0.06271392, 0.06277952, 0.06306276, 0.06361129, 0.06359074, 
    0.06345758, 0.06363223, 0.06368672, 0.06373258, 0.06382364, 0.06386245, 
    0.06398503, 0.06460306, 0.06511065, 0.06550373, 0.0658544, 0.066037, 
    0.06615181, 0.06661721, 0.06738055, 0.06763576, 0.06767426, 0.06749685, 
    0.06762259, 0.06765672, 0.06809366, 0.06855014, 0.06874563, 0.06875528, 
    0.06890777, 0.06900942, 0.06929373, 0.06925418, 0.06863914, 0.06739178, 
    0.06637482, 0.06448451, 0.06217531, 0.05998851, 0.05892765, 0.05821124, 
    0.05739503, 0.05729897, 0.05711105, 0.05716031, 0.05723928, 0.0572053, 
    0.05657799, 0.05550711, 0.05500817, 0.0542099, 0.05344628, 0.05307453, 
    0.05266519, 0.05197578, 0.05140665, 0.0507092, 0.05001444, 0.04912614, 
    0.04791522, 0.04710724, 0.04658544, 0.0464335, 0.04621597, 0.04572408, 
    0.04507176, 0.04435667, 0.04354593, 0.04286818, 0.04243356, 0.04161656, 
    0.04086371, 0.04037502, 0.03987113, 0.03930686, 0.03852613, 0.0379416, 
    0.0373762, 0.03682196, 0.03622298, 0.03566946, 0.0352947, 0.0349003,
  0.03804304, 0.03742401, 0.0370651, 0.03690138, 0.03672415, 0.03679544, 
    0.03701461, 0.03698304, 0.0368804, 0.03683157, 0.03694504, 0.03711885, 
    0.03736461, 0.03748402, 0.03766175, 0.03769658, 0.03796828, 0.03873657, 
    0.03945269, 0.03988828, 0.04043823, 0.04124083, 0.04112763, 0.04089873, 
    0.04080807, 0.04074946, 0.04096385, 0.04145669, 0.04211837, 0.04271647, 
    0.04301239, 0.0431533, 0.0433948, 0.04304988, 0.04292647, 0.04301224, 
    0.04327742, 0.04356101, 0.04391591, 0.04422313, 0.04463364, 0.04480791, 
    0.04513229, 0.04531178, 0.04561678, 0.04604904, 0.04656109, 0.04680054, 
    0.04705026, 0.04679394, 0.04698645, 0.04730386, 0.04733118, 0.04698883, 
    0.04641545, 0.04572592, 0.04513925, 0.04471165, 0.04389476, 0.04336369, 
    0.04300435, 0.04253823, 0.04208874, 0.04156515, 0.04080721, 0.04067596, 
    0.04075441, 0.04073365, 0.04176406, 0.04276173, 0.0432681, 0.04333399, 
    0.04321009, 0.04303782, 0.04298947, 0.0430285, 0.04319805, 0.04313588, 
    0.04323282, 0.04357865, 0.04360349, 0.04350544, 0.04366786, 0.04357556, 
    0.04337215, 0.04362718, 0.04403334, 0.04484391, 0.0455036, 0.0461563, 
    0.0465145, 0.04662334, 0.04685605, 0.04717762, 0.04745653, 0.04779572, 
    0.04848086, 0.04939927, 0.05034859, 0.05137279, 0.05214084, 0.0527276, 
    0.05361392, 0.05468139, 0.0556135, 0.05644172, 0.05753757, 0.05886682, 
    0.06008178, 0.06127164, 0.0625662, 0.06366098, 0.06444879, 0.06491653, 
    0.06532203, 0.06570669, 0.06607872, 0.0666505, 0.06754757, 0.0686939, 
    0.06956228, 0.07013239, 0.07060004, 0.07108226, 0.07140189, 0.0716489, 
    0.07195798, 0.07222632, 0.07268346, 0.07324185, 0.07340546, 0.07359225, 
    0.07363299, 0.07317167, 0.07319608, 0.07351584, 0.07413971, 0.07453872, 
    0.07455256, 0.0741789, 0.07367184, 0.07338757, 0.07329897, 0.07328393, 
    0.07314047, 0.07283886, 0.07273644, 0.07289321, 0.07318913, 0.07338027, 
    0.07367792, 0.07407543, 0.07461215, 0.07517239, 0.07533038, 0.07549812, 
    0.07580248, 0.07632191, 0.07660908, 0.0764365, 0.07628909, 0.07621838, 
    0.07667269, 0.07747933, 0.07794718, 0.07793071, 0.07742289, 0.07728964, 
    0.07686888, 0.07654922, 0.07620319, 0.07594299, 0.07586145, 0.07584605, 
    0.07578507, 0.07579411, 0.07544772, 0.07527171, 0.075297, 0.07542803, 
    0.07559125, 0.07577799, 0.07551306, 0.07483034, 0.07450905, 0.07454892, 
    0.07482185, 0.07494663, 0.07491787, 0.07471037, 0.07413772, 0.07360316, 
    0.07306932, 0.07264394, 0.07185932, 0.07101759, 0.07030987, 0.06945942, 
    0.06872828, 0.06802829, 0.06709869, 0.06622498, 0.06573926, 0.06549429, 
    0.06536016, 0.06507309, 0.06487647, 0.0649252, 0.065431, 0.06555772, 
    0.06558614, 0.06570924, 0.06570154, 0.0658049, 0.06621215, 0.06622984, 
    0.06631827, 0.06670593, 0.06689013, 0.067318, 0.06804023, 0.06814367, 
    0.06803153, 0.06798156, 0.0683377, 0.06855209, 0.06846379, 0.06865131, 
    0.06922374, 0.06981622, 0.07053194, 0.0709556, 0.07114575, 0.07104535, 
    0.07088187, 0.07078777, 0.07078841, 0.07086729, 0.07078031, 0.07020635, 
    0.06884669, 0.06769348, 0.06675801, 0.06583591, 0.06515341, 0.06462964, 
    0.06390324, 0.06344246, 0.06314407, 0.06266377, 0.06229036, 0.06230177, 
    0.06138078, 0.06043986, 0.06016591, 0.0596909, 0.05878086, 0.05767223, 
    0.05729467, 0.05670886, 0.05604247, 0.05527755, 0.05439051, 0.0534327, 
    0.05253805, 0.05170833, 0.05132761, 0.05117302, 0.05101477, 0.05075694, 
    0.05004709, 0.0491364, 0.04812686, 0.04715541, 0.04638002, 0.04569941, 
    0.04512516, 0.04456497, 0.04368536, 0.04277227, 0.04203692, 0.0414518, 
    0.04082381, 0.04004335, 0.03950432, 0.03909428, 0.03884629, 0.03852405,
  0.04192535, 0.04137741, 0.0410756, 0.04076833, 0.04054682, 0.04023853, 
    0.04034231, 0.04038403, 0.04021258, 0.04016866, 0.0402522, 0.04033208, 
    0.04044999, 0.04037668, 0.04067479, 0.04129538, 0.04220284, 0.04325673, 
    0.04438708, 0.04543258, 0.04616658, 0.04622256, 0.04584383, 0.04538612, 
    0.04496576, 0.04498369, 0.04529637, 0.04591251, 0.0466914, 0.04712584, 
    0.04728626, 0.04752605, 0.04757085, 0.0474694, 0.04746151, 0.04748994, 
    0.04757566, 0.04757547, 0.04779377, 0.04812397, 0.04862216, 0.04908158, 
    0.04955081, 0.04956046, 0.04977725, 0.0502341, 0.0508546, 0.05137787, 
    0.05181499, 0.05194798, 0.05206585, 0.05222719, 0.0520012, 0.05167202, 
    0.05146417, 0.05078819, 0.04992525, 0.04919192, 0.04847762, 0.04801961, 
    0.04795017, 0.04777145, 0.04738793, 0.04684557, 0.04618293, 0.04588047, 
    0.0458678, 0.04625244, 0.04723144, 0.04783324, 0.04790273, 0.04751648, 
    0.04719716, 0.04689822, 0.04665574, 0.04684456, 0.04700541, 0.04657385, 
    0.04645832, 0.04654764, 0.04661376, 0.04667945, 0.04671501, 0.04688641, 
    0.04703424, 0.04738382, 0.04737994, 0.04767051, 0.048305, 0.0488169, 
    0.04905622, 0.0491731, 0.0494458, 0.04965826, 0.04979185, 0.05017332, 
    0.05089316, 0.05176155, 0.05264045, 0.0534256, 0.05409556, 0.05493803, 
    0.05598996, 0.05689472, 0.05786118, 0.05906007, 0.0602461, 0.06161423, 
    0.0629014, 0.06432387, 0.06557004, 0.06663901, 0.06728388, 0.06773487, 
    0.06821432, 0.06870976, 0.06934066, 0.07007179, 0.07110272, 0.07216783, 
    0.07319744, 0.07387489, 0.07434718, 0.07506847, 0.07526194, 0.07532202, 
    0.07562566, 0.07601508, 0.07644718, 0.07657588, 0.07683592, 0.07698666, 
    0.07698285, 0.07683054, 0.07687832, 0.07718509, 0.07784899, 0.07782144, 
    0.07721782, 0.07611195, 0.07500025, 0.07447761, 0.07456389, 0.07473589, 
    0.07470131, 0.07461599, 0.07472727, 0.07519562, 0.07568437, 0.07577014, 
    0.07607419, 0.07658307, 0.07732841, 0.07812426, 0.07877626, 0.07908206, 
    0.07930385, 0.07973256, 0.07978582, 0.07960805, 0.07942312, 0.07979049, 
    0.08060174, 0.08132115, 0.08190213, 0.08196346, 0.08163561, 0.0813506, 
    0.0813072, 0.08108528, 0.08058624, 0.08008573, 0.07975788, 0.0795705, 
    0.07953431, 0.07956851, 0.07945707, 0.0793689, 0.07946437, 0.07950891, 
    0.07938002, 0.07935324, 0.07908559, 0.07880829, 0.07858565, 0.07865295, 
    0.07896238, 0.07900869, 0.07872115, 0.07790162, 0.07696028, 0.07599033, 
    0.07502259, 0.07410301, 0.0731569, 0.07257185, 0.07179642, 0.071137, 
    0.07096196, 0.07016298, 0.06917135, 0.06851249, 0.06807762, 0.06777257, 
    0.06754664, 0.0673086, 0.06732306, 0.06757368, 0.06792516, 0.06791894, 
    0.06788676, 0.06797948, 0.06786764, 0.06786208, 0.06800824, 0.06815205, 
    0.06818437, 0.06819587, 0.06807838, 0.06868548, 0.06927547, 0.0692375, 
    0.06891473, 0.06873348, 0.06900457, 0.06930525, 0.06949504, 0.06985664, 
    0.07036558, 0.07074717, 0.07126838, 0.07146756, 0.07121964, 0.07133168, 
    0.07133132, 0.07102118, 0.07079922, 0.0709257, 0.07112642, 0.07082589, 
    0.07053541, 0.0701445, 0.06971724, 0.06921573, 0.06868662, 0.06831164, 
    0.06800386, 0.06779645, 0.06740031, 0.06700161, 0.06682085, 0.06664017, 
    0.06609836, 0.06602528, 0.06606279, 0.06561773, 0.06472514, 0.06392868, 
    0.06314304, 0.06212947, 0.06113055, 0.0602881, 0.05953354, 0.05868088, 
    0.05770938, 0.05685599, 0.05624513, 0.05575117, 0.05588009, 0.05595255, 
    0.05508592, 0.05399831, 0.05283216, 0.05179975, 0.05072517, 0.04989979, 
    0.04932703, 0.0485314, 0.04771719, 0.04700163, 0.04662677, 0.04602889, 
    0.04533372, 0.04454624, 0.04383454, 0.04323443, 0.04271331, 0.04246036,
  0.04622063, 0.04582854, 0.0454906, 0.04496928, 0.04421761, 0.04373695, 
    0.0435851, 0.04365724, 0.04378429, 0.0439101, 0.04411439, 0.04444126, 
    0.04479485, 0.04499601, 0.04534243, 0.04617613, 0.04706084, 0.04805342, 
    0.04921794, 0.05021411, 0.05097008, 0.05087816, 0.05057748, 0.05034653, 
    0.0502113, 0.05007299, 0.05027249, 0.05048389, 0.05077055, 0.05118341, 
    0.05147157, 0.05148965, 0.05124446, 0.0511424, 0.05115011, 0.05108467, 
    0.05123988, 0.05121876, 0.05153633, 0.05161129, 0.0519872, 0.05244878, 
    0.05291903, 0.05334803, 0.0534999, 0.05402167, 0.05488531, 0.05542019, 
    0.05578236, 0.05596539, 0.05587437, 0.05576723, 0.05555925, 0.05543484, 
    0.05554323, 0.05533788, 0.05459944, 0.05387998, 0.05310078, 0.05244778, 
    0.05218395, 0.05211979, 0.0521287, 0.05203538, 0.05168188, 0.05126588, 
    0.05111477, 0.05122399, 0.05123634, 0.05108786, 0.05079253, 0.05055479, 
    0.05010392, 0.04984342, 0.04973444, 0.04987773, 0.04995361, 0.05002646, 
    0.04974598, 0.04963214, 0.04946898, 0.04952817, 0.04989772, 0.0501332, 
    0.05022014, 0.05016281, 0.05014761, 0.05056071, 0.0510579, 0.05157726, 
    0.05183604, 0.0521365, 0.05250075, 0.0529477, 0.05320909, 0.05359781, 
    0.0540508, 0.05483779, 0.0557987, 0.05653816, 0.05726226, 0.05810845, 
    0.05900862, 0.06007407, 0.06122825, 0.06245966, 0.06392868, 0.0651223, 
    0.06604303, 0.06710936, 0.06824283, 0.06954222, 0.07037533, 0.07078745, 
    0.0711809, 0.07160819, 0.07234996, 0.07328033, 0.07442119, 0.07576153, 
    0.07693288, 0.07756614, 0.07790485, 0.07834715, 0.07876921, 0.078892, 
    0.07916807, 0.07959821, 0.08018632, 0.08063292, 0.08089042, 0.08101778, 
    0.08107043, 0.0809069, 0.08093001, 0.08109514, 0.08113437, 0.08040288, 
    0.07911154, 0.07768238, 0.07676136, 0.07615033, 0.07592538, 0.07596354, 
    0.07598857, 0.07615103, 0.07643589, 0.07676519, 0.07696845, 0.0772284, 
    0.07777509, 0.07854991, 0.07953259, 0.08049123, 0.08105835, 0.08147201, 
    0.08171172, 0.08182207, 0.08193486, 0.0824443, 0.08280254, 0.08342649, 
    0.08389085, 0.08422067, 0.08453244, 0.08489847, 0.08492304, 0.08474579, 
    0.08443492, 0.08419997, 0.08387316, 0.08339459, 0.08309496, 0.08316281, 
    0.08331851, 0.0833686, 0.08325203, 0.08312874, 0.08293013, 0.08271218, 
    0.08294129, 0.08324356, 0.08366841, 0.08358316, 0.08322798, 0.08269602, 
    0.08274869, 0.08269735, 0.08192393, 0.08075014, 0.07942277, 0.07814436, 
    0.07711667, 0.07643122, 0.07560398, 0.07495434, 0.07438269, 0.07387569, 
    0.07350563, 0.07269397, 0.07138619, 0.07093831, 0.07047389, 0.07009135, 
    0.06997238, 0.06974076, 0.06974612, 0.06988801, 0.06993968, 0.06976936, 
    0.06964253, 0.06965675, 0.06971432, 0.06966082, 0.06961404, 0.06966413, 
    0.06964652, 0.06964412, 0.06965702, 0.06988205, 0.07005795, 0.07005296, 
    0.07005104, 0.07016114, 0.07036077, 0.07079221, 0.07143381, 0.07164832, 
    0.07156644, 0.07142613, 0.07140836, 0.07102982, 0.07118194, 0.0712593, 
    0.07074569, 0.06993398, 0.0692274, 0.06894713, 0.06894831, 0.06947506, 
    0.07017947, 0.07037859, 0.07039479, 0.07060415, 0.07055131, 0.07079203, 
    0.07103982, 0.07103194, 0.07095318, 0.07074964, 0.07071764, 0.07055364, 
    0.07066095, 0.07050654, 0.07061018, 0.07043698, 0.06996621, 0.06930678, 
    0.06858902, 0.06778411, 0.06694862, 0.06620892, 0.06537756, 0.06433637, 
    0.06305403, 0.06176786, 0.06100503, 0.06052495, 0.06043628, 0.06068183, 
    0.06015207, 0.05918688, 0.05802651, 0.05696782, 0.05589574, 0.05485085, 
    0.05393973, 0.05309669, 0.05241073, 0.05187822, 0.05143174, 0.05064022, 
    0.0498524, 0.04913989, 0.04842126, 0.04779267, 0.04724422, 0.04666673,
  0.05168356, 0.05095723, 0.05029806, 0.04957866, 0.04853281, 0.04806982, 
    0.04788923, 0.04802903, 0.04845442, 0.04873728, 0.0491939, 0.04985449, 
    0.05013811, 0.05036051, 0.0504298, 0.05121019, 0.05231692, 0.05333052, 
    0.05404177, 0.05447168, 0.0546482, 0.05463275, 0.05486056, 0.05477288, 
    0.05428728, 0.05394482, 0.05379143, 0.05390889, 0.05425013, 0.05468408, 
    0.05491545, 0.05477099, 0.05454757, 0.05444471, 0.05440076, 0.05457398, 
    0.05481758, 0.05498273, 0.05528922, 0.05530559, 0.0556968, 0.0561285, 
    0.05658262, 0.05699849, 0.05732155, 0.05786747, 0.05857996, 0.05920678, 
    0.05914962, 0.05919351, 0.0591782, 0.05910439, 0.05882595, 0.05861199, 
    0.05850037, 0.05837318, 0.05833401, 0.05798998, 0.05751476, 0.05700103, 
    0.05623785, 0.05615769, 0.05628692, 0.05632096, 0.05621142, 0.05598987, 
    0.05571958, 0.05534943, 0.05456139, 0.05409384, 0.05360294, 0.05307476, 
    0.05242363, 0.0524695, 0.05259274, 0.05283938, 0.05307491, 0.05335833, 
    0.05335314, 0.0531524, 0.05322323, 0.05333075, 0.05371961, 0.05402047, 
    0.05408639, 0.05407574, 0.0540962, 0.05418532, 0.05448312, 0.05501673, 
    0.05557251, 0.05608542, 0.05652682, 0.05698325, 0.05727739, 0.0577106, 
    0.05844192, 0.05923473, 0.05980014, 0.06041333, 0.06109994, 0.06203387, 
    0.06337175, 0.06467288, 0.06591818, 0.06732293, 0.06864934, 0.06945849, 
    0.07004264, 0.07064736, 0.07157774, 0.07271103, 0.07355082, 0.07404967, 
    0.07425667, 0.07470905, 0.07545925, 0.07672756, 0.07830764, 0.07988118, 
    0.08099619, 0.081671, 0.08219074, 0.08241108, 0.08246598, 0.08266291, 
    0.08308683, 0.08349602, 0.08386675, 0.08430157, 0.08457128, 0.08452885, 
    0.08439062, 0.0842992, 0.08420485, 0.08403093, 0.08355251, 0.08242346, 
    0.08083565, 0.07941731, 0.07891483, 0.07869811, 0.07880348, 0.0789636, 
    0.0787252, 0.07855245, 0.07839158, 0.07826319, 0.07835985, 0.07889058, 
    0.07971054, 0.08063988, 0.08140268, 0.08205372, 0.08240289, 0.082803, 
    0.08337492, 0.0837161, 0.08398082, 0.08450877, 0.08505754, 0.08535006, 
    0.08572666, 0.08615965, 0.08681211, 0.08729137, 0.08753002, 0.08737648, 
    0.08710408, 0.08679095, 0.08629626, 0.08616443, 0.08644711, 0.08677168, 
    0.08690298, 0.08698793, 0.08695877, 0.08683863, 0.08677135, 0.08701906, 
    0.08739063, 0.08772097, 0.08799525, 0.08805276, 0.08756845, 0.08701814, 
    0.08643069, 0.08565848, 0.0844373, 0.08294068, 0.08165792, 0.08052832, 
    0.07985249, 0.07947508, 0.0786464, 0.07753342, 0.0769195, 0.07637715, 
    0.07585469, 0.07539436, 0.07418159, 0.07356001, 0.07316948, 0.07278444, 
    0.07243226, 0.07232823, 0.07230579, 0.07219331, 0.0719621, 0.071876, 
    0.07171579, 0.07165674, 0.07183295, 0.07210307, 0.07216989, 0.07211885, 
    0.07207082, 0.07168494, 0.07149765, 0.07137398, 0.07132009, 0.07138741, 
    0.07142084, 0.0715604, 0.07163464, 0.07172325, 0.07192878, 0.07201994, 
    0.07185299, 0.07169379, 0.07196003, 0.07311614, 0.07379474, 0.07300343, 
    0.07094441, 0.06846996, 0.06621666, 0.06544735, 0.0661663, 0.06718505, 
    0.06820346, 0.06913523, 0.06998863, 0.07076527, 0.07142506, 0.07210582, 
    0.07275324, 0.07324722, 0.07365826, 0.07372876, 0.07365572, 0.07347022, 
    0.07330337, 0.07334227, 0.07358748, 0.07382766, 0.07372715, 0.07338262, 
    0.07301339, 0.07247777, 0.07195199, 0.07119597, 0.07030179, 0.06922013, 
    0.06795763, 0.06680743, 0.06596017, 0.06534162, 0.06555606, 0.06554948, 
    0.06498033, 0.06395428, 0.06292161, 0.06215611, 0.06142632, 0.06037699, 
    0.0595461, 0.05871469, 0.05793237, 0.05721353, 0.05637984, 0.05573533, 
    0.05515965, 0.05460675, 0.05393816, 0.05311039, 0.05237135, 0.05186473,
  0.05732479, 0.0564675, 0.05569776, 0.05498951, 0.05429996, 0.05388044, 
    0.05352598, 0.05351675, 0.05370354, 0.05400915, 0.05487784, 0.05556471, 
    0.05589679, 0.05604652, 0.0563148, 0.05676164, 0.05746994, 0.05823391, 
    0.05868895, 0.05864324, 0.0586715, 0.05867741, 0.05865258, 0.05852604, 
    0.0581805, 0.05770332, 0.05731462, 0.0574667, 0.05790251, 0.05831205, 
    0.05840154, 0.05812863, 0.05780835, 0.05777495, 0.05793913, 0.05828276, 
    0.058743, 0.05936351, 0.05983356, 0.06031668, 0.06069664, 0.06107274, 
    0.06136533, 0.06151125, 0.06168363, 0.06206791, 0.06268696, 0.06330483, 
    0.06338304, 0.06322566, 0.0628344, 0.06264912, 0.06224774, 0.06182804, 
    0.06194305, 0.06174126, 0.06143175, 0.06110984, 0.06093358, 0.06076185, 
    0.06038479, 0.06038155, 0.06058235, 0.06072769, 0.06091523, 0.06084662, 
    0.06018399, 0.05914143, 0.05808134, 0.05719803, 0.05630696, 0.05577537, 
    0.0556959, 0.05605236, 0.05607332, 0.05640454, 0.05685027, 0.05723612, 
    0.05737502, 0.05738281, 0.05759712, 0.05799094, 0.05856158, 0.05872543, 
    0.05867111, 0.05881903, 0.05887241, 0.05881823, 0.05910909, 0.05960939, 
    0.06020072, 0.0607568, 0.06110741, 0.06127272, 0.06134418, 0.06171858, 
    0.06255537, 0.06348313, 0.0643198, 0.06503276, 0.06580611, 0.06688078, 
    0.06821892, 0.06953524, 0.0709404, 0.07229219, 0.07319565, 0.07386751, 
    0.0744903, 0.07505649, 0.07564531, 0.07622731, 0.07649851, 0.0766441, 
    0.07713373, 0.07786535, 0.07915977, 0.08111712, 0.08309017, 0.08453665, 
    0.08586666, 0.08693231, 0.08742191, 0.08734426, 0.08688575, 0.08639047, 
    0.08616822, 0.0862061, 0.08682078, 0.08760014, 0.08799949, 0.08758405, 
    0.08717059, 0.08661538, 0.08575635, 0.08461978, 0.08379867, 0.08273438, 
    0.08158699, 0.08077865, 0.08066012, 0.08070018, 0.08081032, 0.08085415, 
    0.08073223, 0.08067716, 0.07994916, 0.07947608, 0.07945518, 0.08001424, 
    0.08086813, 0.08171496, 0.08227999, 0.082753, 0.0834076, 0.08385185, 
    0.08431387, 0.08496504, 0.08572254, 0.08620641, 0.08657375, 0.0865154, 
    0.08638544, 0.08717875, 0.08792968, 0.08817738, 0.08807351, 0.08785841, 
    0.08807693, 0.08809533, 0.088169, 0.08861102, 0.08955511, 0.09013795, 
    0.09018856, 0.09023948, 0.09036244, 0.09049433, 0.09060326, 0.09077153, 
    0.09118994, 0.09146991, 0.0911348, 0.09067295, 0.09017483, 0.08944231, 
    0.08862963, 0.08745111, 0.08599836, 0.08481255, 0.08391414, 0.08333419, 
    0.08272286, 0.08186343, 0.08095317, 0.07978313, 0.07900525, 0.07846968, 
    0.07831256, 0.07722636, 0.07667537, 0.07634978, 0.07591098, 0.07561699, 
    0.07513591, 0.07494812, 0.07492874, 0.074786, 0.07437966, 0.07411475, 
    0.07390973, 0.07389805, 0.07428148, 0.07472847, 0.07456253, 0.07413399, 
    0.07373451, 0.0735811, 0.07338055, 0.07334534, 0.07339204, 0.07352301, 
    0.0732807, 0.07304379, 0.07275812, 0.07247297, 0.07281753, 0.07282107, 
    0.07283082, 0.07384189, 0.07707109, 0.07888362, 0.07663137, 0.07445381, 
    0.06958426, 0.06511424, 0.06257841, 0.06114026, 0.06145536, 0.06312685, 
    0.06510013, 0.06683175, 0.06864964, 0.07002418, 0.07112905, 0.0720919, 
    0.0732107, 0.07419542, 0.07481534, 0.07508763, 0.07540607, 0.07559458, 
    0.07579139, 0.07622673, 0.07646702, 0.07650013, 0.07697162, 0.07726675, 
    0.07690626, 0.07592712, 0.07513031, 0.07438136, 0.07323386, 0.07226414, 
    0.07148046, 0.0709808, 0.07057185, 0.06998225, 0.06974053, 0.06927747, 
    0.06867328, 0.06791673, 0.0671061, 0.06680437, 0.06672389, 0.06587181, 
    0.06497452, 0.06407885, 0.0632323, 0.06242102, 0.06179468, 0.06128073, 
    0.06076967, 0.06018225, 0.05953986, 0.05886944, 0.05831846, 0.05785649,
  0.06256698, 0.06171935, 0.061253, 0.0607293, 0.06041761, 0.05991105, 
    0.05921807, 0.05898522, 0.05893499, 0.05953984, 0.06036354, 0.0606995, 
    0.06115626, 0.06132721, 0.06140768, 0.0615277, 0.06202979, 0.06249066, 
    0.06245782, 0.06255668, 0.06269597, 0.06293473, 0.06314382, 0.06294645, 
    0.0623986, 0.06199137, 0.06189479, 0.06223579, 0.06260629, 0.06279074, 
    0.06260444, 0.06213503, 0.06180189, 0.06183839, 0.06256279, 0.06345406, 
    0.06429965, 0.06542195, 0.0662582, 0.0668147, 0.06687758, 0.06673229, 
    0.06671011, 0.06670702, 0.06656247, 0.06680825, 0.06708004, 0.06728809, 
    0.06746425, 0.06740604, 0.06690899, 0.06642933, 0.06589393, 0.06540801, 
    0.06522922, 0.06518637, 0.06498163, 0.06475325, 0.06478848, 0.06475733, 
    0.06479932, 0.06496416, 0.06514021, 0.06525785, 0.06564005, 0.06552965, 
    0.06479286, 0.06358419, 0.06229648, 0.06111048, 0.0601283, 0.05964454, 
    0.05968687, 0.05995141, 0.06017669, 0.06054996, 0.06077686, 0.0610457, 
    0.06134218, 0.06135359, 0.06189937, 0.06246527, 0.06306628, 0.06327301, 
    0.06370986, 0.06400102, 0.06418271, 0.0639314, 0.06398134, 0.06445903, 
    0.06489006, 0.06529082, 0.06581476, 0.06599713, 0.06628425, 0.06670326, 
    0.06736925, 0.06803212, 0.06889427, 0.06987546, 0.07092775, 0.07199954, 
    0.07294334, 0.07414852, 0.0754459, 0.07642752, 0.07714967, 0.07778874, 
    0.078477, 0.07879668, 0.07905435, 0.07954402, 0.07973012, 0.07995974, 
    0.081069, 0.08257904, 0.08421592, 0.08626886, 0.0878573, 0.08890712, 
    0.08995146, 0.09063525, 0.09116536, 0.09103604, 0.09024594, 0.08959755, 
    0.08874839, 0.08871255, 0.08928164, 0.09003446, 0.09039371, 0.09017525, 
    0.08928271, 0.08797464, 0.0863156, 0.0843898, 0.08308765, 0.08221766, 
    0.08163331, 0.08124296, 0.08110754, 0.0812232, 0.08145104, 0.08153205, 
    0.08136156, 0.08081914, 0.08010872, 0.07918885, 0.07901102, 0.0796297, 
    0.08054506, 0.08163118, 0.08220319, 0.08273839, 0.08327757, 0.08378104, 
    0.08412672, 0.08484256, 0.08593567, 0.08668573, 0.08691219, 0.08699055, 
    0.08688726, 0.08726376, 0.08787554, 0.08779702, 0.08808252, 0.088333, 
    0.08851428, 0.08875366, 0.08939648, 0.09038783, 0.09133994, 0.09202015, 
    0.09208048, 0.09196217, 0.09198228, 0.09209266, 0.09252833, 0.09296484, 
    0.09313561, 0.09289572, 0.09220868, 0.09183598, 0.09121551, 0.09058031, 
    0.08980551, 0.08877924, 0.08787551, 0.08697894, 0.08622141, 0.08564302, 
    0.08501093, 0.08415233, 0.08326153, 0.08246444, 0.08173903, 0.08108927, 
    0.07997171, 0.07881552, 0.07819062, 0.07808259, 0.07759637, 0.07739299, 
    0.0768456, 0.07636254, 0.07617708, 0.0761281, 0.07591651, 0.07593729, 
    0.0760817, 0.07620405, 0.07630589, 0.07640983, 0.0760618, 0.07556701, 
    0.07510181, 0.07495099, 0.07515854, 0.07555107, 0.07580722, 0.07579004, 
    0.07532887, 0.07460251, 0.07350798, 0.07347163, 0.07401678, 0.07473786, 
    0.07748538, 0.08251489, 0.08796172, 0.08378556, 0.08602515, 0.06504515, 
    0.05505193, 0.05300327, 0.0525586, 0.0534696, 0.0552515, 0.05767124, 
    0.0603369, 0.06284728, 0.06510016, 0.06706386, 0.06858042, 0.07006063, 
    0.07196048, 0.07358589, 0.07481843, 0.07551794, 0.07655165, 0.07720421, 
    0.07791177, 0.07863212, 0.07885166, 0.07928605, 0.08109448, 0.08210643, 
    0.08112339, 0.07950925, 0.07689162, 0.07578676, 0.07469923, 0.07390611, 
    0.07399055, 0.07427846, 0.07444084, 0.07441799, 0.07411408, 0.07333332, 
    0.0730126, 0.07234602, 0.07172296, 0.07143049, 0.07121551, 0.07062372, 
    0.06963024, 0.0687331, 0.0680094, 0.06721107, 0.06677759, 0.06648861, 
    0.06610418, 0.06558894, 0.06501736, 0.06449538, 0.0641875, 0.06349691,
  0.06806134, 0.06740931, 0.06705514, 0.06664153, 0.06582879, 0.06576285, 
    0.06561683, 0.06526808, 0.06501165, 0.06528362, 0.06567392, 0.06575344, 
    0.06583317, 0.06580048, 0.06567184, 0.06578294, 0.06629737, 0.06700783, 
    0.06727972, 0.06747789, 0.0676175, 0.06778198, 0.06799834, 0.06797657, 
    0.06761001, 0.06740601, 0.06750973, 0.06793903, 0.06801483, 0.06780653, 
    0.06751138, 0.06709523, 0.06704251, 0.06747796, 0.06824985, 0.06914188, 
    0.07039863, 0.07162985, 0.07272203, 0.07289065, 0.07269058, 0.07232094, 
    0.0718931, 0.07168407, 0.07145401, 0.07141257, 0.07149577, 0.07155646, 
    0.07138167, 0.07101388, 0.07061836, 0.0702697, 0.06991863, 0.06980985, 
    0.0698796, 0.06984349, 0.06964695, 0.0694336, 0.06889427, 0.06879278, 
    0.06912401, 0.06967606, 0.06987571, 0.06992538, 0.07015511, 0.06998895, 
    0.06911223, 0.06782978, 0.06664832, 0.06582653, 0.06527828, 0.06489662, 
    0.0647845, 0.06487384, 0.06495707, 0.06510586, 0.06550911, 0.06582361, 
    0.06590076, 0.06593717, 0.0661976, 0.06676598, 0.06742856, 0.06816713, 
    0.0687812, 0.06907488, 0.06909344, 0.0688476, 0.06861315, 0.06888337, 
    0.06941988, 0.06968229, 0.07022041, 0.07074702, 0.07148981, 0.07229571, 
    0.07288975, 0.07352956, 0.07431571, 0.07506927, 0.07583243, 0.0766645, 
    0.07765286, 0.07853811, 0.07969337, 0.08038899, 0.08079008, 0.08122237, 
    0.0817768, 0.08209747, 0.08244532, 0.08307625, 0.08372396, 0.08447056, 
    0.08566868, 0.08731471, 0.08886446, 0.09035873, 0.09148843, 0.09219324, 
    0.09305675, 0.09348878, 0.09319473, 0.09233054, 0.09155183, 0.09109038, 
    0.09075706, 0.09052895, 0.09058864, 0.09125611, 0.09178153, 0.09125734, 
    0.08971639, 0.0878066, 0.0858531, 0.08388223, 0.0825287, 0.08201642, 
    0.08155931, 0.08100096, 0.08066264, 0.0809243, 0.08170802, 0.08176305, 
    0.0812574, 0.08033015, 0.07918061, 0.07827457, 0.07795445, 0.07891393, 
    0.07993556, 0.08091882, 0.08184322, 0.08258206, 0.08312693, 0.0836629, 
    0.08413009, 0.08449972, 0.08514835, 0.08569495, 0.08603552, 0.08643541, 
    0.08672217, 0.08682501, 0.08695109, 0.08726407, 0.08783388, 0.08831132, 
    0.0886613, 0.08930682, 0.09023092, 0.09130507, 0.09196554, 0.09196093, 
    0.09215076, 0.09225952, 0.09229033, 0.09266848, 0.0932799, 0.09356654, 
    0.09345627, 0.09319876, 0.09290278, 0.09244081, 0.09179983, 0.09102453, 
    0.09046876, 0.09010201, 0.08948001, 0.08880928, 0.08815995, 0.08742609, 
    0.08683135, 0.08572839, 0.08436718, 0.08359836, 0.08292649, 0.08220651, 
    0.08128446, 0.08034316, 0.0797166, 0.07961614, 0.07930772, 0.07867365, 
    0.07788885, 0.07724971, 0.07699104, 0.07716993, 0.07731662, 0.07732151, 
    0.07746303, 0.07725689, 0.07689362, 0.07670841, 0.07654, 0.07634008, 
    0.07625858, 0.0763776, 0.0767061, 0.07704721, 0.07722884, 0.07702154, 
    0.07639589, 0.07545763, 0.07494725, 0.07529034, 0.07605702, 0.08022449, 
    0.08592824, 0.09363875, 0.1019042, 0.09950979, 0.1044423, 0.07421599, 
    0.04689812, 0.04113439, 0.04320152, 0.04590088, 0.04953572, 0.05307405, 
    0.05616447, 0.05887133, 0.0610564, 0.06287903, 0.06476977, 0.06690748, 
    0.06922752, 0.07155862, 0.07358623, 0.07532881, 0.07702346, 0.07837212, 
    0.07915644, 0.07969977, 0.08015843, 0.08152297, 0.08446294, 0.08649807, 
    0.09129975, 0.0787135, 0.07138932, 0.07481938, 0.07590976, 0.07665044, 
    0.07758323, 0.07832618, 0.07873099, 0.07890669, 0.078522, 0.07773478, 
    0.07712864, 0.07672771, 0.07639007, 0.07607478, 0.07558529, 0.07495158, 
    0.07411992, 0.07321382, 0.07239285, 0.07183213, 0.0714839, 0.0708723, 
    0.0705783, 0.07009558, 0.06972662, 0.06972323, 0.06958476, 0.0689189,
  0.07337572, 0.07283019, 0.07232457, 0.07169212, 0.07110767, 0.07099082, 
    0.07113343, 0.07078948, 0.07034048, 0.07035414, 0.07064754, 0.07072832, 
    0.0706535, 0.07055888, 0.07050177, 0.07072945, 0.0711967, 0.07188333, 
    0.07239498, 0.07287421, 0.07314754, 0.07324475, 0.0734882, 0.07337161, 
    0.07329581, 0.07381033, 0.07388162, 0.07360305, 0.0734401, 0.07317028, 
    0.07278913, 0.07259177, 0.07275829, 0.07317067, 0.07371955, 0.07459721, 
    0.07544976, 0.07626171, 0.07698738, 0.07732667, 0.077191, 0.07687231, 
    0.07657649, 0.07638243, 0.07618608, 0.07596626, 0.07581647, 0.07572379, 
    0.07544321, 0.07498036, 0.07460632, 0.07425337, 0.07401963, 0.07399662, 
    0.07416471, 0.07420664, 0.07422273, 0.07430726, 0.07488269, 0.07317839, 
    0.07182629, 0.0733, 0.07390771, 0.07417233, 0.07435854, 0.07392618, 
    0.07308682, 0.07217287, 0.07142436, 0.07104339, 0.07085268, 0.07051222, 
    0.07016663, 0.06990945, 0.06960276, 0.06970296, 0.07028548, 0.07092187, 
    0.07118867, 0.07118145, 0.07142123, 0.07159768, 0.07187421, 0.07223666, 
    0.07250652, 0.07276461, 0.07276661, 0.07251565, 0.07270616, 0.07311692, 
    0.07393426, 0.07476689, 0.07528424, 0.07568152, 0.07634897, 0.07699663, 
    0.07751552, 0.07787579, 0.07838649, 0.07891341, 0.07975578, 0.08091308, 
    0.08197637, 0.08291267, 0.08390099, 0.08433002, 0.08480892, 0.08522782, 
    0.08541131, 0.08556934, 0.0859174, 0.0866247, 0.08741527, 0.08834068, 
    0.08924648, 0.09022579, 0.09182201, 0.09296963, 0.09363904, 0.09393954, 
    0.0939279, 0.09378619, 0.09314933, 0.09240656, 0.09193244, 0.09171375, 
    0.09133981, 0.09098416, 0.09101299, 0.09114538, 0.09112324, 0.09001194, 
    0.08818067, 0.0864659, 0.08480431, 0.08385074, 0.08296225, 0.08221979, 
    0.08114321, 0.07996953, 0.07958801, 0.07988668, 0.08018683, 0.08014327, 
    0.0797631, 0.07906517, 0.07836809, 0.07801796, 0.07794608, 0.07844695, 
    0.07922879, 0.0799107, 0.08105768, 0.08195537, 0.08253591, 0.08315843, 
    0.08427762, 0.08402446, 0.08406643, 0.08449899, 0.08521932, 0.08565859, 
    0.08577579, 0.08591423, 0.08630079, 0.08667697, 0.08674049, 0.08704229, 
    0.08733392, 0.08876913, 0.09010131, 0.09126376, 0.09161533, 0.09129664, 
    0.09122329, 0.09101073, 0.09105546, 0.09145906, 0.09210225, 0.09245103, 
    0.09278666, 0.09240049, 0.09196616, 0.09139363, 0.09087373, 0.09045669, 
    0.09028686, 0.08981647, 0.08930201, 0.08911468, 0.08879901, 0.0883059, 
    0.0875541, 0.08643416, 0.08527692, 0.08460747, 0.08389877, 0.08284971, 
    0.08172645, 0.08089836, 0.0802486, 0.08002068, 0.07951036, 0.07883902, 
    0.07846586, 0.07841606, 0.07852836, 0.07880757, 0.07885379, 0.07874059, 
    0.07843313, 0.07777379, 0.07726865, 0.07704227, 0.07689136, 0.07686687, 
    0.07703566, 0.07724949, 0.07769797, 0.07802013, 0.07794928, 0.07747667, 
    0.07702038, 0.0762972, 0.07629004, 0.07659528, 0.08022255, 0.08832441, 
    0.09684066, 0.1094571, 0.09946714, 0.07516374, 0.06194755, 0.04495496, 
    0.03452629, 0.0363835, 0.03835746, 0.04188551, 0.04663786, 0.05129994, 
    0.05470608, 0.05657831, 0.05787846, 0.05970144, 0.06190778, 0.06431046, 
    0.06668399, 0.06914704, 0.07201184, 0.07459979, 0.07684799, 0.07865213, 
    0.0798685, 0.08049888, 0.08137257, 0.08306353, 0.08510944, 0.08735839, 
    0.08930041, 0.07904446, 0.07518626, 0.07819644, 0.07998858, 0.08139712, 
    0.08275791, 0.08376948, 0.08397204, 0.08395049, 0.08352853, 0.08272943, 
    0.0821086, 0.08184277, 0.08159645, 0.0814226, 0.08078713, 0.07993644, 
    0.07901045, 0.077991, 0.07717556, 0.07654062, 0.07611383, 0.07575481, 
    0.07538966, 0.07490289, 0.07467635, 0.07477357, 0.07464437, 0.07410867,
  0.07789245, 0.07732895, 0.07686903, 0.07652632, 0.07623029, 0.07592928, 
    0.07585824, 0.07545927, 0.07469437, 0.0742876, 0.07476608, 0.07541133, 
    0.07585364, 0.07586996, 0.07586712, 0.07632104, 0.07675857, 0.07704373, 
    0.0772625, 0.07753681, 0.07787567, 0.07816294, 0.07875451, 0.07912112, 
    0.0793743, 0.07970412, 0.07956451, 0.07915526, 0.07882924, 0.07846312, 
    0.07804953, 0.07805208, 0.07806899, 0.07832414, 0.07871748, 0.07936385, 
    0.07999695, 0.08056888, 0.0811561, 0.08141378, 0.08118799, 0.08059953, 
    0.08032553, 0.08007689, 0.07998664, 0.08009383, 0.08007728, 0.0799135, 
    0.07965873, 0.07951508, 0.0794113, 0.07908072, 0.07866536, 0.0782735, 
    0.07842858, 0.0783594, 0.07841121, 0.07856178, 0.07801881, 0.07675281, 
    0.07639888, 0.07734012, 0.07839107, 0.07941551, 0.07965139, 0.07900756, 
    0.07792888, 0.07700249, 0.07671987, 0.07652374, 0.07601357, 0.07552087, 
    0.07531676, 0.07512216, 0.07457595, 0.07435455, 0.07457123, 0.07517117, 
    0.07567219, 0.07594217, 0.07622416, 0.07619605, 0.07624951, 0.07615262, 
    0.07606707, 0.07602559, 0.07604899, 0.07634833, 0.07700412, 0.07786725, 
    0.07877883, 0.07936051, 0.07983369, 0.08027014, 0.08071213, 0.08107193, 
    0.08162611, 0.08235281, 0.08317192, 0.08401726, 0.0848882, 0.08588769, 
    0.08676789, 0.08746694, 0.08825386, 0.08882863, 0.08882124, 0.08869908, 
    0.08871593, 0.08869965, 0.08920228, 0.089895, 0.09054573, 0.09101911, 
    0.09174495, 0.09299257, 0.09406397, 0.09455057, 0.09449789, 0.09389322, 
    0.0932373, 0.09271928, 0.09237967, 0.09221556, 0.09187242, 0.09171216, 
    0.09110349, 0.09062253, 0.09047281, 0.09010853, 0.0894953, 0.08840226, 
    0.08668796, 0.0852988, 0.08456109, 0.08429953, 0.08326753, 0.08178665, 
    0.08024342, 0.07895651, 0.07831518, 0.07801188, 0.07791584, 0.07789974, 
    0.07774116, 0.07748588, 0.07740244, 0.07785054, 0.07808018, 0.07823153, 
    0.07836513, 0.07881551, 0.07985163, 0.08086005, 0.08149998, 0.08225995, 
    0.08264431, 0.08260883, 0.08260661, 0.08287623, 0.08335177, 0.08370106, 
    0.08378258, 0.08432986, 0.08495793, 0.08527696, 0.08539689, 0.0857688, 
    0.08655777, 0.08790441, 0.08911826, 0.08970215, 0.08972915, 0.08947691, 
    0.08904425, 0.08851852, 0.08859511, 0.08889199, 0.08962338, 0.0905193, 
    0.09108662, 0.09108599, 0.09073385, 0.09025905, 0.08961163, 0.08940243, 
    0.08914375, 0.08868088, 0.08821744, 0.08792516, 0.0880101, 0.08794978, 
    0.08712026, 0.08600456, 0.08526009, 0.08509982, 0.08454841, 0.08350812, 
    0.0821532, 0.08115946, 0.08028206, 0.07981696, 0.07978888, 0.0797277, 
    0.07952093, 0.07967541, 0.08016721, 0.08055689, 0.08059601, 0.08036412, 
    0.0802437, 0.07984814, 0.07953654, 0.07904474, 0.07871332, 0.07871277, 
    0.07863104, 0.07845516, 0.07860153, 0.07855622, 0.07831165, 0.07806005, 
    0.07749475, 0.07707615, 0.077489, 0.07949936, 0.0864793, 0.09768684, 
    0.1121858, 0.1121673, 0.07887954, 0.05868736, 0.04526193, 0.03507347, 
    0.0326783, 0.03415642, 0.03696572, 0.04155983, 0.04696572, 0.0517223, 
    0.05248553, 0.05284446, 0.05352128, 0.05580293, 0.058958, 0.06193439, 
    0.06483237, 0.06802142, 0.07144821, 0.0747446, 0.07735375, 0.07925189, 
    0.08100129, 0.08246371, 0.08380911, 0.08503735, 0.08615035, 0.08714493, 
    0.0871741, 0.08551953, 0.08444006, 0.08463348, 0.08592907, 0.08765235, 
    0.08861599, 0.08925955, 0.08910784, 0.08860446, 0.08829936, 0.08767304, 
    0.08687496, 0.08634038, 0.0860569, 0.08593006, 0.08549458, 0.08474601, 
    0.0837848, 0.08267386, 0.08208505, 0.08140977, 0.08083028, 0.08053894, 
    0.08022323, 0.07990091, 0.07943536, 0.0793508, 0.0791246, 0.07850116,
  0.08237836, 0.08166405, 0.08101422, 0.08059917, 0.08038256, 0.08031027, 
    0.08008474, 0.07950689, 0.07901601, 0.07898573, 0.07941543, 0.07992294, 
    0.08056317, 0.08138371, 0.08186392, 0.08203905, 0.08205466, 0.08180404, 
    0.08238147, 0.08287677, 0.08343059, 0.08387041, 0.08425239, 0.0846225, 
    0.08465684, 0.0844866, 0.08418418, 0.08397845, 0.08360139, 0.08308744, 
    0.08275896, 0.08252551, 0.08257703, 0.08289043, 0.0834192, 0.08376554, 
    0.08446287, 0.08525193, 0.08550932, 0.08516643, 0.08454049, 0.0839924, 
    0.08373251, 0.08377306, 0.08399115, 0.08422547, 0.08437829, 0.08422828, 
    0.08363733, 0.08334547, 0.08318198, 0.08307061, 0.08280596, 0.08327606, 
    0.08396889, 0.08359285, 0.08282278, 0.08248869, 0.08154651, 0.08094104, 
    0.08096482, 0.08169097, 0.08313065, 0.08450146, 0.08458692, 0.08404312, 
    0.08303789, 0.08215879, 0.08186476, 0.08183523, 0.08157077, 0.08150634, 
    0.08135869, 0.08084545, 0.07996863, 0.07928787, 0.07916924, 0.07928804, 
    0.07944921, 0.07971487, 0.07994499, 0.08011428, 0.0798387, 0.07956952, 
    0.07955173, 0.08002186, 0.08037786, 0.08077965, 0.08156813, 0.08246481, 
    0.08278801, 0.08311599, 0.08338346, 0.08367033, 0.08417239, 0.0851215, 
    0.08624268, 0.08735946, 0.08808334, 0.08862008, 0.08915728, 0.08992755, 
    0.09065818, 0.09123292, 0.09148982, 0.09132193, 0.09121072, 0.09169743, 
    0.09180073, 0.09181572, 0.09180415, 0.09166762, 0.09149554, 0.09150778, 
    0.0920799, 0.09323913, 0.09375553, 0.09332987, 0.0923402, 0.09129446, 
    0.09079707, 0.09060019, 0.09042372, 0.08989398, 0.08945626, 0.08901022, 
    0.0887433, 0.08867352, 0.08865863, 0.08864326, 0.08835009, 0.08739282, 
    0.08573765, 0.08325138, 0.08317333, 0.08316156, 0.0822735, 0.08108376, 
    0.08005924, 0.07888716, 0.07731164, 0.07630005, 0.07599144, 0.07569794, 
    0.07535314, 0.07553163, 0.07654639, 0.07769413, 0.07817631, 0.07833929, 
    0.07781468, 0.07772458, 0.07831115, 0.07918617, 0.07998908, 0.0805205, 
    0.08070833, 0.08136361, 0.08194952, 0.08212893, 0.08222739, 0.082601, 
    0.08261961, 0.08335988, 0.0840513, 0.08437428, 0.08447545, 0.08485638, 
    0.0859124, 0.0868454, 0.08722138, 0.08722069, 0.08712935, 0.08726998, 
    0.08732723, 0.08732987, 0.08740386, 0.08786561, 0.0886111, 0.08928584, 
    0.08982162, 0.08999125, 0.08975096, 0.0898146, 0.08917509, 0.08851171, 
    0.08842605, 0.08799406, 0.08760475, 0.08719535, 0.08711869, 0.0872084, 
    0.08708948, 0.0866171, 0.08611717, 0.0855248, 0.08474807, 0.08381609, 
    0.08284973, 0.08213962, 0.08148207, 0.08121964, 0.08150946, 0.08175866, 
    0.08152039, 0.08157881, 0.08176822, 0.08218428, 0.08204649, 0.08227928, 
    0.08222597, 0.08195116, 0.08154426, 0.08087457, 0.08053102, 0.08051176, 
    0.08032705, 0.07983468, 0.07976769, 0.0800001, 0.07970288, 0.07927412, 
    0.07866924, 0.07877296, 0.07991998, 0.0835269, 0.09436967, 0.1082954, 
    0.1216911, 0.1144317, 0.0661028, 0.04579524, 0.03833617, 0.03353801, 
    0.03197777, 0.0328017, 0.03677171, 0.04182606, 0.04607497, 0.04974676, 
    0.04979283, 0.0468232, 0.04762188, 0.05201374, 0.0560099, 0.05980418, 
    0.06323992, 0.06666386, 0.07020491, 0.07351279, 0.07683269, 0.07954957, 
    0.08175254, 0.08357085, 0.08524344, 0.08660218, 0.08784099, 0.08875765, 
    0.0891517, 0.08955332, 0.08994929, 0.0904491, 0.09116187, 0.09164412, 
    0.09228486, 0.0928598, 0.09265498, 0.09202062, 0.09136017, 0.09079387, 
    0.09020106, 0.08955279, 0.08905008, 0.08890638, 0.08872293, 0.08801588, 
    0.08717289, 0.0865124, 0.08608135, 0.0855296, 0.08493327, 0.08425699, 
    0.08394345, 0.08390253, 0.08381157, 0.08383109, 0.08341973, 0.0829315,
  0.08651438, 0.08615573, 0.08551817, 0.0848859, 0.0847014, 0.08474758, 
    0.08466142, 0.08432296, 0.08412202, 0.08398408, 0.08420206, 0.08478817, 
    0.08599009, 0.08708552, 0.08755268, 0.08747056, 0.08707496, 0.08709219, 
    0.08780308, 0.08828142, 0.08847144, 0.08869421, 0.08872809, 0.0887157, 
    0.08861738, 0.08843447, 0.08819719, 0.08816931, 0.08784224, 0.08712886, 
    0.08691046, 0.08704636, 0.08692774, 0.08728367, 0.08796676, 0.08822878, 
    0.0883257, 0.08848018, 0.08846049, 0.08832305, 0.08785429, 0.08747424, 
    0.08744083, 0.08743245, 0.08775008, 0.08788832, 0.08803885, 0.08799688, 
    0.08776385, 0.08764007, 0.08758137, 0.08753272, 0.08785044, 0.08975343, 
    0.09125609, 0.08912952, 0.08489758, 0.08683483, 0.08623222, 0.08533001, 
    0.08563346, 0.08657019, 0.08791094, 0.08880384, 0.08909228, 0.08882708, 
    0.08824991, 0.08771799, 0.08718205, 0.08678633, 0.08663564, 0.08662771, 
    0.08591676, 0.08507627, 0.0842424, 0.08363544, 0.08347557, 0.08314869, 
    0.08290432, 0.08279274, 0.08257873, 0.08255327, 0.08240711, 0.08262752, 
    0.08338301, 0.08406446, 0.08433668, 0.08472587, 0.08586565, 0.08644207, 
    0.08634291, 0.08640271, 0.0867534, 0.08723843, 0.0879218, 0.08907537, 
    0.09059999, 0.09179859, 0.09226141, 0.0925373, 0.09259424, 0.09255663, 
    0.09283794, 0.09310365, 0.09326392, 0.09309936, 0.09325852, 0.09346122, 
    0.09351535, 0.09322163, 0.09248461, 0.09192038, 0.09141851, 0.0912461, 
    0.09135275, 0.09119418, 0.09094165, 0.08981181, 0.08855351, 0.0878097, 
    0.08761611, 0.0873346, 0.08682435, 0.08644545, 0.08622828, 0.08606946, 
    0.08601721, 0.08664192, 0.0872832, 0.0873106, 0.08681305, 0.08584233, 
    0.08446331, 0.08154812, 0.08122627, 0.08153011, 0.08077153, 0.07960535, 
    0.0785792, 0.07753149, 0.0760266, 0.07479198, 0.07406046, 0.0735135, 
    0.07373122, 0.07441954, 0.07598968, 0.07734761, 0.07826222, 0.07818815, 
    0.07749303, 0.07699486, 0.07711571, 0.0777325, 0.07847199, 0.0787223, 
    0.07948102, 0.08023686, 0.080876, 0.08141091, 0.08192233, 0.08246024, 
    0.08280375, 0.08289757, 0.08283441, 0.08289447, 0.0829244, 0.08336956, 
    0.08437078, 0.08508046, 0.08530325, 0.08540776, 0.08559761, 0.08610903, 
    0.08634825, 0.08678745, 0.08733262, 0.08793636, 0.08848931, 0.08896621, 
    0.08954695, 0.08969549, 0.08938741, 0.08921908, 0.08909058, 0.08850656, 
    0.08823262, 0.08860551, 0.08855426, 0.08783704, 0.08763808, 0.08753639, 
    0.08757622, 0.08756985, 0.08713961, 0.08627649, 0.08534054, 0.08465767, 
    0.08412824, 0.08421498, 0.08413723, 0.08356449, 0.08354549, 0.08343948, 
    0.08345036, 0.08362322, 0.0833277, 0.08343023, 0.08359063, 0.08386716, 
    0.08362292, 0.08322414, 0.08252542, 0.08182439, 0.08176289, 0.08175104, 
    0.08157325, 0.08136256, 0.08159181, 0.08181423, 0.08136245, 0.08032846, 
    0.07938161, 0.07935778, 0.08087881, 0.08728927, 0.10323, 0.1179559, 
    0.1489135, 0.1237568, 0.05953136, 0.03541905, 0.03613668, 0.03161893, 
    0.03026233, 0.03110863, 0.03470659, 0.03947055, 0.04224958, 0.04291156, 
    0.04289018, 0.04319024, 0.04609917, 0.05005176, 0.05400314, 0.05799688, 
    0.06162178, 0.06495519, 0.06787009, 0.07115107, 0.07482085, 0.07813961, 
    0.08069851, 0.08267333, 0.08440614, 0.08610315, 0.08832569, 0.09024616, 
    0.0917234, 0.09283505, 0.09376859, 0.09394685, 0.09335171, 0.09320239, 
    0.09335381, 0.09348825, 0.0936042, 0.0935962, 0.09333474, 0.09290937, 
    0.09242625, 0.09185044, 0.09079182, 0.09045919, 0.09047891, 0.09005911, 
    0.08926842, 0.0886024, 0.0883493, 0.08785024, 0.08746511, 0.08730144, 
    0.0873438, 0.0873955, 0.08748318, 0.08739983, 0.08711667, 0.08670703,
  0.08978042, 0.08970959, 0.08956942, 0.08956465, 0.08976822, 0.08965601, 
    0.08935209, 0.08903031, 0.08892362, 0.08894137, 0.08919089, 0.08996013, 
    0.09097699, 0.09171399, 0.09174911, 0.09162979, 0.09157933, 0.09179706, 
    0.09230111, 0.09246063, 0.09251787, 0.09234859, 0.09206304, 0.09182683, 
    0.09191052, 0.09183732, 0.09168259, 0.09136517, 0.09093513, 0.09040648, 
    0.09020063, 0.09062961, 0.09112937, 0.09152758, 0.09168541, 0.09142861, 
    0.09106745, 0.09081682, 0.09056016, 0.09033883, 0.09025232, 0.09045392, 
    0.09044997, 0.09025891, 0.09032156, 0.09037922, 0.0905313, 0.09069614, 
    0.09074598, 0.09113268, 0.09151736, 0.09184116, 0.09239297, 0.0948035, 
    0.09970434, 0.1019035, 0.08454322, 0.08579364, 0.08849458, 0.08911245, 
    0.08987064, 0.09104627, 0.09205203, 0.092583, 0.09306057, 0.09315464, 
    0.09297573, 0.09262571, 0.09239547, 0.09173841, 0.09115112, 0.09068158, 
    0.08994744, 0.08912782, 0.08805894, 0.08735421, 0.08672407, 0.08604588, 
    0.08562486, 0.08549607, 0.08560871, 0.08592609, 0.08621387, 0.08672719, 
    0.0871321, 0.08760331, 0.08804365, 0.08865989, 0.08912092, 0.08912434, 
    0.08922961, 0.08973885, 0.09046826, 0.09092385, 0.09151389, 0.09239765, 
    0.09381109, 0.09475125, 0.09504318, 0.09472679, 0.09447706, 0.09419568, 
    0.09425298, 0.09429454, 0.09411081, 0.09387833, 0.09377386, 0.09364455, 
    0.09344935, 0.09302501, 0.09220693, 0.09141782, 0.09051649, 0.08954571, 
    0.0885931, 0.08753571, 0.08667263, 0.08562349, 0.08491885, 0.08477619, 
    0.08470687, 0.08447669, 0.08380744, 0.08338166, 0.08344231, 0.08414945, 
    0.08453671, 0.08517043, 0.08570254, 0.08492193, 0.08339816, 0.08237337, 
    0.08142226, 0.08081114, 0.08013757, 0.07916419, 0.07722056, 0.0758537, 
    0.07482377, 0.07425831, 0.07398937, 0.07392564, 0.07338408, 0.07259564, 
    0.07258566, 0.07279064, 0.07392608, 0.07564951, 0.07692189, 0.0770476, 
    0.07648742, 0.07545953, 0.07589785, 0.07669248, 0.07749154, 0.07802192, 
    0.078502, 0.07908884, 0.07966472, 0.08064318, 0.08146139, 0.08160932, 
    0.08167936, 0.08159273, 0.08184575, 0.08159608, 0.08146637, 0.08196392, 
    0.08301498, 0.08355278, 0.08369369, 0.08410104, 0.08470563, 0.08511787, 
    0.08502679, 0.08551773, 0.0860014, 0.08694158, 0.08747501, 0.08780077, 
    0.08798026, 0.08804366, 0.08854233, 0.08914319, 0.08904579, 0.08909751, 
    0.08921452, 0.08946281, 0.08951664, 0.08915903, 0.08861395, 0.08810633, 
    0.0876283, 0.0872642, 0.08675753, 0.08671907, 0.08677902, 0.08686138, 
    0.08667805, 0.08669353, 0.08673832, 0.0861065, 0.08538531, 0.08496646, 
    0.08487647, 0.08482428, 0.08465341, 0.08479101, 0.08504008, 0.08525673, 
    0.08500752, 0.0845107, 0.0837841, 0.08348586, 0.08406261, 0.08436076, 
    0.08386768, 0.08409918, 0.08441886, 0.08404575, 0.08309239, 0.08125268, 
    0.07940818, 0.07903851, 0.08083935, 0.08976487, 0.1080244, 0.1342885, 
    0.1668117, 0.1272506, 0.05683933, 0.03242402, 0.03417606, 0.03091573, 
    0.0284386, 0.02986961, 0.03301746, 0.03666428, 0.03937807, 0.0407583, 
    0.04152657, 0.04308715, 0.04578581, 0.04919145, 0.05296407, 0.0569345, 
    0.05987194, 0.06254881, 0.06561752, 0.06904542, 0.07280244, 0.07605915, 
    0.07826427, 0.08010244, 0.08229244, 0.08480225, 0.0875609, 0.0898255, 
    0.09176359, 0.09283457, 0.09336456, 0.09328987, 0.09349602, 0.0937521, 
    0.09394151, 0.09425072, 0.09464611, 0.09501065, 0.09481774, 0.09456095, 
    0.09378082, 0.09319232, 0.09247623, 0.09199946, 0.09179983, 0.09165099, 
    0.09129237, 0.09080993, 0.09024004, 0.08942853, 0.0894875, 0.08978668, 
    0.09017385, 0.09011526, 0.09002693, 0.08998621, 0.0900576, 0.08974352,
  0.09394465, 0.09415449, 0.09425548, 0.09402498, 0.0938654, 0.09359621, 
    0.09336862, 0.09333852, 0.0935747, 0.09377171, 0.09394965, 0.09434994, 
    0.09493764, 0.09492588, 0.09470655, 0.09455246, 0.09460099, 0.09465277, 
    0.09466013, 0.09480828, 0.09505805, 0.09490859, 0.09464736, 0.0947677, 
    0.0946514, 0.0940666, 0.09353562, 0.09296552, 0.09240498, 0.09214155, 
    0.09270577, 0.09354252, 0.09419981, 0.09425371, 0.09414105, 0.09402873, 
    0.09368403, 0.09310432, 0.09273292, 0.0927977, 0.09303751, 0.0933229, 
    0.0931391, 0.09302097, 0.0931573, 0.09325114, 0.09339151, 0.09332064, 
    0.09300707, 0.09295526, 0.09329545, 0.09367626, 0.09405366, 0.09542084, 
    0.09911446, 0.09595216, 0.08773614, 0.08850186, 0.09161483, 0.09325694, 
    0.09443737, 0.09546566, 0.0959807, 0.09637181, 0.09695439, 0.09711993, 
    0.09722062, 0.09713959, 0.09668594, 0.09581685, 0.09488797, 0.09429301, 
    0.09362593, 0.09278512, 0.0918151, 0.09090321, 0.08985317, 0.08908124, 
    0.08892542, 0.08912406, 0.08953308, 0.09002164, 0.09017055, 0.09047269, 
    0.09062566, 0.09085751, 0.09168457, 0.09206786, 0.09184802, 0.09175646, 
    0.09255408, 0.0932492, 0.09361685, 0.09411688, 0.09482666, 0.09579161, 
    0.09647597, 0.09635928, 0.09551642, 0.09499077, 0.09461819, 0.09434875, 
    0.09418178, 0.09400278, 0.09361756, 0.09290447, 0.0921382, 0.09179763, 
    0.09130984, 0.09066517, 0.08954091, 0.08798473, 0.08626635, 0.08499949, 
    0.08391778, 0.08280587, 0.08157824, 0.0807436, 0.08041133, 0.08040775, 
    0.0804966, 0.08049211, 0.07981886, 0.07923746, 0.07960531, 0.08064, 
    0.08165782, 0.08213234, 0.08177785, 0.08067387, 0.07971647, 0.07904299, 
    0.07987174, 0.08133099, 0.07992844, 0.07542653, 0.07093282, 0.06837218, 
    0.06766902, 0.06871224, 0.0702633, 0.07145684, 0.07157438, 0.07105389, 
    0.07063252, 0.07047024, 0.07110138, 0.07260317, 0.0741438, 0.07490046, 
    0.0750117, 0.07488348, 0.07556249, 0.07645097, 0.07705043, 0.07720593, 
    0.07710412, 0.07786477, 0.07926188, 0.08045945, 0.08078649, 0.08039434, 
    0.08017158, 0.08055878, 0.08075023, 0.08041014, 0.08036629, 0.08142336, 
    0.08258374, 0.0834421, 0.08369999, 0.0838981, 0.08405121, 0.08401883, 
    0.08409278, 0.08478418, 0.08517347, 0.08577432, 0.08578579, 0.08595516, 
    0.08634264, 0.08680368, 0.08752975, 0.08817457, 0.08849549, 0.08872008, 
    0.08886469, 0.08870663, 0.08876608, 0.08890066, 0.08881757, 0.08817777, 
    0.08762132, 0.08713833, 0.08683412, 0.08696972, 0.08755331, 0.08815789, 
    0.08797082, 0.08769568, 0.0878441, 0.08778644, 0.0871224, 0.08626296, 
    0.08565418, 0.08563188, 0.08554459, 0.08586296, 0.08606308, 0.08686855, 
    0.0870225, 0.08606386, 0.08544738, 0.08597939, 0.08690374, 0.0869264, 
    0.08623277, 0.08619417, 0.08627128, 0.08582995, 0.08440871, 0.08174785, 
    0.07959991, 0.07903264, 0.08039398, 0.08827855, 0.1084586, 0.1383864, 
    0.1816737, 0.1518816, 0.07795779, 0.0320515, 0.02993213, 0.02935719, 
    0.02747638, 0.02842366, 0.03022252, 0.03362906, 0.03682893, 0.03854083, 
    0.03956473, 0.04136844, 0.04462387, 0.04879975, 0.05246795, 0.05594195, 
    0.05925098, 0.06210763, 0.06513906, 0.06837921, 0.07138971, 0.07359643, 
    0.07562845, 0.07776955, 0.0809159, 0.08430675, 0.08675003, 0.08882698, 
    0.09048963, 0.09136705, 0.09226894, 0.09304228, 0.09381858, 0.09439672, 
    0.09471379, 0.09493434, 0.09521964, 0.09550751, 0.09547639, 0.09520816, 
    0.09471788, 0.09445875, 0.09421626, 0.09370369, 0.09359149, 0.0936598, 
    0.09389564, 0.09369735, 0.0928141, 0.09188332, 0.09183286, 0.09228213, 
    0.09271741, 0.09305036, 0.09372086, 0.09415276, 0.09405933, 0.09387358,
  0.09857439, 0.09842835, 0.09812576, 0.09742013, 0.09720101, 0.09713096, 
    0.09738433, 0.09745998, 0.09773131, 0.09774744, 0.09788687, 0.09828811, 
    0.09829192, 0.0978576, 0.09713884, 0.09618182, 0.09556183, 0.09552336, 
    0.09586006, 0.09575731, 0.09570223, 0.09589835, 0.09588721, 0.09595615, 
    0.09555621, 0.09470534, 0.09383331, 0.0933034, 0.09326348, 0.09367196, 
    0.09477805, 0.09487641, 0.09617464, 0.09616395, 0.09590517, 0.09607298, 
    0.09584005, 0.0955051, 0.09548774, 0.0955219, 0.09525411, 0.09524631, 
    0.09545031, 0.09610895, 0.09643009, 0.09644343, 0.09642357, 0.09586149, 
    0.09513458, 0.09462744, 0.09467368, 0.0947077, 0.09481163, 0.09533565, 
    0.0963333, 0.09574659, 0.09456883, 0.09516189, 0.09669615, 0.09846347, 
    0.0995111, 0.09970227, 0.09957407, 0.09966083, 0.09995074, 0.09999688, 
    0.09999367, 0.09982815, 0.0989744, 0.09816942, 0.09742773, 0.09655743, 
    0.09571484, 0.0950071, 0.09399274, 0.09281535, 0.09227305, 0.09209776, 
    0.09208291, 0.09241796, 0.09298616, 0.09339474, 0.0935123, 0.09355674, 
    0.09365218, 0.09401201, 0.09429093, 0.09405444, 0.09378162, 0.09390783, 
    0.09458748, 0.09501678, 0.09552993, 0.09601219, 0.09649146, 0.09666932, 
    0.09631031, 0.09583681, 0.09534319, 0.09474345, 0.09376816, 0.09303298, 
    0.0926671, 0.09227141, 0.09130231, 0.08972041, 0.08867987, 0.08839253, 
    0.08785883, 0.08646342, 0.08469529, 0.0829534, 0.08127745, 0.08023975, 
    0.07937814, 0.07847712, 0.07670866, 0.07592357, 0.07542475, 0.0752171, 
    0.07479957, 0.07464917, 0.07463602, 0.07470063, 0.0752756, 0.07619721, 
    0.07716738, 0.07763531, 0.07722201, 0.07706822, 0.0773807, 0.07913157, 
    0.084043, 0.08588705, 0.08193773, 0.07478771, 0.06675847, 0.06077832, 
    0.05888785, 0.06114268, 0.06421143, 0.06688786, 0.06851561, 0.06887596, 
    0.06813341, 0.06779432, 0.06826209, 0.0699188, 0.07194716, 0.07361024, 
    0.074108, 0.07406018, 0.07481171, 0.07541111, 0.07604199, 0.07669666, 
    0.0772201, 0.07827725, 0.07924296, 0.07985757, 0.07986207, 0.07934539, 
    0.07888917, 0.07905762, 0.07918241, 0.07980122, 0.08093935, 0.08219214, 
    0.08307014, 0.08353719, 0.08361515, 0.08350147, 0.08326329, 0.08344629, 
    0.08400214, 0.08472607, 0.08478121, 0.08428393, 0.08455887, 0.08498191, 
    0.08596388, 0.08703528, 0.0867053, 0.08641991, 0.08674078, 0.08716416, 
    0.08765855, 0.08792145, 0.08783134, 0.08840811, 0.08876491, 0.08829068, 
    0.08752571, 0.08756805, 0.08780403, 0.08800367, 0.08805816, 0.08847464, 
    0.08823721, 0.08799388, 0.08834247, 0.08863566, 0.0882731, 0.0873671, 
    0.08651858, 0.08626604, 0.08663285, 0.08719832, 0.08755644, 0.08803823, 
    0.087983, 0.08736667, 0.08734799, 0.08841041, 0.0892816, 0.08888123, 
    0.08796892, 0.08768472, 0.08775707, 0.08740027, 0.08549173, 0.08228504, 
    0.07967659, 0.07840982, 0.079381, 0.08464764, 0.1022568, 0.1257857, 
    0.1514178, 0.15887, 0.08325969, 0.03587619, 0.02937425, 0.02610229, 
    0.02645755, 0.02530406, 0.02739497, 0.0312156, 0.03440825, 0.03641104, 
    0.03819103, 0.04048014, 0.04414225, 0.04842519, 0.05235491, 0.05628391, 
    0.05991371, 0.0628602, 0.06555031, 0.06791662, 0.0703459, 0.07230099, 
    0.07491133, 0.07771509, 0.08046828, 0.08330735, 0.08529721, 0.08704474, 
    0.08877341, 0.08970817, 0.09097635, 0.09218456, 0.0931995, 0.09404638, 
    0.09427631, 0.09432004, 0.09473765, 0.09494574, 0.09542194, 0.09584898, 
    0.09591227, 0.09607488, 0.0961618, 0.09605696, 0.09609, 0.09603713, 
    0.09588216, 0.09574585, 0.09543895, 0.09531783, 0.09543559, 0.09623075, 
    0.09691887, 0.09748652, 0.09828062, 0.0986701, 0.09894374, 0.09883436,
  0.1031936, 0.1029851, 0.1023275, 0.1014831, 0.1011543, 0.1011179, 
    0.1010242, 0.1007497, 0.1007011, 0.1008387, 0.1006777, 0.1003119, 
    0.09986497, 0.09920169, 0.09817994, 0.09715004, 0.09631265, 0.0962641, 
    0.09586731, 0.0954284, 0.09542916, 0.09568864, 0.09585084, 0.0954752, 
    0.09535499, 0.09513781, 0.09482308, 0.09510252, 0.09562333, 0.09635644, 
    0.09685527, 0.0960485, 0.09635383, 0.09669092, 0.09696946, 0.09745366, 
    0.09768816, 0.09758707, 0.09746812, 0.09738747, 0.09767038, 0.09757553, 
    0.09698089, 0.09736018, 0.09785475, 0.09816565, 0.09828524, 0.09817069, 
    0.09793028, 0.09759113, 0.0974061, 0.0973246, 0.09736148, 0.09772467, 
    0.0986746, 0.09939045, 0.09996053, 0.1008264, 0.101736, 0.1023785, 
    0.102599, 0.1026823, 0.1022593, 0.1020668, 0.1019119, 0.1019721, 
    0.1017901, 0.1015088, 0.1009828, 0.1004749, 0.09987727, 0.0989937, 
    0.0979738, 0.09709077, 0.09608252, 0.09509224, 0.09458531, 0.09418676, 
    0.09430278, 0.09472836, 0.09462172, 0.09477161, 0.0951473, 0.09527407, 
    0.09524941, 0.09534539, 0.09523088, 0.09475128, 0.09461535, 0.09500061, 
    0.09516062, 0.09499827, 0.09508544, 0.09508474, 0.09471527, 0.09400469, 
    0.09390349, 0.09411823, 0.09414003, 0.09331145, 0.09237221, 0.09179855, 
    0.09118589, 0.09015126, 0.08831524, 0.08685773, 0.08617365, 0.08569074, 
    0.08443782, 0.0825941, 0.08043136, 0.07837266, 0.07688872, 0.07616333, 
    0.07524719, 0.07410899, 0.07282111, 0.07125211, 0.07015585, 0.06920336, 
    0.06783549, 0.06732823, 0.06788542, 0.06897526, 0.07055993, 0.07170854, 
    0.07211728, 0.07263371, 0.0734849, 0.07445064, 0.07646168, 0.08167376, 
    0.08918386, 0.09200042, 0.07582452, 0.06628764, 0.06377492, 0.06066344, 
    0.05466107, 0.05366819, 0.05641648, 0.05945259, 0.06253986, 0.06487659, 
    0.06565029, 0.06626386, 0.06686625, 0.06848803, 0.07061692, 0.07272029, 
    0.07388281, 0.07387409, 0.07378466, 0.07410187, 0.07496177, 0.07590546, 
    0.07711395, 0.0779806, 0.07817683, 0.07846121, 0.07792205, 0.07711276, 
    0.0775736, 0.07803927, 0.0791546, 0.08041359, 0.08121756, 0.08140842, 
    0.08221062, 0.08265452, 0.08261601, 0.08266959, 0.08275017, 0.08309925, 
    0.0835124, 0.08332222, 0.08261178, 0.08241633, 0.08276278, 0.08341537, 
    0.08442587, 0.08515389, 0.08451561, 0.08409631, 0.08532995, 0.08654179, 
    0.08723567, 0.08719807, 0.08686998, 0.08709756, 0.08774304, 0.08772475, 
    0.08770664, 0.08805855, 0.08863916, 0.08876232, 0.08809944, 0.08785969, 
    0.08794282, 0.08846708, 0.08907062, 0.08910172, 0.08853272, 0.08792845, 
    0.08756976, 0.08778512, 0.08826671, 0.08862168, 0.08879145, 0.08920974, 
    0.08914813, 0.08960881, 0.09054005, 0.09147605, 0.09139562, 0.09053271, 
    0.08948483, 0.08884326, 0.08815209, 0.08721326, 0.08510046, 0.08206135, 
    0.07967997, 0.07856295, 0.0795188, 0.08350105, 0.09849945, 0.1254447, 
    0.1622182, 0.166753, 0.09173462, 0.04059599, 0.02826942, 0.02578347, 
    0.0248029, 0.02551026, 0.02676919, 0.02971107, 0.03255831, 0.03467054, 
    0.03716472, 0.04026932, 0.04454298, 0.04945083, 0.0536074, 0.05721096, 
    0.0603411, 0.06253909, 0.06475983, 0.06740627, 0.06983084, 0.07221203, 
    0.07513735, 0.07829095, 0.08114372, 0.08312344, 0.08475021, 0.08626867, 
    0.08801251, 0.08911408, 0.09006489, 0.09104617, 0.09201016, 0.09278612, 
    0.09339446, 0.09385663, 0.09443801, 0.09475376, 0.09507612, 0.09582657, 
    0.09636557, 0.09659602, 0.09687956, 0.09713712, 0.0973532, 0.09726942, 
    0.09718286, 0.09720697, 0.09763681, 0.0979504, 0.09881604, 0.1002919, 
    0.1014636, 0.1019849, 0.1027858, 0.103176, 0.1034102, 0.1033906,
  0.1064515, 0.1060823, 0.1053942, 0.1047048, 0.1045251, 0.1044558, 0.104067, 
    0.1038546, 0.1036617, 0.1034298, 0.1025715, 0.1019324, 0.1008265, 
    0.09970604, 0.09860425, 0.09776329, 0.09704068, 0.09639689, 0.09539986, 
    0.09497661, 0.09479834, 0.09465985, 0.09470971, 0.0949352, 0.0950744, 
    0.09542356, 0.09588772, 0.09642934, 0.09662444, 0.0968511, 0.09730342, 
    0.09737984, 0.09752264, 0.09778148, 0.09822369, 0.09885208, 0.09933176, 
    0.09919398, 0.09865232, 0.09814845, 0.09793692, 0.0977229, 0.09791488, 
    0.0988158, 0.099411, 0.1001661, 0.1006813, 0.1010538, 0.1012127, 
    0.1009056, 0.1001619, 0.09973275, 0.0996047, 0.1000677, 0.1008632, 
    0.1019731, 0.1029549, 0.1035621, 0.1038656, 0.1037703, 0.1032923, 
    0.1031029, 0.10279, 0.1027812, 0.1028405, 0.1026749, 0.1023644, 
    0.1023449, 0.1027408, 0.1029852, 0.1024687, 0.1018497, 0.1009722, 
    0.1000487, 0.09925077, 0.09855675, 0.0979876, 0.09760506, 0.09730837, 
    0.0967049, 0.09542299, 0.09470569, 0.09471889, 0.09498473, 0.09522875, 
    0.09518571, 0.09481233, 0.09447537, 0.09416284, 0.09330764, 0.09273833, 
    0.0928769, 0.09287912, 0.09243847, 0.09165923, 0.09122425, 0.0917757, 
    0.09229435, 0.09169395, 0.09033044, 0.08970851, 0.08913206, 0.08786397, 
    0.08644343, 0.08491597, 0.08406623, 0.08347377, 0.08193728, 0.07987779, 
    0.07783595, 0.0756235, 0.07365775, 0.07209583, 0.07097249, 0.07008953, 
    0.069089, 0.06738099, 0.0657901, 0.06437789, 0.06271479, 0.06154275, 
    0.06148971, 0.06244195, 0.06360768, 0.06511056, 0.06677417, 0.06797215, 
    0.06896655, 0.07052588, 0.07190644, 0.07412539, 0.08042246, 0.08896365, 
    0.1339529, 0.141304, 0.06973366, 0.05638203, 0.062353, 0.05572077, 
    0.04712097, 0.04848031, 0.05255414, 0.05694947, 0.0608555, 0.06299537, 
    0.06466027, 0.06641451, 0.06838325, 0.07071299, 0.07308355, 0.07438916, 
    0.07374257, 0.07265975, 0.07247002, 0.07323238, 0.07459164, 0.07608477, 
    0.07630806, 0.07655972, 0.07666156, 0.07595386, 0.07644682, 0.07759799, 
    0.07884704, 0.07976299, 0.08031411, 0.08018988, 0.0807325, 0.08133402, 
    0.08162224, 0.08168428, 0.08176098, 0.08226402, 0.08281987, 0.08220473, 
    0.08122252, 0.08022126, 0.0801682, 0.08060667, 0.08145218, 0.08217312, 
    0.08245341, 0.08291926, 0.08351446, 0.08495966, 0.08664458, 0.0873511, 
    0.0867968, 0.08612221, 0.08628448, 0.0869931, 0.08794535, 0.08844183, 
    0.08832433, 0.0884015, 0.08809642, 0.08760022, 0.08720584, 0.08755472, 
    0.08814745, 0.08868307, 0.08871779, 0.08832671, 0.08791514, 0.0882991, 
    0.08885501, 0.08880492, 0.08850101, 0.08872537, 0.08941416, 0.09022329, 
    0.09108359, 0.09159639, 0.09199727, 0.09141636, 0.09048351, 0.08988539, 
    0.08892315, 0.08768765, 0.08689028, 0.08511876, 0.08313663, 0.0808405, 
    0.07954992, 0.07944558, 0.08177457, 0.09168822, 0.1114117, 0.1354681, 
    0.1530843, 0.1115091, 0.04868823, 0.02942186, 0.02862966, 0.02573816, 
    0.02572985, 0.02703739, 0.02884442, 0.03106147, 0.033692, 0.03714924, 
    0.04098555, 0.04589662, 0.05144423, 0.05563278, 0.05867279, 0.06070134, 
    0.06235941, 0.06502479, 0.06719292, 0.06949814, 0.07245541, 0.07548717, 
    0.07848845, 0.0806369, 0.08234552, 0.08390832, 0.08618098, 0.08818665, 
    0.08914802, 0.08953227, 0.09047607, 0.09195542, 0.09298877, 0.09381185, 
    0.09451804, 0.09463101, 0.09475534, 0.09455846, 0.09498288, 0.09566668, 
    0.09611636, 0.09660962, 0.09675959, 0.09691557, 0.09704977, 0.09743605, 
    0.09783833, 0.09870434, 0.09979547, 0.1010992, 0.1025485, 0.1039205, 
    0.1049286, 0.1057724, 0.1060732, 0.1067925, 0.1068742,
  0.1052529, 0.1051694, 0.1051322, 0.1054614, 0.1064182, 0.1072796, 0.107411, 
    0.1069844, 0.1058513, 0.1043677, 0.1031853, 0.1016807, 0.09987183, 
    0.09839228, 0.09755302, 0.0967335, 0.09590418, 0.09496406, 0.09398929, 
    0.09304249, 0.09238733, 0.09201447, 0.09193853, 0.09216296, 0.09243609, 
    0.09340554, 0.09451057, 0.09526037, 0.09564864, 0.09600832, 0.096319, 
    0.09672701, 0.09777679, 0.09890297, 0.09966365, 0.1001515, 0.1005578, 
    0.100185, 0.09929891, 0.09884788, 0.0986855, 0.09894248, 0.09978247, 
    0.1006743, 0.1011879, 0.1016511, 0.1022023, 0.1029006, 0.1027123, 
    0.1020085, 0.1013068, 0.1008054, 0.1004928, 0.1004397, 0.1006371, 
    0.1011767, 0.1016171, 0.1011878, 0.1008347, 0.1005874, 0.1005322, 
    0.1003864, 0.09997261, 0.09994912, 0.1001803, 0.1000908, 0.1000107, 
    0.1004543, 0.1010315, 0.1010787, 0.1002728, 0.09948875, 0.09891798, 
    0.09856229, 0.09876405, 0.09911863, 0.09937787, 0.09935594, 0.09881903, 
    0.09834084, 0.09722586, 0.09609812, 0.09493624, 0.09431112, 0.0937179, 
    0.09305555, 0.09268481, 0.09242992, 0.09102175, 0.0901079, 0.08992977, 
    0.09002609, 0.0898452, 0.08923727, 0.08848131, 0.08793072, 0.08763317, 
    0.08775914, 0.08724041, 0.08646758, 0.08572852, 0.08423736, 0.08287027, 
    0.08175304, 0.08076369, 0.07992408, 0.07852241, 0.07659132, 0.07480108, 
    0.07285393, 0.07070889, 0.06896075, 0.06738167, 0.06565234, 0.06505606, 
    0.06623369, 0.06430859, 0.06092646, 0.05966797, 0.05725782, 0.0554802, 
    0.05528731, 0.05651195, 0.05821643, 0.05991443, 0.06222693, 0.06427916, 
    0.0655823, 0.06619686, 0.06691166, 0.06855982, 0.07289712, 0.0819823, 
    0.09356494, 0.1609716, 0.1302008, 0.06781556, 0.0609307, 0.06155775, 
    0.04735088, 0.04368578, 0.04762947, 0.051635, 0.05579432, 0.0592312, 
    0.06291161, 0.06557854, 0.06782064, 0.06995285, 0.07178622, 0.07300548, 
    0.07292296, 0.07248972, 0.07250204, 0.07258772, 0.07253598, 0.07326256, 
    0.07422005, 0.07472987, 0.07529038, 0.07596625, 0.07653834, 0.07744345, 
    0.0782925, 0.07851738, 0.07871681, 0.0797914, 0.08104185, 0.08140446, 
    0.08126879, 0.0812301, 0.0813075, 0.08202952, 0.0821726, 0.08107883, 
    0.07966588, 0.07865438, 0.07885614, 0.07884205, 0.07943809, 0.08058516, 
    0.08144057, 0.0824766, 0.08393764, 0.0853802, 0.08618726, 0.08665141, 
    0.08663645, 0.08636802, 0.08729843, 0.08802458, 0.08831923, 0.08802028, 
    0.08726471, 0.08705152, 0.08690619, 0.08701653, 0.08697976, 0.08729325, 
    0.08798199, 0.08817136, 0.0883285, 0.08792949, 0.08752064, 0.08759014, 
    0.0873592, 0.0864434, 0.08593104, 0.08633035, 0.08692359, 0.08787429, 
    0.08748234, 0.08685818, 0.08729523, 0.08747631, 0.0869085, 0.08649305, 
    0.08582072, 0.08562125, 0.08553182, 0.08485667, 0.08373833, 0.08217415, 
    0.08077736, 0.07943439, 0.07858645, 0.08274037, 0.09845033, 0.120726, 
    0.1402615, 0.1302348, 0.06041735, 0.03058477, 0.02723201, 0.02568763, 
    0.02530115, 0.02636037, 0.02911539, 0.03133242, 0.03434628, 0.03829387, 
    0.04244073, 0.04712678, 0.05198684, 0.05588685, 0.05862356, 0.06042261, 
    0.06234725, 0.06488024, 0.06719004, 0.07017512, 0.07367948, 0.07642858, 
    0.07846519, 0.08005885, 0.08190205, 0.08416314, 0.08652822, 0.0886599, 
    0.0895128, 0.08971217, 0.09028305, 0.0910996, 0.09158071, 0.0922189, 
    0.09293773, 0.09332018, 0.09357281, 0.09397069, 0.0945319, 0.09492112, 
    0.09510692, 0.09518865, 0.09507912, 0.09516507, 0.09540135, 0.09609109, 
    0.09742392, 0.09877497, 0.1004464, 0.1018906, 0.1028911, 0.1034264, 
    0.1037578, 0.1041128, 0.1043991, 0.1048624, 0.1051157,
  0.1043559, 0.1039006, 0.1029436, 0.1021681, 0.102027, 0.1021124, 0.1015303, 
    0.1012669, 0.1014788, 0.101576, 0.1011831, 0.1002197, 0.09859096, 
    0.09719981, 0.09599231, 0.09439225, 0.09267248, 0.09071404, 0.0890791, 
    0.08789837, 0.08711001, 0.08672254, 0.08732191, 0.08797863, 0.08866365, 
    0.08975974, 0.09113386, 0.09250326, 0.0931795, 0.09370192, 0.09436221, 
    0.09566598, 0.09750358, 0.09909033, 0.1005022, 0.1011919, 0.1014503, 
    0.1010662, 0.100757, 0.1005054, 0.1000048, 0.09971049, 0.1000975, 
    0.1005115, 0.1004259, 0.1009085, 0.1019061, 0.1025048, 0.1020804, 
    0.1007724, 0.09923429, 0.09767935, 0.09682285, 0.09705874, 0.09758688, 
    0.09804427, 0.09911548, 0.09963538, 0.09966909, 0.1000551, 0.1003647, 
    0.1001397, 0.09997647, 0.1000302, 0.09995749, 0.09970381, 0.09966332, 
    0.09985562, 0.09999532, 0.09974824, 0.09939879, 0.09841587, 0.09744329, 
    0.0965157, 0.09520593, 0.09392856, 0.09299792, 0.09287427, 0.09338405, 
    0.09423447, 0.09482435, 0.09508097, 0.09493313, 0.09458131, 0.09335749, 
    0.09166605, 0.0896119, 0.08787835, 0.0872723, 0.08714209, 0.0870674, 
    0.08670183, 0.08585837, 0.08501597, 0.08410488, 0.08304558, 0.08223712, 
    0.08187784, 0.08132572, 0.08091926, 0.08025132, 0.0786353, 0.07710732, 
    0.07589131, 0.07476074, 0.07329194, 0.07143764, 0.06996451, 0.06942269, 
    0.0677482, 0.06575849, 0.06429008, 0.0626207, 0.06032604, 0.06203784, 
    0.06659, 0.06438754, 0.05605858, 0.05135712, 0.05497998, 0.05178996, 
    0.05074969, 0.05257937, 0.05529448, 0.05778017, 0.05915312, 0.06012306, 
    0.06096733, 0.06173262, 0.06314642, 0.06531592, 0.06752499, 0.07298624, 
    0.08280866, 0.08531059, 0.122235, 0.1153603, 0.07260208, 0.05592127, 
    0.05290536, 0.04723158, 0.04587452, 0.04939336, 0.05283854, 0.05652107, 
    0.06017359, 0.06228128, 0.06370118, 0.06511221, 0.06659313, 0.0684259, 
    0.069872, 0.07074932, 0.07170022, 0.07207847, 0.07182046, 0.07247756, 
    0.07332216, 0.07394903, 0.07497715, 0.07582105, 0.07648115, 0.07715637, 
    0.07723583, 0.07766058, 0.0784276, 0.07961212, 0.08061641, 0.08048654, 
    0.08014464, 0.08011362, 0.08043487, 0.08040322, 0.07998373, 0.07942366, 
    0.07867087, 0.07824412, 0.07806697, 0.07823603, 0.07945065, 0.0811548, 
    0.08263138, 0.08364443, 0.08444269, 0.0854215, 0.08605679, 0.08598223, 
    0.08592197, 0.08608595, 0.08692395, 0.08772086, 0.08773334, 0.08672892, 
    0.0864116, 0.0865199, 0.08655588, 0.08693784, 0.0870426, 0.08729333, 
    0.08731642, 0.08717111, 0.08710904, 0.08663086, 0.08648888, 0.08663944, 
    0.08613542, 0.08619533, 0.08652955, 0.08682757, 0.08750454, 0.08777124, 
    0.08672843, 0.08626977, 0.08689885, 0.0874007, 0.08684449, 0.08528303, 
    0.08331431, 0.08179466, 0.08025091, 0.07914819, 0.07875496, 0.07833866, 
    0.07704723, 0.07523559, 0.07367146, 0.07568484, 0.0875513, 0.1066597, 
    0.1266831, 0.1214492, 0.06493197, 0.03465516, 0.02825518, 0.02844644, 
    0.02812879, 0.02754634, 0.03000611, 0.0326227, 0.03524816, 0.03899799, 
    0.04271964, 0.04701262, 0.051463, 0.05438754, 0.05687812, 0.05937037, 
    0.06197771, 0.06471971, 0.06753701, 0.07108641, 0.07470818, 0.07756282, 
    0.07934642, 0.08048446, 0.08223983, 0.08443794, 0.08658102, 0.08830007, 
    0.08898807, 0.08949687, 0.0895995, 0.08969752, 0.08994596, 0.09087923, 
    0.09232297, 0.09274466, 0.09252971, 0.09259371, 0.09317645, 0.09373663, 
    0.09422116, 0.09433512, 0.09457219, 0.09533278, 0.0962548, 0.09769382, 
    0.09923267, 0.1003732, 0.1014134, 0.1024035, 0.1030928, 0.1037707, 
    0.1041699, 0.1042951, 0.1046387, 0.1043529, 0.1042832,
  0.1048808, 0.1047617, 0.1042518, 0.1035377, 0.1023816, 0.1003675, 
    0.0966199, 0.09368556, 0.09193732, 0.09100705, 0.09131593, 0.09259554, 
    0.09364659, 0.09353951, 0.09250959, 0.0900823, 0.08700501, 0.08394171, 
    0.08136193, 0.07949591, 0.07846037, 0.07900565, 0.08011009, 0.08108332, 
    0.08237303, 0.08418754, 0.08584069, 0.08786074, 0.08983866, 0.0913877, 
    0.0926849, 0.09449408, 0.09664311, 0.09865301, 0.1007041, 0.1015624, 
    0.1012626, 0.1008825, 0.1004835, 0.09979695, 0.09863176, 0.09799389, 
    0.09804624, 0.09904706, 0.09974782, 0.1003127, 0.1006313, 0.09984033, 
    0.09839296, 0.09711805, 0.09614605, 0.09518667, 0.09462673, 0.09517401, 
    0.0959308, 0.0963093, 0.09701022, 0.09744855, 0.09759057, 0.09788598, 
    0.09822614, 0.09837365, 0.09816574, 0.0975455, 0.09674018, 0.09657395, 
    0.09643333, 0.09619242, 0.09633838, 0.09648243, 0.09634984, 0.09592266, 
    0.09574533, 0.0956547, 0.09461822, 0.09365229, 0.09278546, 0.09183517, 
    0.0904532, 0.08912825, 0.08766315, 0.08640549, 0.08611222, 0.08701718, 
    0.08792184, 0.08798351, 0.08725108, 0.08608713, 0.08541421, 0.08437525, 
    0.08289143, 0.08179474, 0.08105326, 0.08043282, 0.07899438, 0.07763522, 
    0.07680286, 0.07632462, 0.07584673, 0.07505005, 0.07363129, 0.07183931, 
    0.0704774, 0.06917679, 0.06803887, 0.06677984, 0.06568313, 0.0651083, 
    0.06398759, 0.06216236, 0.06040816, 0.05877671, 0.05661431, 0.05468797, 
    0.05903532, 0.06774233, 0.08821402, 0.07097789, 0.04221059, 0.04998564, 
    0.04772335, 0.04663793, 0.04941809, 0.05275708, 0.05493198, 0.05579012, 
    0.05647922, 0.05762505, 0.0592289, 0.06045853, 0.06236347, 0.06414872, 
    0.06507248, 0.06905304, 0.07577496, 0.07788715, 0.09243691, 0.1076553, 
    0.08228552, 0.05689548, 0.05197773, 0.04792977, 0.04851501, 0.0509438, 
    0.05437728, 0.0575651, 0.06013104, 0.06228074, 0.06369431, 0.0647646, 
    0.06654891, 0.06724291, 0.067077, 0.06748016, 0.0678836, 0.06892792, 
    0.07132713, 0.07337808, 0.07514341, 0.07553672, 0.07571952, 0.07598022, 
    0.07577056, 0.07586449, 0.07665435, 0.07699921, 0.07735547, 0.07761259, 
    0.07761753, 0.07754578, 0.07840046, 0.07919016, 0.07927502, 0.07887457, 
    0.07836883, 0.07817048, 0.07817194, 0.07841206, 0.07972226, 0.08128427, 
    0.08292749, 0.08409718, 0.08504311, 0.08516346, 0.08529022, 0.0856763, 
    0.08565236, 0.08545574, 0.08535918, 0.08604708, 0.08617072, 0.08555688, 
    0.08534684, 0.08628047, 0.08679152, 0.08668929, 0.08723789, 0.08799216, 
    0.08742232, 0.08662128, 0.08644705, 0.08636129, 0.08632512, 0.08604981, 
    0.08578192, 0.08559059, 0.08604381, 0.086731, 0.08649541, 0.08673768, 
    0.08635992, 0.0855008, 0.08528949, 0.08603333, 0.087006, 0.08712895, 
    0.08611979, 0.08437604, 0.08277648, 0.08108989, 0.07978328, 0.07808708, 
    0.0753909, 0.07092445, 0.06640546, 0.06422763, 0.06621536, 0.07824462, 
    0.1033728, 0.1160055, 0.120162, 0.06087315, 0.03841541, 0.03109176, 
    0.02856586, 0.03172616, 0.03005616, 0.03010749, 0.03327208, 0.03635944, 
    0.03878304, 0.04247433, 0.04650601, 0.05046311, 0.05311745, 0.05593539, 
    0.05865619, 0.06217188, 0.06591342, 0.06965147, 0.07331643, 0.07613213, 
    0.07841627, 0.08025671, 0.08172763, 0.08366095, 0.08535206, 0.0860928, 
    0.08610605, 0.08665948, 0.08785817, 0.08878682, 0.08901956, 0.08963924, 
    0.09050025, 0.09096177, 0.09097143, 0.09155942, 0.09220115, 0.09306311, 
    0.09408044, 0.09487908, 0.09554304, 0.09583509, 0.09618612, 0.09742577, 
    0.09925304, 0.1006054, 0.1013051, 0.1021168, 0.1026409, 0.1027712, 
    0.1030505, 0.1034117, 0.1038487, 0.1043243, 0.104601, 0.1048465,
  0.1016575, 0.1012448, 0.1004824, 0.09999525, 0.09934866, 0.09770201, 
    0.09581348, 0.09411186, 0.09244762, 0.09032816, 0.08739479, 0.08430003, 
    0.08064181, 0.07839784, 0.07800891, 0.07820418, 0.07767434, 0.07657074, 
    0.07415229, 0.07175796, 0.07077564, 0.07099993, 0.07207295, 0.07384757, 
    0.07608304, 0.07897162, 0.08161071, 0.0844209, 0.08617242, 0.08829214, 
    0.09085938, 0.09312501, 0.09539819, 0.09783816, 0.09917516, 0.09962144, 
    0.09957387, 0.09851923, 0.09721052, 0.09656531, 0.09614745, 0.09616467, 
    0.09631559, 0.0964308, 0.09584645, 0.09564212, 0.09542113, 0.09504683, 
    0.09456984, 0.0942027, 0.09383832, 0.09285445, 0.09272622, 0.09305155, 
    0.09313714, 0.09321383, 0.09344945, 0.09403027, 0.09446826, 0.09463866, 
    0.09479544, 0.09461078, 0.09415091, 0.09337664, 0.09180375, 0.09133632, 
    0.09159765, 0.09155874, 0.09138516, 0.09120147, 0.09134119, 0.09130856, 
    0.09113313, 0.09087195, 0.09024235, 0.08979971, 0.08951585, 0.08924002, 
    0.0886131, 0.0878882, 0.08689582, 0.0851455, 0.0824203, 0.08001104, 
    0.07817371, 0.07727095, 0.07826773, 0.08018421, 0.08111075, 0.08062987, 
    0.0788535, 0.07675032, 0.07489412, 0.07299016, 0.07095131, 0.06966571, 
    0.06958907, 0.06949445, 0.06875885, 0.06768437, 0.06631621, 0.06452629, 
    0.06316186, 0.06242042, 0.06187109, 0.06115131, 0.06057293, 0.05975516, 
    0.05824348, 0.05635517, 0.05453274, 0.05277749, 0.0512225, 0.05046682, 
    0.05397432, 0.05877188, 0.07377037, 0.0540522, 0.04027283, 0.04020741, 
    0.0420859, 0.04398601, 0.04745313, 0.05051496, 0.05250211, 0.05295541, 
    0.05392906, 0.05592959, 0.05762574, 0.05828022, 0.05960139, 0.06109372, 
    0.06239522, 0.06326564, 0.06464641, 0.07115206, 0.07760837, 0.09570821, 
    0.09905957, 0.05854176, 0.05601693, 0.05076209, 0.05001368, 0.04939095, 
    0.05145134, 0.0542065, 0.05747608, 0.06041011, 0.06227343, 0.062925, 
    0.06516688, 0.06693394, 0.06725395, 0.06691287, 0.06611213, 0.06625192, 
    0.06800795, 0.06975886, 0.07223064, 0.07367367, 0.07438273, 0.07510692, 
    0.07542575, 0.07569384, 0.07573905, 0.07520153, 0.07514844, 0.07499868, 
    0.07535214, 0.07638246, 0.07730024, 0.07791807, 0.07838556, 0.07826207, 
    0.07763177, 0.07768687, 0.07852839, 0.07976443, 0.08129203, 0.08300012, 
    0.08398238, 0.08361832, 0.08329757, 0.08303186, 0.08342087, 0.08458617, 
    0.08481344, 0.08484784, 0.08451004, 0.08493261, 0.08532848, 0.08540972, 
    0.08617017, 0.08735154, 0.08709648, 0.08657406, 0.08633702, 0.08608545, 
    0.08519354, 0.08420005, 0.08452667, 0.08492529, 0.08541885, 0.08529633, 
    0.08462287, 0.08455314, 0.08518384, 0.08583891, 0.08555692, 0.08484969, 
    0.08434072, 0.0840276, 0.08390664, 0.08442146, 0.08467232, 0.08425873, 
    0.08329667, 0.0820894, 0.08033976, 0.07879355, 0.07746635, 0.07567766, 
    0.0730404, 0.06918739, 0.0648877, 0.06246483, 0.06213764, 0.06817145, 
    0.08526935, 0.1046792, 0.1142608, 0.06305353, 0.03750234, 0.02873678, 
    0.02731201, 0.03033053, 0.03113335, 0.0318093, 0.03418366, 0.03647788, 
    0.03865141, 0.04240292, 0.0464298, 0.05036061, 0.05338623, 0.05688212, 
    0.06004949, 0.06511325, 0.06946008, 0.0727654, 0.07515306, 0.07745379, 
    0.08032203, 0.08243988, 0.08409344, 0.08504949, 0.08548433, 0.08529013, 
    0.08470275, 0.08524033, 0.08692883, 0.08774322, 0.08872467, 0.08936976, 
    0.08973558, 0.08946542, 0.08993103, 0.09153137, 0.09248251, 0.09340423, 
    0.09445257, 0.09491779, 0.09522337, 0.09567182, 0.0965962, 0.0980915, 
    0.09930622, 0.1001573, 0.1007732, 0.1011892, 0.1009007, 0.1002599, 
    0.1000569, 0.1003253, 0.1010439, 0.1018794, 0.1019243, 0.1017914,
  0.09660977, 0.09567353, 0.09494478, 0.09422018, 0.09313025, 0.09177291, 
    0.09076886, 0.08983535, 0.08815137, 0.08563716, 0.08313514, 0.07980895, 
    0.07562955, 0.0716288, 0.06712534, 0.06319969, 0.06188773, 0.06273939, 
    0.064191, 0.06529538, 0.06537922, 0.06501161, 0.06529768, 0.06673744, 
    0.06886729, 0.07253312, 0.07592269, 0.07919779, 0.0818314, 0.08554823, 
    0.08866104, 0.09096674, 0.09225765, 0.09385917, 0.09432085, 0.09417411, 
    0.0938348, 0.09342644, 0.0927927, 0.09300859, 0.09248219, 0.09164511, 
    0.09177746, 0.09205402, 0.09167144, 0.091481, 0.09102405, 0.09051597, 
    0.0903302, 0.08988713, 0.08922949, 0.08865686, 0.08877263, 0.08891384, 
    0.08839892, 0.08784823, 0.0878839, 0.08838137, 0.08906882, 0.08944001, 
    0.0895041, 0.08886908, 0.08852955, 0.08805725, 0.08724529, 0.08711543, 
    0.08727378, 0.08697397, 0.08669654, 0.08638109, 0.08709688, 0.08670699, 
    0.08611034, 0.08564369, 0.08501709, 0.084636, 0.0846101, 0.08417153, 
    0.08297268, 0.0821138, 0.08191179, 0.08115682, 0.07966975, 0.07872717, 
    0.07771753, 0.07568646, 0.0723763, 0.06967818, 0.06869853, 0.06913406, 
    0.07024524, 0.07023046, 0.06870341, 0.06552707, 0.0629916, 0.06209164, 
    0.06254873, 0.06230493, 0.06159604, 0.06059026, 0.05933502, 0.05698559, 
    0.0559471, 0.05585868, 0.05574984, 0.05495639, 0.05361366, 0.05231192, 
    0.05105852, 0.05035106, 0.04980325, 0.04904296, 0.04811101, 0.04728258, 
    0.04955816, 0.05105603, 0.04746997, 0.03922731, 0.03617804, 0.0366033, 
    0.03872707, 0.04188641, 0.04546362, 0.04870104, 0.05087307, 0.05208442, 
    0.05324687, 0.05506372, 0.05622339, 0.05744154, 0.05864168, 0.05923832, 
    0.05994165, 0.0615032, 0.06343409, 0.06587771, 0.07145349, 0.0745601, 
    0.06841794, 0.05488643, 0.06344981, 0.05257602, 0.05446158, 0.04963245, 
    0.050104, 0.05375773, 0.05686731, 0.05887576, 0.06030115, 0.06138483, 
    0.06310081, 0.06491087, 0.0656175, 0.06589112, 0.06596564, 0.06709974, 
    0.06937213, 0.07009717, 0.06969466, 0.06897182, 0.07010447, 0.07262652, 
    0.0749655, 0.07596301, 0.07554519, 0.07518691, 0.07441389, 0.07332245, 
    0.07386778, 0.07542512, 0.07633148, 0.07656582, 0.07664623, 0.07689379, 
    0.07740139, 0.0782728, 0.07941352, 0.08062356, 0.08158536, 0.08162528, 
    0.08089998, 0.08032635, 0.08020528, 0.08065353, 0.0816208, 0.08285707, 
    0.08327145, 0.08408743, 0.08463681, 0.08564008, 0.08569451, 0.08591321, 
    0.08668648, 0.08679623, 0.08636784, 0.08553569, 0.08450017, 0.08446812, 
    0.08454937, 0.08377817, 0.08392535, 0.08421227, 0.08428555, 0.08375657, 
    0.0837148, 0.08408292, 0.0845975, 0.084926, 0.08379474, 0.0833002, 
    0.08300089, 0.08314456, 0.08305054, 0.08220939, 0.08090792, 0.07978477, 
    0.07949767, 0.07851594, 0.07630724, 0.07411995, 0.07238759, 0.07079229, 
    0.06896629, 0.06581815, 0.0618961, 0.05972012, 0.05990234, 0.06378244, 
    0.07935536, 0.1050245, 0.1092527, 0.05136082, 0.03406808, 0.0277479, 
    0.02795392, 0.0304528, 0.0311307, 0.03222317, 0.03489354, 0.03789275, 
    0.04058728, 0.04423102, 0.04824495, 0.05263509, 0.05569297, 0.05905489, 
    0.06364797, 0.06940048, 0.07341121, 0.07674018, 0.07900207, 0.0812067, 
    0.0835132, 0.08614781, 0.08714125, 0.08717397, 0.08668986, 0.08587506, 
    0.08589356, 0.08709067, 0.08805826, 0.08895988, 0.08951356, 0.08919874, 
    0.08936131, 0.08993057, 0.09165269, 0.09320597, 0.09360091, 0.09347913, 
    0.09347397, 0.09370691, 0.09385923, 0.09444461, 0.09573914, 0.09723209, 
    0.09753493, 0.09773806, 0.09768997, 0.09705333, 0.09685157, 0.09624866, 
    0.09665041, 0.09718546, 0.09743374, 0.09770362, 0.09749351, 0.09710503,
  0.09097243, 0.09010272, 0.08918638, 0.08798145, 0.08625594, 0.0847158, 
    0.08329359, 0.08135711, 0.07909768, 0.07662567, 0.07428151, 0.07057763, 
    0.06600998, 0.06298071, 0.06072685, 0.0583999, 0.05609186, 0.05325726, 
    0.05155309, 0.05202583, 0.05399761, 0.05706125, 0.05893335, 0.0598706, 
    0.06168333, 0.06538146, 0.06984853, 0.07488052, 0.07876448, 0.08208807, 
    0.08471967, 0.08687191, 0.08774021, 0.08741954, 0.08732595, 0.08778432, 
    0.08806194, 0.08769077, 0.08649882, 0.08609973, 0.08692249, 0.08792079, 
    0.08909491, 0.08928804, 0.08883031, 0.08869064, 0.08827033, 0.08816756, 
    0.08757041, 0.08615892, 0.08472714, 0.08403009, 0.08382385, 0.08356209, 
    0.08302665, 0.08317126, 0.08288469, 0.08314312, 0.08299056, 0.08310942, 
    0.08314231, 0.08265306, 0.08234485, 0.08238943, 0.0822373, 0.08229882, 
    0.08231886, 0.08190783, 0.08222017, 0.08218612, 0.0824468, 0.08220864, 
    0.08200393, 0.08147858, 0.08104055, 0.08062957, 0.07974187, 0.07883313, 
    0.07732941, 0.07649597, 0.0763469, 0.07572271, 0.07499323, 0.0743404, 
    0.07297495, 0.07144509, 0.06975299, 0.06804789, 0.0652603, 0.06082706, 
    0.05754733, 0.05653692, 0.05687717, 0.0573754, 0.05764512, 0.05700889, 
    0.05609485, 0.05539171, 0.05488187, 0.05386989, 0.05244191, 0.05063473, 
    0.05028407, 0.05035964, 0.05012493, 0.04877369, 0.04752802, 0.0465315, 
    0.04608195, 0.0458215, 0.04549759, 0.04542098, 0.04640034, 0.04722583, 
    0.04708885, 0.04634964, 0.0463179, 0.0433266, 0.03914295, 0.03684871, 
    0.03751597, 0.04037694, 0.04400199, 0.04682408, 0.04882933, 0.05023975, 
    0.05169161, 0.05377595, 0.05523967, 0.0567822, 0.05805548, 0.05837768, 
    0.05821466, 0.05975913, 0.0621174, 0.06396568, 0.06583363, 0.06828123, 
    0.06922294, 0.06875319, 0.0831484, 0.05718783, 0.0547337, 0.05300613, 
    0.05158471, 0.05387468, 0.05598542, 0.05717695, 0.05831517, 0.0600086, 
    0.06234477, 0.06408992, 0.06429382, 0.06465344, 0.06579739, 0.06675309, 
    0.06840709, 0.06889398, 0.06935202, 0.06957946, 0.07070401, 0.07084297, 
    0.07067353, 0.07132514, 0.07263528, 0.07351506, 0.0731305, 0.07203568, 
    0.07236739, 0.07348016, 0.07458876, 0.07493845, 0.07536062, 0.07676208, 
    0.07792384, 0.07930593, 0.08000658, 0.07972288, 0.0792373, 0.07831369, 
    0.07652678, 0.07585106, 0.07835687, 0.08064085, 0.08204117, 0.08344086, 
    0.08337081, 0.08322009, 0.0845222, 0.08575459, 0.08581634, 0.08549891, 
    0.08586059, 0.085279, 0.08424104, 0.08319149, 0.08287381, 0.08379401, 
    0.08418241, 0.08397242, 0.08408901, 0.08388475, 0.08386682, 0.08332811, 
    0.08311519, 0.0830095, 0.08256255, 0.08203626, 0.08142861, 0.08089937, 
    0.08063693, 0.08046073, 0.07984339, 0.0781019, 0.07643551, 0.07566669, 
    0.075363, 0.07398048, 0.07194614, 0.0701297, 0.06836317, 0.06657917, 
    0.06462082, 0.06176312, 0.05812076, 0.05519219, 0.05469303, 0.05742316, 
    0.069823, 0.09015346, 0.1082382, 0.04848315, 0.03234425, 0.02704077, 
    0.02557584, 0.02791062, 0.03083177, 0.0356421, 0.0399116, 0.04371881, 
    0.04595926, 0.04816438, 0.0516497, 0.05543461, 0.0584091, 0.06280926, 
    0.06805262, 0.07270054, 0.0758373, 0.07856311, 0.08028988, 0.08242253, 
    0.08451438, 0.08686779, 0.08737388, 0.08724057, 0.08731854, 0.08802065, 
    0.08848449, 0.08868621, 0.08816543, 0.08862375, 0.08955508, 0.08990753, 
    0.09056257, 0.09236322, 0.09373177, 0.09413356, 0.09318163, 0.09230664, 
    0.09155399, 0.09112889, 0.09127008, 0.09207054, 0.09336013, 0.09422787, 
    0.09437867, 0.0945114, 0.09428868, 0.09355156, 0.09328783, 0.09328602, 
    0.09334381, 0.09350959, 0.09329072, 0.09321406, 0.09290144, 0.0919018,
  0.0849475, 0.08404753, 0.08267838, 0.08115455, 0.07939229, 0.07758544, 
    0.07522574, 0.07294028, 0.07036273, 0.06758594, 0.06448735, 0.0603269, 
    0.05617282, 0.05427799, 0.05262692, 0.05087641, 0.05015748, 0.04944422, 
    0.04846861, 0.04597153, 0.04331251, 0.04420101, 0.04809611, 0.05300026, 
    0.05741162, 0.06151565, 0.06610417, 0.07121264, 0.07438307, 0.07737085, 
    0.07982484, 0.08101673, 0.08120434, 0.08111706, 0.08123681, 0.08153505, 
    0.08132023, 0.08091161, 0.0812619, 0.08282104, 0.08432069, 0.0850808, 
    0.08608329, 0.08665229, 0.08652994, 0.08664285, 0.08606732, 0.08517604, 
    0.08344711, 0.08148933, 0.08035772, 0.07983626, 0.07982268, 0.07983282, 
    0.07998919, 0.07987034, 0.07933182, 0.07865628, 0.07784215, 0.07789569, 
    0.07838301, 0.07848722, 0.0783766, 0.07808888, 0.07791373, 0.07782501, 
    0.0778667, 0.0777093, 0.07799003, 0.07747624, 0.07761593, 0.07789516, 
    0.07796413, 0.0778944, 0.07695442, 0.07564554, 0.07468405, 0.07372455, 
    0.07268136, 0.07205715, 0.07162714, 0.07071663, 0.07003186, 0.06851253, 
    0.06655584, 0.06479616, 0.06295531, 0.06146652, 0.0598087, 0.05730652, 
    0.05448538, 0.05077325, 0.04737612, 0.04651807, 0.04835973, 0.05055214, 
    0.05158609, 0.05045922, 0.04875173, 0.04725783, 0.04624391, 0.0452354, 
    0.04464712, 0.04404991, 0.0435665, 0.04372785, 0.0437619, 0.04308277, 
    0.0421054, 0.04182247, 0.04206044, 0.0435359, 0.04538681, 0.04510228, 
    0.04395961, 0.04238943, 0.04463357, 0.04350134, 0.0436651, 0.04155881, 
    0.03941543, 0.03950677, 0.04243838, 0.04524701, 0.04740106, 0.04901477, 
    0.05090083, 0.05216412, 0.05357613, 0.05516503, 0.05773211, 0.05872145, 
    0.05845213, 0.05919578, 0.06101574, 0.06291988, 0.06440969, 0.06526925, 
    0.0677436, 0.07002786, 0.0879856, 0.06499833, 0.05895932, 0.05269568, 
    0.05315664, 0.05380256, 0.05503404, 0.0564198, 0.0576392, 0.05912603, 
    0.0615527, 0.06291341, 0.06271765, 0.0636003, 0.06510248, 0.06559151, 
    0.06592195, 0.06601418, 0.06665598, 0.06856308, 0.07028463, 0.07161669, 
    0.07173239, 0.06955173, 0.06741702, 0.06787565, 0.07040132, 0.07359304, 
    0.07527738, 0.07468852, 0.07387129, 0.0739091, 0.07542005, 0.07767514, 
    0.07887446, 0.07916557, 0.07871973, 0.07824952, 0.07728394, 0.07580565, 
    0.0749339, 0.07623099, 0.08002794, 0.0828356, 0.0834531, 0.08316543, 
    0.08217224, 0.08187003, 0.0839309, 0.08552367, 0.08503269, 0.08438246, 
    0.08403666, 0.08298758, 0.08197597, 0.08124875, 0.08202811, 0.08348642, 
    0.08347458, 0.08310244, 0.08302964, 0.08290442, 0.08310541, 0.0822566, 
    0.08189134, 0.08108478, 0.07980126, 0.07859965, 0.07741969, 0.07641356, 
    0.07544719, 0.07437785, 0.07379723, 0.07349994, 0.07288028, 0.07245476, 
    0.07145641, 0.06983162, 0.06811041, 0.06676418, 0.06530277, 0.06330397, 
    0.06133512, 0.05851917, 0.05458274, 0.05082867, 0.04951073, 0.05156819, 
    0.05947275, 0.0774074, 0.09072009, 0.04989616, 0.03185646, 0.03082661, 
    0.02619834, 0.02691924, 0.0309147, 0.03606096, 0.04389112, 0.04862172, 
    0.05156999, 0.05310371, 0.05588616, 0.05887249, 0.0618352, 0.06594339, 
    0.07024579, 0.07433233, 0.07704655, 0.07893602, 0.08024503, 0.08144267, 
    0.08309377, 0.08537991, 0.08647978, 0.08585993, 0.08606817, 0.08715018, 
    0.08756237, 0.08740497, 0.0870854, 0.08854473, 0.09028994, 0.09160573, 
    0.09250214, 0.09347853, 0.09335454, 0.09293936, 0.09243978, 0.09141158, 
    0.09020647, 0.0901092, 0.09034124, 0.09115089, 0.09174199, 0.09199771, 
    0.09169114, 0.09125227, 0.09021746, 0.08934315, 0.08893253, 0.08845635, 
    0.08821272, 0.08795203, 0.087655, 0.08720198, 0.08650668, 0.08564406,
  0.07722271, 0.07642183, 0.07504508, 0.07368824, 0.07175418, 0.06968913, 
    0.06742353, 0.06536022, 0.06248115, 0.05913899, 0.05473649, 0.05058029, 
    0.04751911, 0.0458152, 0.04446734, 0.04289975, 0.04253962, 0.04268413, 
    0.04226666, 0.04206443, 0.04128618, 0.04094674, 0.04119468, 0.04493441, 
    0.05220056, 0.06065689, 0.06564958, 0.06744168, 0.06868234, 0.07041777, 
    0.07209752, 0.07395075, 0.07541482, 0.07582169, 0.07548815, 0.07616618, 
    0.07666046, 0.07652324, 0.07743312, 0.07943957, 0.08073512, 0.08158176, 
    0.08320336, 0.08332283, 0.08289038, 0.08252966, 0.08160248, 0.08077921, 
    0.0789692, 0.07743204, 0.07708911, 0.07769115, 0.07761207, 0.07723949, 
    0.07673556, 0.07567174, 0.07487647, 0.07450021, 0.07412457, 0.07419129, 
    0.07432259, 0.07466231, 0.0748328, 0.07454564, 0.07403837, 0.07360753, 
    0.07341506, 0.07348901, 0.0736193, 0.07335181, 0.07332465, 0.07347605, 
    0.07364876, 0.07332321, 0.07204067, 0.07022756, 0.06916962, 0.0689041, 
    0.06846157, 0.0682131, 0.06756415, 0.06584833, 0.06393637, 0.06214784, 
    0.05987447, 0.05788986, 0.05628305, 0.05459618, 0.05296405, 0.05107098, 
    0.04880388, 0.04705559, 0.04558842, 0.04392466, 0.04170498, 0.04113057, 
    0.04292356, 0.04465836, 0.04473582, 0.04288564, 0.04154401, 0.04047982, 
    0.03982107, 0.03916403, 0.03925358, 0.03981658, 0.03971656, 0.03974001, 
    0.03954742, 0.03917035, 0.0396135, 0.04104297, 0.04318659, 0.04133756, 
    0.04126063, 0.04176069, 0.04813465, 0.05339178, 0.04781285, 0.04636665, 
    0.04193028, 0.03912099, 0.03991593, 0.04298554, 0.0462101, 0.04844694, 
    0.04966429, 0.05048419, 0.05219517, 0.05408694, 0.05689101, 0.05811473, 
    0.0584726, 0.05932946, 0.06096002, 0.06287645, 0.06365912, 0.06314308, 
    0.06352653, 0.06428477, 0.06508679, 0.05593518, 0.05617008, 0.05114882, 
    0.05214931, 0.05368159, 0.05459053, 0.05617876, 0.05740725, 0.05870784, 
    0.06039441, 0.06124526, 0.06124224, 0.06174879, 0.06241177, 0.06296282, 
    0.06333109, 0.06329178, 0.0642853, 0.06632724, 0.06797922, 0.06970056, 
    0.0698958, 0.06913964, 0.0694626, 0.06961481, 0.06946439, 0.07175997, 
    0.07460533, 0.07589106, 0.07567725, 0.07560087, 0.07708534, 0.07938244, 
    0.08011932, 0.07937139, 0.07843924, 0.0784592, 0.07779804, 0.07749583, 
    0.07754028, 0.07910214, 0.0819497, 0.08281033, 0.08245564, 0.0820396, 
    0.08132465, 0.08163613, 0.08379558, 0.0850156, 0.0848133, 0.0841372, 
    0.08313919, 0.08161179, 0.08085775, 0.08076904, 0.08152319, 0.08217123, 
    0.08226273, 0.08173047, 0.08183751, 0.08176875, 0.08190095, 0.08110667, 
    0.08012215, 0.07875939, 0.07739859, 0.0756327, 0.07389499, 0.07222909, 
    0.0700239, 0.06845383, 0.06882058, 0.06936871, 0.06986502, 0.06940742, 
    0.06782094, 0.06592172, 0.06453592, 0.06358627, 0.06220653, 0.06008536, 
    0.05810526, 0.05539298, 0.05134307, 0.04722347, 0.0447466, 0.04494606, 
    0.05219097, 0.07092249, 0.07846493, 0.04542774, 0.02510133, 0.03398706, 
    0.0287483, 0.02873345, 0.03528626, 0.04100126, 0.0450488, 0.04765913, 
    0.05355732, 0.05933696, 0.06211841, 0.06365834, 0.06446138, 0.06620824, 
    0.06901908, 0.07328413, 0.07711945, 0.07897525, 0.07926681, 0.08087118, 
    0.08233166, 0.08368769, 0.08401033, 0.0842976, 0.08496174, 0.08599571, 
    0.0866958, 0.08820774, 0.08911292, 0.09049495, 0.09109735, 0.09086405, 
    0.09157492, 0.09211335, 0.09196139, 0.09195861, 0.09103575, 0.09037776, 
    0.09017994, 0.09009644, 0.08992882, 0.08963145, 0.08956639, 0.08938162, 
    0.08850314, 0.08753351, 0.0857785, 0.08469096, 0.08392901, 0.08337053, 
    0.0826624, 0.08187149, 0.08101787, 0.08012865, 0.07934166, 0.07826101,
  0.07023544, 0.06885382, 0.06720921, 0.06534814, 0.0633698, 0.06115085, 
    0.05907097, 0.05677119, 0.05376897, 0.04999521, 0.04595699, 0.04259839, 
    0.03983187, 0.03779909, 0.03667708, 0.0364653, 0.03556585, 0.03566348, 
    0.03548701, 0.03538482, 0.03605164, 0.03834274, 0.04182617, 0.0459836, 
    0.04950938, 0.05470349, 0.06046396, 0.06367906, 0.06451631, 0.0655875, 
    0.06771818, 0.06984708, 0.07084271, 0.07125507, 0.07172504, 0.07137314, 
    0.0709473, 0.07128419, 0.07286795, 0.07574357, 0.07724618, 0.07869145, 
    0.07972421, 0.07935835, 0.0785338, 0.07826865, 0.0774614, 0.07657076, 
    0.07516599, 0.07498614, 0.07574081, 0.07628977, 0.07570487, 0.07451674, 
    0.07320349, 0.07206599, 0.07140952, 0.07149882, 0.07148906, 0.07104938, 
    0.07027781, 0.0699339, 0.07013986, 0.06994478, 0.06937068, 0.06875844, 
    0.06882333, 0.06907357, 0.06926534, 0.0689854, 0.06869456, 0.06852541, 
    0.06841619, 0.06769349, 0.06641466, 0.06541491, 0.06494546, 0.06513294, 
    0.06474688, 0.06343637, 0.06225665, 0.06069154, 0.05848727, 0.05655874, 
    0.0545158, 0.05277639, 0.05106416, 0.04946483, 0.04753385, 0.04494193, 
    0.04271924, 0.04172048, 0.04183623, 0.04195067, 0.04199992, 0.03981547, 
    0.03643275, 0.03564513, 0.03758945, 0.03895723, 0.03828655, 0.03739585, 
    0.03680074, 0.03617768, 0.03611757, 0.03637474, 0.03602713, 0.03603146, 
    0.0365159, 0.03663436, 0.0365514, 0.03672541, 0.03559422, 0.03372362, 
    0.03402193, 0.03667345, 0.04189462, 0.04830359, 0.05433666, 0.05232687, 
    0.04301395, 0.03970662, 0.03802025, 0.04142454, 0.04625695, 0.04815363, 
    0.04865111, 0.05001363, 0.05166795, 0.05295268, 0.05470516, 0.05601644, 
    0.05838574, 0.06032318, 0.06157047, 0.0620312, 0.06145896, 0.06135183, 
    0.05958357, 0.05753564, 0.05666695, 0.05400784, 0.05212419, 0.05164812, 
    0.05259966, 0.05450341, 0.05523964, 0.0565365, 0.05764972, 0.0582615, 
    0.0591814, 0.05942952, 0.05937814, 0.05936828, 0.06016916, 0.06126632, 
    0.06192649, 0.06234334, 0.06346259, 0.06446306, 0.06558809, 0.06754855, 
    0.0681073, 0.06909389, 0.07055537, 0.07268934, 0.0754248, 0.07646495, 
    0.07336411, 0.07241628, 0.0756654, 0.07901634, 0.08020309, 0.08080125, 
    0.08053721, 0.08018919, 0.08152898, 0.08248952, 0.08184025, 0.08109754, 
    0.08021974, 0.08136424, 0.0823601, 0.08189335, 0.08147887, 0.08190887, 
    0.08242994, 0.08260749, 0.08384395, 0.08427876, 0.08389372, 0.08400158, 
    0.08278257, 0.08138464, 0.08120763, 0.08107773, 0.08023985, 0.07996966, 
    0.08054458, 0.08061402, 0.0801149, 0.07960152, 0.07935684, 0.07853371, 
    0.07699304, 0.07538255, 0.07437566, 0.07322507, 0.07167345, 0.06987727, 
    0.0671903, 0.06623878, 0.06694148, 0.06700069, 0.06713825, 0.06630224, 
    0.06493194, 0.06332485, 0.06129784, 0.06038133, 0.05852766, 0.05589771, 
    0.05330696, 0.05118326, 0.04765492, 0.04333454, 0.03876887, 0.03676192, 
    0.04240471, 0.05915494, 0.06661139, 0.05922033, 0.02106018, 0.03526829, 
    0.03203103, 0.03073285, 0.03783694, 0.04538295, 0.05096617, 0.0531594, 
    0.05374767, 0.05740988, 0.06356777, 0.06528842, 0.06449814, 0.0645408, 
    0.06718042, 0.07215655, 0.07657793, 0.07880271, 0.07923146, 0.07975172, 
    0.08097292, 0.08260524, 0.0839199, 0.08498192, 0.08515375, 0.08663879, 
    0.08885434, 0.09067371, 0.09090459, 0.09033871, 0.08928143, 0.08872133, 
    0.08950545, 0.08980088, 0.08971068, 0.08906607, 0.08838293, 0.08818446, 
    0.08785816, 0.08693688, 0.08625965, 0.08624543, 0.08616079, 0.08554847, 
    0.08431493, 0.08254111, 0.08055693, 0.07894821, 0.07785474, 0.07734399, 
    0.07597134, 0.07442379, 0.0735447, 0.07279694, 0.07213561, 0.07131772,
  0.06291283, 0.06140506, 0.05930307, 0.05753453, 0.05601272, 0.05403116, 
    0.05152553, 0.04851944, 0.04501898, 0.04114662, 0.03766362, 0.03467453, 
    0.03234181, 0.0311241, 0.03182321, 0.0322375, 0.03255949, 0.0326036, 
    0.03217177, 0.03310249, 0.0339936, 0.0368659, 0.04115454, 0.04699035, 
    0.05158698, 0.05432254, 0.05483, 0.05744825, 0.06125991, 0.06315448, 
    0.0651275, 0.06683479, 0.06818601, 0.06695462, 0.06627274, 0.06597507, 
    0.06632453, 0.06773895, 0.06964992, 0.07198462, 0.07418065, 0.07547362, 
    0.07572357, 0.07537185, 0.07431024, 0.07378949, 0.07341307, 0.07282251, 
    0.0724195, 0.07293037, 0.07384485, 0.07382009, 0.07239237, 0.07017253, 
    0.06898501, 0.06789608, 0.06737877, 0.06754266, 0.06754258, 0.06676517, 
    0.06642488, 0.06583293, 0.0659263, 0.06610314, 0.066067, 0.06564569, 
    0.06596335, 0.06587442, 0.06584872, 0.06554184, 0.06458981, 0.06383094, 
    0.06319005, 0.062466, 0.06157952, 0.06149727, 0.0618835, 0.06167687, 
    0.06064466, 0.05927922, 0.05782432, 0.05641215, 0.05439695, 0.05197697, 
    0.04985309, 0.04829676, 0.0463539, 0.04462437, 0.04233457, 0.03938578, 
    0.03728221, 0.03803956, 0.03798974, 0.03734728, 0.03897993, 0.03953604, 
    0.03740773, 0.03508116, 0.0318098, 0.03137541, 0.03285549, 0.03319631, 
    0.03337953, 0.03340819, 0.03363194, 0.03340204, 0.03294702, 0.03323161, 
    0.0328468, 0.03154271, 0.03136558, 0.03038845, 0.02934268, 0.02904453, 
    0.03017602, 0.03266352, 0.0375807, 0.04174961, 0.04648653, 0.04776336, 
    0.04470874, 0.0409826, 0.037545, 0.04101574, 0.04536813, 0.04722737, 
    0.04809007, 0.04888117, 0.04986216, 0.05086978, 0.05245376, 0.05513138, 
    0.05812472, 0.06068604, 0.06108036, 0.05995626, 0.05916841, 0.05949154, 
    0.06009579, 0.05626046, 0.0530788, 0.05316966, 0.05342867, 0.05306619, 
    0.05356281, 0.05485344, 0.05524974, 0.05634784, 0.05706305, 0.05665937, 
    0.05677452, 0.05768031, 0.05797414, 0.05845304, 0.05965931, 0.06116777, 
    0.06209864, 0.06317597, 0.06422029, 0.0649998, 0.06537592, 0.06654548, 
    0.06848659, 0.07070444, 0.07223324, 0.07524708, 0.07873914, 0.07949506, 
    0.07807072, 0.07577667, 0.07436682, 0.07693561, 0.07942925, 0.07959625, 
    0.08130447, 0.08335737, 0.08509208, 0.08448729, 0.08355346, 0.08286266, 
    0.08201879, 0.08273394, 0.08288279, 0.08192986, 0.08287437, 0.08419095, 
    0.08408975, 0.08395745, 0.08449476, 0.08434779, 0.08358263, 0.08320887, 
    0.08218079, 0.08101089, 0.08074158, 0.08022905, 0.07897431, 0.0784161, 
    0.07839819, 0.07760607, 0.07656406, 0.07632769, 0.07627214, 0.07512955, 
    0.07383922, 0.07257619, 0.07163544, 0.07021936, 0.06859129, 0.06681804, 
    0.06548952, 0.0656218, 0.06595282, 0.06560177, 0.06502318, 0.06415108, 
    0.06287495, 0.0610732, 0.0587747, 0.05712978, 0.05429686, 0.05126087, 
    0.04842239, 0.04630058, 0.04317604, 0.03820593, 0.03263792, 0.02956671, 
    0.03377076, 0.04807251, 0.05264362, 0.05486443, 0.02356225, 0.03589718, 
    0.03196509, 0.03297251, 0.04023553, 0.04862014, 0.05319139, 0.05556589, 
    0.05809092, 0.06101074, 0.063366, 0.06539758, 0.06505997, 0.06396898, 
    0.0670101, 0.07178506, 0.07638099, 0.07800471, 0.07799222, 0.07907521, 
    0.08091157, 0.08241427, 0.08427305, 0.08554738, 0.08587245, 0.08704408, 
    0.08805223, 0.08827971, 0.08841044, 0.0889391, 0.08884466, 0.08849941, 
    0.08817011, 0.08752937, 0.08702868, 0.08650339, 0.08596557, 0.0849489, 
    0.08322801, 0.08213181, 0.08153185, 0.08140768, 0.0808363, 0.08020444, 
    0.0780604, 0.07587575, 0.07377147, 0.07145529, 0.07070497, 0.07012102, 
    0.06860659, 0.06738196, 0.06660115, 0.06556889, 0.06463242, 0.06391609,
  0.05646552, 0.05488382, 0.05303685, 0.05151913, 0.04986242, 0.04815671, 
    0.04535489, 0.04180434, 0.03805419, 0.03426609, 0.03094873, 0.0280635, 
    0.0255968, 0.02574733, 0.02797746, 0.03371486, 0.03416029, 0.03246179, 
    0.03366059, 0.0370671, 0.03784421, 0.03960926, 0.04196113, 0.04580785, 
    0.05018642, 0.05496043, 0.05792172, 0.05782519, 0.05746127, 0.06155952, 
    0.06319612, 0.06361862, 0.06333997, 0.06127627, 0.06031211, 0.06118312, 
    0.06303917, 0.06524941, 0.06725073, 0.06914637, 0.07205167, 0.07268833, 
    0.07115395, 0.07058477, 0.07034291, 0.07015818, 0.07032238, 0.07021037, 
    0.06998874, 0.06952503, 0.06927053, 0.06832828, 0.06643901, 0.06470852, 
    0.06401266, 0.06387284, 0.06387191, 0.06330156, 0.06259169, 0.06198689, 
    0.06134689, 0.06095939, 0.06095221, 0.06133728, 0.06178909, 0.06186989, 
    0.06235583, 0.06244259, 0.06242759, 0.06142091, 0.06044, 0.05959029, 
    0.05876683, 0.05848834, 0.0581285, 0.05814673, 0.05772922, 0.0570611, 
    0.05598725, 0.05451858, 0.05295498, 0.05189385, 0.05041442, 0.04891006, 
    0.04692652, 0.04500511, 0.04254982, 0.04024456, 0.03735356, 0.03463112, 
    0.03297187, 0.03334822, 0.03379084, 0.03233641, 0.0309325, 0.03376953, 
    0.03550357, 0.03370478, 0.0317612, 0.03025268, 0.02891058, 0.03000726, 
    0.03062974, 0.03093944, 0.03096176, 0.03098052, 0.03080782, 0.03076873, 
    0.02923195, 0.02736243, 0.02799571, 0.02615953, 0.02581712, 0.02663545, 
    0.0270407, 0.02829512, 0.03365646, 0.03931425, 0.03947297, 0.04477476, 
    0.049466, 0.04387086, 0.03857264, 0.03958718, 0.04299824, 0.04539126, 
    0.04673642, 0.04734343, 0.04836803, 0.04913374, 0.05056666, 0.05326793, 
    0.05594919, 0.0578402, 0.05773927, 0.05800405, 0.05784583, 0.05761624, 
    0.05523285, 0.05299219, 0.05306131, 0.05309838, 0.05389026, 0.05339313, 
    0.05309723, 0.05380519, 0.05451205, 0.05513908, 0.05522167, 0.05467838, 
    0.05524373, 0.0569314, 0.05816669, 0.0595905, 0.06015798, 0.06152707, 
    0.06233719, 0.06410858, 0.06578068, 0.06643952, 0.06660192, 0.0678982, 
    0.07006511, 0.0725015, 0.07435717, 0.07843043, 0.0808392, 0.08004336, 
    0.07933944, 0.08047717, 0.08027038, 0.07843748, 0.07655431, 0.08008192, 
    0.08336323, 0.08612072, 0.08677068, 0.08577277, 0.08471034, 0.08390757, 
    0.08339511, 0.08330079, 0.08232754, 0.0827355, 0.08460863, 0.08497209, 
    0.0848866, 0.08610704, 0.0863739, 0.08463264, 0.08359856, 0.08308005, 
    0.08130071, 0.07890845, 0.07713584, 0.07583447, 0.07538436, 0.07506873, 
    0.07529393, 0.07481521, 0.07406016, 0.0737973, 0.07291484, 0.0714896, 
    0.07041065, 0.06950935, 0.06818563, 0.06640259, 0.06477717, 0.06363364, 
    0.06285007, 0.06275816, 0.06292865, 0.0625569, 0.06269152, 0.06197431, 
    0.06071116, 0.05878194, 0.05564252, 0.05299602, 0.05077795, 0.04753631, 
    0.04374937, 0.04120007, 0.03861739, 0.03398795, 0.0280983, 0.02412704, 
    0.02754722, 0.03571382, 0.03931714, 0.03981484, 0.03135405, 0.04139589, 
    0.03152223, 0.03737077, 0.04464443, 0.04978801, 0.05449588, 0.05745789, 
    0.06151031, 0.0655253, 0.06791964, 0.06842314, 0.06613731, 0.06473267, 
    0.06712022, 0.07024665, 0.07290427, 0.07508208, 0.07646704, 0.07853376, 
    0.08141261, 0.08289905, 0.08422504, 0.08561922, 0.08528077, 0.08525734, 
    0.08597966, 0.08564066, 0.08601654, 0.08721187, 0.0872746, 0.08675659, 
    0.08538289, 0.0844302, 0.08316117, 0.08211531, 0.08129863, 0.07959109, 
    0.07749285, 0.0762803, 0.07529752, 0.07485148, 0.07444426, 0.0733538, 
    0.07089391, 0.06895778, 0.06746825, 0.06597507, 0.06526329, 0.06403146, 
    0.06222933, 0.06106682, 0.06019891, 0.05885177, 0.05798738, 0.05722944,
  0.05009723, 0.04825538, 0.0468139, 0.04576305, 0.04417444, 0.04281224, 
    0.04012829, 0.03618461, 0.03249981, 0.02882227, 0.02518133, 0.02219445, 
    0.01977493, 0.02066116, 0.02637091, 0.03802929, 0.03284981, 0.03635469, 
    0.04308147, 0.04973105, 0.05212095, 0.05399465, 0.05005227, 0.04617238, 
    0.04861457, 0.05306479, 0.05656699, 0.05814305, 0.05653227, 0.0593471, 
    0.05919492, 0.0581486, 0.05678073, 0.05557397, 0.05544647, 0.05688041, 
    0.05966328, 0.06177514, 0.06371703, 0.06603619, 0.06738813, 0.06701638, 
    0.06628371, 0.06606611, 0.06680671, 0.06697898, 0.06629713, 0.06612313, 
    0.06604073, 0.06539005, 0.06497761, 0.06412856, 0.0630962, 0.06221316, 
    0.061594, 0.06077827, 0.06031124, 0.0593976, 0.05808998, 0.05766927, 
    0.05737054, 0.05722351, 0.05703782, 0.05692199, 0.0570778, 0.05698805, 
    0.05705789, 0.05695986, 0.05625546, 0.05609497, 0.05561111, 0.05536083, 
    0.05470511, 0.05445923, 0.05438904, 0.05387258, 0.05270416, 0.05157828, 
    0.05074459, 0.04957616, 0.0483163, 0.04768847, 0.04677845, 0.04588646, 
    0.04431275, 0.04172751, 0.03942699, 0.03656133, 0.03308599, 0.03073754, 
    0.02947646, 0.03012263, 0.03062014, 0.0282812, 0.02563057, 0.02770988, 
    0.02956483, 0.02859677, 0.02685993, 0.02840919, 0.02750536, 0.02859866, 
    0.02864011, 0.02877109, 0.02887611, 0.02870153, 0.02878747, 0.02795907, 
    0.02578416, 0.02597679, 0.02571578, 0.02430908, 0.02478853, 0.02608556, 
    0.02550782, 0.02635323, 0.02975509, 0.03520599, 0.03789774, 0.0430024, 
    0.05135653, 0.04531474, 0.03914118, 0.0378013, 0.03996799, 0.0425605, 
    0.04425692, 0.04624663, 0.0477214, 0.04809797, 0.04939035, 0.05119885, 
    0.05318596, 0.05508868, 0.05553301, 0.05656708, 0.05601998, 0.05496029, 
    0.05397822, 0.05386559, 0.05398499, 0.05332118, 0.05329105, 0.0528404, 
    0.05273624, 0.05326969, 0.05374209, 0.05391279, 0.05407829, 0.05464447, 
    0.05594247, 0.0583231, 0.0602652, 0.06139642, 0.06241095, 0.06360831, 
    0.06456832, 0.066059, 0.06785089, 0.06861681, 0.06920738, 0.07098773, 
    0.07329702, 0.07528688, 0.07746376, 0.081077, 0.08240084, 0.08164378, 
    0.08116963, 0.08286574, 0.08310381, 0.08112949, 0.07851005, 0.08297799, 
    0.08537248, 0.08815697, 0.08903979, 0.08818282, 0.08574506, 0.08491272, 
    0.08466329, 0.08350211, 0.08279792, 0.08359611, 0.0849677, 0.08515209, 
    0.08554592, 0.08690903, 0.08573344, 0.08314839, 0.08150385, 0.08047426, 
    0.07762697, 0.07473046, 0.07308203, 0.07281506, 0.07248472, 0.07194576, 
    0.07206486, 0.07230849, 0.07184542, 0.07061134, 0.06903785, 0.06785075, 
    0.0669058, 0.06570246, 0.06418649, 0.06253438, 0.06136835, 0.06051058, 
    0.05987489, 0.05896971, 0.05785127, 0.05793422, 0.05881231, 0.05855582, 
    0.05715173, 0.05479677, 0.05119447, 0.04835059, 0.04600757, 0.04292816, 
    0.03909914, 0.03649976, 0.03429344, 0.03068315, 0.02478469, 0.02074901, 
    0.02327061, 0.02829061, 0.0302895, 0.02530064, 0.03643785, 0.0455179, 
    0.03093897, 0.03890213, 0.04890992, 0.05207647, 0.0563864, 0.05963483, 
    0.06317116, 0.06648789, 0.06841182, 0.06844728, 0.06736229, 0.06732206, 
    0.06834376, 0.06793644, 0.06986132, 0.07267211, 0.07460877, 0.07650483, 
    0.07876755, 0.08059691, 0.0819184, 0.08200856, 0.08091494, 0.08145444, 
    0.08297909, 0.08369099, 0.08475787, 0.08522282, 0.08371659, 0.0822218, 
    0.08047138, 0.07876663, 0.07729504, 0.07631664, 0.07503694, 0.07332188, 
    0.07182848, 0.070428, 0.0692529, 0.06812052, 0.06656545, 0.06464588, 
    0.06308647, 0.0618298, 0.06098982, 0.06034945, 0.05978825, 0.05857685, 
    0.0566221, 0.05545526, 0.05478361, 0.05335178, 0.05257867, 0.05183084,
  0.04434489, 0.04303698, 0.04201306, 0.04102902, 0.03916942, 0.0369927, 
    0.03452403, 0.03133078, 0.02797988, 0.02418906, 0.02058717, 0.01791774, 
    0.01625111, 0.01772723, 0.02241903, 0.02597683, 0.02250087, 0.02359114, 
    0.02628646, 0.03640921, 0.04551125, 0.06631233, 0.08539375, 0.06180593, 
    0.05006064, 0.05077011, 0.05380644, 0.05595932, 0.0543359, 0.05536061, 
    0.05400068, 0.05223833, 0.05124375, 0.05030601, 0.05081256, 0.05301802, 
    0.05519689, 0.05737836, 0.05911346, 0.05984361, 0.06025182, 0.0606863, 
    0.06165579, 0.06329238, 0.06351518, 0.0626233, 0.06189824, 0.06236318, 
    0.0634436, 0.06375823, 0.06364285, 0.0623704, 0.06140519, 0.06102259, 
    0.05982312, 0.05778624, 0.05674074, 0.05569638, 0.05442778, 0.05397409, 
    0.05413542, 0.05413748, 0.05403295, 0.05401774, 0.05369005, 0.05326863, 
    0.05289298, 0.05242087, 0.05180129, 0.052177, 0.05184121, 0.05214225, 
    0.05176319, 0.0509026, 0.05015957, 0.04957566, 0.04878448, 0.04766237, 
    0.04678546, 0.04603225, 0.0453401, 0.04532568, 0.0445031, 0.04389852, 
    0.04216198, 0.03965168, 0.037227, 0.0338737, 0.03031201, 0.02803191, 
    0.02695967, 0.02791511, 0.02759248, 0.02601346, 0.0237676, 0.02344375, 
    0.02405442, 0.02356716, 0.02182949, 0.02346784, 0.02440904, 0.02590906, 
    0.02663042, 0.02717938, 0.02712123, 0.02667532, 0.02595851, 0.02483222, 
    0.02354732, 0.0239002, 0.02401466, 0.02260133, 0.02341529, 0.02511549, 
    0.02477665, 0.02570563, 0.02735115, 0.03237943, 0.03602684, 0.03942185, 
    0.04485283, 0.04536593, 0.04193942, 0.03942534, 0.03861495, 0.04117913, 
    0.04326736, 0.04571196, 0.04787603, 0.04882874, 0.04990782, 0.05010743, 
    0.05129013, 0.0527767, 0.05409381, 0.05492714, 0.05449834, 0.05354809, 
    0.05311113, 0.05390656, 0.05535165, 0.05586438, 0.05499395, 0.05381751, 
    0.05321247, 0.05277694, 0.05325601, 0.05363061, 0.0545933, 0.0565544, 
    0.05847486, 0.06062792, 0.06213834, 0.0626214, 0.06411857, 0.06611208, 
    0.0670067, 0.06841265, 0.07010167, 0.07114403, 0.07239871, 0.07464217, 
    0.0768002, 0.07832694, 0.08025054, 0.08275412, 0.08245707, 0.08164856, 
    0.08259636, 0.08455136, 0.08437325, 0.08291161, 0.08145377, 0.08576205, 
    0.08648975, 0.08824443, 0.08836125, 0.08649766, 0.08423248, 0.08387384, 
    0.08341844, 0.08211682, 0.08218488, 0.08366906, 0.08473422, 0.08516514, 
    0.08540757, 0.08533537, 0.08352548, 0.08069175, 0.07783904, 0.07550863, 
    0.07334772, 0.07197709, 0.07094858, 0.07083288, 0.0702349, 0.06946417, 
    0.06921463, 0.06941649, 0.06859627, 0.06698796, 0.06510682, 0.06334731, 
    0.06183065, 0.06070565, 0.05969427, 0.05872708, 0.05817417, 0.05722877, 
    0.05618708, 0.05532315, 0.05458473, 0.05384159, 0.05374433, 0.0533187, 
    0.05194182, 0.04909578, 0.04565611, 0.0427313, 0.04070891, 0.03850028, 
    0.03504923, 0.03232558, 0.03073835, 0.0281161, 0.02273135, 0.01833546, 
    0.01956693, 0.02294568, 0.02302288, 0.02006494, 0.03187482, 0.04487762, 
    0.03058671, 0.0375715, 0.05407305, 0.0578569, 0.05971576, 0.06088721, 
    0.06227547, 0.06514405, 0.06643306, 0.06772323, 0.0699634, 0.07080843, 
    0.06752906, 0.06633175, 0.06797643, 0.07111686, 0.07232209, 0.07249194, 
    0.073451, 0.07516474, 0.07530151, 0.07453579, 0.07487323, 0.07718848, 
    0.08002352, 0.08244094, 0.08311007, 0.08195473, 0.07931379, 0.07682829, 
    0.07519215, 0.07346849, 0.07161348, 0.07069211, 0.06924861, 0.06786512, 
    0.06670333, 0.06573582, 0.06345691, 0.06093107, 0.05885021, 0.05725177, 
    0.0557177, 0.05449351, 0.0537771, 0.05395316, 0.05349327, 0.05259077, 
    0.05061788, 0.04920329, 0.0485587, 0.04838426, 0.04807606, 0.04641441,
  0.04046791, 0.03972591, 0.03894617, 0.03764922, 0.03529968, 0.03293922, 
    0.03057666, 0.02780556, 0.02445517, 0.02053225, 0.01715463, 0.01471442, 
    0.01446936, 0.01666714, 0.01901149, 0.0201802, 0.01720011, 0.0180404, 
    0.0211501, 0.02736978, 0.03236744, 0.04366936, 0.07023285, 0.09358442, 
    0.06636291, 0.05273835, 0.05292089, 0.05402118, 0.05168428, 0.05171654, 
    0.04973021, 0.04824969, 0.04704541, 0.04599415, 0.04690372, 0.04932515, 
    0.05069274, 0.05324045, 0.05386632, 0.05427925, 0.0555887, 0.05652783, 
    0.0586582, 0.05999026, 0.05975566, 0.05923506, 0.05834496, 0.05895472, 
    0.06012397, 0.06025216, 0.06016766, 0.0590206, 0.05852948, 0.05756428, 
    0.05571266, 0.05384781, 0.05292322, 0.05192299, 0.05065608, 0.0500562, 
    0.05051535, 0.05092486, 0.05107114, 0.05134035, 0.05106087, 0.04977807, 
    0.04918025, 0.04898929, 0.04846286, 0.04851362, 0.04839154, 0.0484996, 
    0.0482446, 0.04750378, 0.04679509, 0.04631758, 0.04591978, 0.04495284, 
    0.04379591, 0.0432937, 0.04306433, 0.04299991, 0.04224579, 0.04147092, 
    0.03979804, 0.03791215, 0.03577856, 0.0324129, 0.0290981, 0.0265103, 
    0.02555376, 0.02600791, 0.0258322, 0.02399679, 0.02248041, 0.02245699, 
    0.02218397, 0.02191707, 0.020899, 0.02122102, 0.02039796, 0.02125765, 
    0.02214237, 0.02361334, 0.02397007, 0.02313352, 0.02251844, 0.02204486, 
    0.02185898, 0.0224956, 0.02195629, 0.02074096, 0.02222914, 0.02360528, 
    0.02431563, 0.02529015, 0.02663783, 0.03116667, 0.03585432, 0.0377423, 
    0.04116587, 0.05607709, 0.04664142, 0.04286829, 0.03980561, 0.04166039, 
    0.0430022, 0.04504405, 0.0470386, 0.04790343, 0.04823763, 0.04897306, 
    0.04933326, 0.05039539, 0.05213923, 0.05264903, 0.05262973, 0.05211738, 
    0.05222617, 0.05353488, 0.05628813, 0.0577919, 0.05674966, 0.0549751, 
    0.05381008, 0.05269466, 0.053097, 0.05377642, 0.05579009, 0.05855334, 
    0.06034875, 0.06180588, 0.06256254, 0.06279182, 0.06459416, 0.06676894, 
    0.0679618, 0.06970374, 0.07182378, 0.07357176, 0.07606014, 0.07750121, 
    0.07861326, 0.08057629, 0.08306112, 0.0836952, 0.08222325, 0.08090813, 
    0.08228531, 0.08491593, 0.08510043, 0.08349283, 0.0824149, 0.08617873, 
    0.08628348, 0.08650747, 0.08421488, 0.08225904, 0.08120138, 0.08104807, 
    0.0810842, 0.08036114, 0.0802215, 0.08148499, 0.08275469, 0.08356731, 
    0.08507864, 0.08449492, 0.08117326, 0.07770313, 0.0741715, 0.07144038, 
    0.0701955, 0.06981473, 0.06952453, 0.06873029, 0.06768368, 0.06701289, 
    0.06622035, 0.06446842, 0.06361044, 0.06216269, 0.06055096, 0.05840344, 
    0.05609652, 0.05493, 0.05440679, 0.05458271, 0.05483958, 0.05398679, 
    0.05277056, 0.05238572, 0.05146147, 0.05016831, 0.04914394, 0.04792076, 
    0.04645105, 0.0440456, 0.04107119, 0.03847502, 0.03690247, 0.03506214, 
    0.032106, 0.0296691, 0.02812453, 0.0259541, 0.02063701, 0.01560741, 
    0.01598103, 0.01734561, 0.017658, 0.01598318, 0.02534452, 0.04037343, 
    0.03488794, 0.03757016, 0.05682986, 0.06147002, 0.06287482, 0.0607161, 
    0.06033128, 0.06364353, 0.06543058, 0.06871989, 0.06960709, 0.07481536, 
    0.06973985, 0.06758568, 0.06804308, 0.0670855, 0.06765879, 0.06799698, 
    0.06778548, 0.06835962, 0.06821334, 0.06960631, 0.0715284, 0.07478642, 
    0.07756142, 0.08025893, 0.07953977, 0.07723886, 0.0739549, 0.071226, 
    0.07001133, 0.06809188, 0.06590103, 0.06467571, 0.06285477, 0.06091328, 
    0.05942031, 0.0578498, 0.05516559, 0.0527919, 0.05117867, 0.05040769, 
    0.04915642, 0.04806963, 0.04708369, 0.04729633, 0.04716419, 0.04597819, 
    0.04425895, 0.04334394, 0.04318891, 0.0434239, 0.04345318, 0.04225869,
  0.03801444, 0.03693331, 0.0357765, 0.03406218, 0.03189616, 0.03025011, 
    0.02793494, 0.02493106, 0.02154191, 0.01759303, 0.0146462, 0.01275718, 
    0.01372907, 0.01526279, 0.01631864, 0.01625866, 0.01615216, 0.01663751, 
    0.01920195, 0.02384556, 0.02844699, 0.0320764, 0.04401091, 0.08130051, 
    0.09496748, 0.06312338, 0.05366001, 0.05177745, 0.04850277, 0.04762901, 
    0.04590651, 0.04457593, 0.04300296, 0.04149963, 0.04177821, 0.04363793, 
    0.04538726, 0.04831761, 0.04999032, 0.05182226, 0.05340048, 0.05482413, 
    0.05555231, 0.05565714, 0.05564762, 0.05536718, 0.05485033, 0.05474653, 
    0.05496112, 0.05500307, 0.05533165, 0.05494627, 0.05480532, 0.05378525, 
    0.05189622, 0.05031508, 0.04947857, 0.04895538, 0.04834516, 0.04736557, 
    0.04735215, 0.04766265, 0.04813104, 0.04914832, 0.04912059, 0.04807913, 
    0.0472487, 0.04670004, 0.04629073, 0.0456128, 0.0453412, 0.04506131, 
    0.04450002, 0.04432287, 0.04471658, 0.04456148, 0.04412177, 0.04310863, 
    0.04208121, 0.04197387, 0.04155358, 0.04125603, 0.04060834, 0.03967606, 
    0.03835117, 0.03655827, 0.03437927, 0.03119326, 0.02806987, 0.0250071, 
    0.02407542, 0.02383184, 0.02361655, 0.02203682, 0.02170354, 0.02184444, 
    0.02189865, 0.0217351, 0.02049001, 0.02090981, 0.01906198, 0.01887143, 
    0.01944616, 0.02068674, 0.02115911, 0.02074532, 0.02099916, 0.02109395, 
    0.02078863, 0.02139008, 0.02077153, 0.02088866, 0.02263384, 0.02350949, 
    0.02508045, 0.02634194, 0.02766141, 0.03122787, 0.03586777, 0.03814568, 
    0.03856385, 0.06160086, 0.05121303, 0.04705741, 0.04197826, 0.0418694, 
    0.04307009, 0.04538937, 0.04640681, 0.04621563, 0.04617507, 0.04760531, 
    0.04777173, 0.04851407, 0.05001158, 0.05033593, 0.04960506, 0.05016211, 
    0.05182016, 0.05289089, 0.05516123, 0.0576941, 0.05794677, 0.05650388, 
    0.05524815, 0.05340168, 0.05320315, 0.05496255, 0.05753418, 0.05989856, 
    0.06039452, 0.06121036, 0.06179073, 0.06266654, 0.06456631, 0.06632295, 
    0.06879519, 0.07183286, 0.07389954, 0.07638019, 0.0787168, 0.07930025, 
    0.08034443, 0.08318348, 0.0855357, 0.08471528, 0.08309023, 0.08185685, 
    0.0830447, 0.08557189, 0.08558641, 0.08378962, 0.08263811, 0.08512443, 
    0.0845649, 0.08309572, 0.07973988, 0.07883769, 0.07852065, 0.07881395, 
    0.0786913, 0.07866311, 0.07869224, 0.07972203, 0.08090521, 0.08247899, 
    0.08370255, 0.0819103, 0.07772419, 0.07391268, 0.07129771, 0.06940874, 
    0.06861888, 0.06807732, 0.06762657, 0.0653102, 0.06342696, 0.06232085, 
    0.06034773, 0.05858946, 0.05750163, 0.05597575, 0.05487362, 0.05322203, 
    0.0511407, 0.04981032, 0.04959395, 0.05037857, 0.05089334, 0.04997954, 
    0.04918541, 0.04876716, 0.04744974, 0.04646779, 0.04533774, 0.04387889, 
    0.04278182, 0.04116945, 0.03868508, 0.03657072, 0.03521387, 0.03348898, 
    0.03095781, 0.02841548, 0.02607672, 0.02369983, 0.01899512, 0.0140515, 
    0.01356368, 0.01346805, 0.01387773, 0.01120309, 0.02254648, 0.04290273, 
    0.04193874, 0.04405, 0.05461711, 0.06252508, 0.06253952, 0.06032073, 
    0.05803727, 0.06172846, 0.06454249, 0.06804719, 0.06956445, 0.07386719, 
    0.07830095, 0.07784571, 0.07359929, 0.06698851, 0.06354292, 0.06297375, 
    0.06244524, 0.06320654, 0.06454473, 0.06758156, 0.0706754, 0.07268862, 
    0.07449757, 0.07552392, 0.07471975, 0.07203914, 0.068454, 0.06597931, 
    0.0645676, 0.06184706, 0.0594348, 0.05768955, 0.05517516, 0.05313643, 
    0.05149586, 0.0501002, 0.04805828, 0.04636217, 0.04497568, 0.04378957, 
    0.04312261, 0.04292961, 0.04204106, 0.04154602, 0.04132384, 0.0402068, 
    0.03952423, 0.03930355, 0.03912808, 0.03959444, 0.03951573, 0.03889898,
  0.03561168, 0.03456685, 0.03334856, 0.03196467, 0.02970018, 0.02828603, 
    0.02625371, 0.02301549, 0.01912425, 0.01524964, 0.01270474, 0.01210845, 
    0.01383477, 0.01388592, 0.01314798, 0.01384266, 0.0155061, 0.017523, 
    0.02070261, 0.02579466, 0.03131165, 0.03863021, 0.05200509, 0.06604155, 
    0.1039955, 0.07683556, 0.05665555, 0.04956791, 0.0455026, 0.04413506, 
    0.04186158, 0.03908851, 0.03752442, 0.03602117, 0.03606259, 0.03795921, 
    0.04070925, 0.04418104, 0.04689618, 0.04939668, 0.05088307, 0.05221175, 
    0.05264067, 0.05277425, 0.052284, 0.05205033, 0.05206655, 0.05250084, 
    0.05263276, 0.0521108, 0.05133225, 0.05065966, 0.05050385, 0.04991328, 
    0.04855728, 0.04733396, 0.04687513, 0.04714348, 0.04664389, 0.04538513, 
    0.04539124, 0.0460869, 0.04675614, 0.04809348, 0.04825102, 0.04775947, 
    0.046774, 0.04551578, 0.04455337, 0.04298117, 0.04213685, 0.04193091, 
    0.0418952, 0.042536, 0.04363713, 0.04323598, 0.04248884, 0.04148721, 
    0.04042256, 0.04045776, 0.04103662, 0.04031654, 0.03989512, 0.03904955, 
    0.03778039, 0.03595995, 0.03311532, 0.02969847, 0.02689642, 0.02392423, 
    0.0227922, 0.02151058, 0.02122357, 0.02039175, 0.02098212, 0.02109834, 
    0.02147112, 0.02121904, 0.0200204, 0.02024334, 0.01964481, 0.0198137, 
    0.02081766, 0.02123943, 0.02167849, 0.02152132, 0.02147803, 0.02115996, 
    0.02050101, 0.02119676, 0.02062068, 0.02122799, 0.0226792, 0.02418341, 
    0.02589772, 0.02730653, 0.02917171, 0.03229078, 0.03574111, 0.03843241, 
    0.03671027, 0.05695035, 0.05284373, 0.04882844, 0.04266375, 0.04137386, 
    0.04252382, 0.04447405, 0.04510625, 0.04458484, 0.04420561, 0.04512872, 
    0.04589358, 0.04707024, 0.04858223, 0.04869254, 0.04797331, 0.04923162, 
    0.05178349, 0.05225689, 0.05353646, 0.05686268, 0.0584223, 0.05736323, 
    0.05576707, 0.05385214, 0.05388542, 0.05686777, 0.05992995, 0.06109048, 
    0.06114043, 0.0617512, 0.06205963, 0.06308626, 0.06567336, 0.06869423, 
    0.07220876, 0.07476652, 0.07630499, 0.07892647, 0.08132531, 0.08166023, 
    0.08251514, 0.08543327, 0.08681653, 0.08617797, 0.08479133, 0.08405481, 
    0.08404411, 0.08526422, 0.08441155, 0.08272433, 0.08116842, 0.08314031, 
    0.08221149, 0.07902832, 0.07712439, 0.07715587, 0.07739382, 0.0773926, 
    0.07754279, 0.07844786, 0.07955366, 0.07963304, 0.07995051, 0.07998458, 
    0.07963088, 0.07754511, 0.07408211, 0.07104973, 0.06883722, 0.06690339, 
    0.06557716, 0.06425617, 0.06291784, 0.06030788, 0.0581147, 0.05642244, 
    0.05457958, 0.05284798, 0.05130619, 0.04996267, 0.04906916, 0.04815659, 
    0.04694843, 0.04641949, 0.04674829, 0.04731417, 0.046884, 0.04583847, 
    0.04488769, 0.04443308, 0.04397603, 0.04310672, 0.04194304, 0.04060969, 
    0.040186, 0.03911919, 0.03746468, 0.03620315, 0.03487875, 0.03305429, 
    0.0304184, 0.02744344, 0.02485898, 0.02239036, 0.0184669, 0.01372283, 
    0.01261922, 0.01148909, 0.0108266, 0.007752086, 0.0161257, 0.04585078, 
    0.04234697, 0.04966583, 0.04874856, 0.05762375, 0.06107855, 0.05932807, 
    0.05738733, 0.0609698, 0.06621126, 0.06888533, 0.07250831, 0.07813696, 
    0.08363084, 0.09290542, 0.08426791, 0.07074475, 0.06118139, 0.05886712, 
    0.05873052, 0.06033977, 0.0633715, 0.06699691, 0.0699724, 0.07110511, 
    0.07207099, 0.07159481, 0.07013247, 0.06672069, 0.06299698, 0.06017376, 
    0.0587418, 0.05585678, 0.05299811, 0.05059197, 0.04828598, 0.04666345, 
    0.04592726, 0.04453994, 0.04237193, 0.04148399, 0.04044877, 0.03912216, 
    0.03835365, 0.03865179, 0.03824621, 0.03786885, 0.03795744, 0.03739479, 
    0.03682577, 0.03663252, 0.03647249, 0.03706732, 0.03710379, 0.03638629,
  0.03442005, 0.03362681, 0.03257553, 0.03085538, 0.02846509, 0.02664528, 
    0.0243247, 0.02109625, 0.01696389, 0.01311749, 0.0112826, 0.01211682, 
    0.01377901, 0.01639711, 0.01394393, 0.01438416, 0.01641477, 0.01871964, 
    0.02156846, 0.02770958, 0.03459489, 0.04184636, 0.05114914, 0.06693549, 
    0.08590247, 0.08798744, 0.06149957, 0.04825206, 0.04269538, 0.04049462, 
    0.03696923, 0.03379878, 0.03292992, 0.03175092, 0.03204667, 0.0338148, 
    0.03724299, 0.04079964, 0.04361335, 0.04585797, 0.04707728, 0.04924018, 
    0.05073616, 0.05083901, 0.04992836, 0.04928222, 0.04993642, 0.0514015, 
    0.05038707, 0.0494338, 0.04787219, 0.047787, 0.04702932, 0.04605465, 
    0.04580334, 0.04461573, 0.0443984, 0.04452821, 0.04326051, 0.04251988, 
    0.04329104, 0.04374393, 0.04390926, 0.04450012, 0.0451725, 0.04495947, 
    0.04426958, 0.04359526, 0.04285183, 0.0414776, 0.04084674, 0.04067835, 
    0.04087105, 0.04213056, 0.04382492, 0.04353068, 0.04175669, 0.0407968, 
    0.04006208, 0.04049424, 0.04111971, 0.04053669, 0.03986467, 0.03914993, 
    0.03770584, 0.03502577, 0.03206804, 0.02865496, 0.02553882, 0.02281111, 
    0.02123704, 0.01941187, 0.0192688, 0.01911195, 0.02024697, 0.02084633, 
    0.02119444, 0.02067383, 0.02018948, 0.02018778, 0.02007309, 0.02100669, 
    0.0217814, 0.02216519, 0.02320749, 0.02323467, 0.02262583, 0.02183928, 
    0.02101802, 0.0209738, 0.02099868, 0.0214445, 0.02259726, 0.02430667, 
    0.02603122, 0.02794559, 0.03100309, 0.03333884, 0.03564256, 0.03877708, 
    0.03649515, 0.04784991, 0.05335807, 0.04812131, 0.04249554, 0.04076478, 
    0.04182451, 0.04346414, 0.04380918, 0.04265701, 0.04197742, 0.04265043, 
    0.0437898, 0.04531893, 0.04671777, 0.04744532, 0.04786022, 0.04977339, 
    0.05185847, 0.05260511, 0.0540027, 0.05693339, 0.05855308, 0.05792309, 
    0.05685043, 0.05550105, 0.05605827, 0.05913027, 0.06169106, 0.06221395, 
    0.06287036, 0.06403089, 0.06469674, 0.06621175, 0.06896032, 0.07157969, 
    0.07518975, 0.07814111, 0.07986098, 0.08200852, 0.08374265, 0.08405223, 
    0.08398798, 0.0856552, 0.08599631, 0.0858373, 0.085785, 0.08500771, 
    0.08404179, 0.08284589, 0.08130142, 0.07975275, 0.07813537, 0.08009306, 
    0.07875405, 0.07604239, 0.07515381, 0.07528792, 0.07577728, 0.07705238, 
    0.07782189, 0.07848064, 0.07839844, 0.07736315, 0.07559362, 0.07455673, 
    0.07427981, 0.07292067, 0.06958365, 0.06655958, 0.06418792, 0.06163172, 
    0.06003724, 0.05909136, 0.05763299, 0.05524776, 0.05265728, 0.05114492, 
    0.04943432, 0.04783889, 0.0462809, 0.04534056, 0.04485798, 0.04383033, 
    0.04298518, 0.04297516, 0.04344577, 0.04410319, 0.04389989, 0.04286854, 
    0.04187016, 0.04100247, 0.04108113, 0.04020856, 0.0390006, 0.03851321, 
    0.03823194, 0.03789232, 0.03709248, 0.03640524, 0.0351647, 0.03319244, 
    0.03002105, 0.02675187, 0.02404969, 0.02154324, 0.01846255, 0.0144901, 
    0.01276988, 0.01065724, 0.008580913, 0.005480625, 0.009972958, 
    0.03190566, 0.04816747, 0.06303232, 0.05419995, 0.05312287, 0.05886551, 
    0.05979476, 0.05840078, 0.06132501, 0.067771, 0.06923093, 0.07001521, 
    0.07395138, 0.07620046, 0.08854299, 0.1029517, 0.07634201, 0.06059472, 
    0.05645877, 0.05674396, 0.05851787, 0.06249007, 0.06645827, 0.06939568, 
    0.07078595, 0.07088441, 0.06911128, 0.06670339, 0.06245113, 0.05757727, 
    0.05470742, 0.05338996, 0.04996698, 0.04747171, 0.04549638, 0.04394568, 
    0.04323654, 0.04225411, 0.04025894, 0.03833045, 0.03825314, 0.03767233, 
    0.0363955, 0.03648369, 0.03650692, 0.03572647, 0.03563115, 0.03594492, 
    0.03615433, 0.03536955, 0.03538787, 0.03570077, 0.03576579, 0.03564753, 
    0.03519304,
  0.03487609, 0.0336972, 0.03261575, 0.03105533, 0.02821223, 0.02529845, 
    0.02238746, 0.01872925, 0.01445663, 0.01116388, 0.009720857, 0.009897351, 
    0.01101078, 0.01529255, 0.01522771, 0.01679246, 0.01854667, 0.02107035, 
    0.02511777, 0.02937201, 0.03302105, 0.03927018, 0.04554712, 0.05563445, 
    0.07811719, 0.08251715, 0.06149194, 0.04655168, 0.03808176, 0.03470761, 
    0.03212807, 0.0302724, 0.02867968, 0.02779311, 0.02806813, 0.02991863, 
    0.03369474, 0.03767631, 0.04055323, 0.04235986, 0.04371528, 0.04599641, 
    0.04760671, 0.04832613, 0.04783401, 0.0470011, 0.0474017, 0.04804922, 
    0.04680266, 0.0456651, 0.04451391, 0.04475111, 0.04477232, 0.04398501, 
    0.04288102, 0.04194681, 0.04187828, 0.04169849, 0.04033854, 0.03978553, 
    0.03966091, 0.03889428, 0.03893502, 0.03996173, 0.04020378, 0.04063431, 
    0.04088524, 0.04064261, 0.04065864, 0.04080709, 0.0407841, 0.04017413, 
    0.03962546, 0.04101379, 0.04276475, 0.04286881, 0.04159604, 0.04121399, 
    0.04174572, 0.04173204, 0.04187519, 0.04110736, 0.04031245, 0.03910609, 
    0.03730243, 0.0337224, 0.02982446, 0.02613344, 0.02288063, 0.02039521, 
    0.01908872, 0.01743084, 0.01766446, 0.0185154, 0.01990576, 0.02049538, 
    0.02104661, 0.02080221, 0.02073409, 0.02078207, 0.02037323, 0.02122149, 
    0.02193985, 0.02340668, 0.02465681, 0.02409115, 0.02345003, 0.02263437, 
    0.02170995, 0.02145494, 0.02151441, 0.02252946, 0.02340303, 0.02527625, 
    0.02763266, 0.03030455, 0.03357549, 0.03527061, 0.03736822, 0.04025666, 
    0.03934183, 0.04707418, 0.05104423, 0.04804245, 0.04259893, 0.04108493, 
    0.04215604, 0.04305313, 0.04284781, 0.04177564, 0.0409601, 0.04147261, 
    0.04246322, 0.04419295, 0.04585146, 0.04759575, 0.04843046, 0.05034126, 
    0.05227856, 0.05427327, 0.05616039, 0.05826133, 0.05938024, 0.059822, 
    0.05950039, 0.05924181, 0.05985816, 0.06257677, 0.06450398, 0.06493065, 
    0.06598678, 0.06733546, 0.06833307, 0.06972937, 0.07257892, 0.07495366, 
    0.07829454, 0.08104306, 0.08191616, 0.08237537, 0.08334229, 0.08356382, 
    0.08363716, 0.08399043, 0.08341283, 0.08343764, 0.0845648, 0.08382331, 
    0.08213056, 0.07992245, 0.07790166, 0.07628188, 0.07509666, 0.07711942, 
    0.07576606, 0.07437709, 0.07363847, 0.07443802, 0.07618611, 0.0769593, 
    0.07717586, 0.0763042, 0.07472097, 0.07184494, 0.0694202, 0.06776974, 
    0.06725347, 0.06593344, 0.06276804, 0.06048221, 0.05741171, 0.05595075, 
    0.05513329, 0.05406914, 0.0518268, 0.04963252, 0.04795229, 0.04720241, 
    0.045673, 0.04435995, 0.04295651, 0.04195289, 0.04121154, 0.04020682, 
    0.03954157, 0.03935109, 0.03994957, 0.0406565, 0.04005292, 0.03914873, 
    0.03900115, 0.0388648, 0.03851212, 0.03798449, 0.03754424, 0.03738103, 
    0.03727164, 0.03754586, 0.037382, 0.03637135, 0.03517913, 0.03332065, 
    0.03015145, 0.02693804, 0.02411, 0.0215465, 0.01890413, 0.01577174, 
    0.01365295, 0.01114494, 0.009022705, 0.004076272, 0.007682013, 
    0.01909484, 0.04126217, 0.06917354, 0.05657956, 0.0535538, 0.05831766, 
    0.06005362, 0.0592302, 0.06190902, 0.0669781, 0.06648931, 0.06572721, 
    0.06674829, 0.06611262, 0.0908094, 0.121093, 0.08395054, 0.06126992, 
    0.05673385, 0.0571302, 0.05894173, 0.06242991, 0.06578933, 0.06774884, 
    0.06811274, 0.06643335, 0.0638365, 0.06117542, 0.0573321, 0.05230356, 
    0.04944621, 0.047587, 0.0448202, 0.04291006, 0.04149823, 0.04074167, 
    0.03977996, 0.03868364, 0.03652443, 0.03551091, 0.03568668, 0.03540586, 
    0.03478209, 0.03472901, 0.03434366, 0.03350008, 0.0332594, 0.03338157, 
    0.03410072, 0.03453421, 0.03524571, 0.03555839, 0.03559536, 0.03549613, 
    0.03537912,
  0.03494225, 0.03413526, 0.03276469, 0.03086545, 0.02765453, 0.02446694, 
    0.02060946, 0.01632937, 0.01214262, 0.009415447, 0.008231718, 
    0.008146871, 0.008969445, 0.01400861, 0.01572562, 0.01616269, 0.01826923, 
    0.02154004, 0.02695071, 0.03000444, 0.03457859, 0.04244332, 0.05043481, 
    0.0529406, 0.07568757, 0.07531705, 0.05737424, 0.04297162, 0.03392418, 
    0.03011602, 0.02827924, 0.02701639, 0.02517118, 0.02393262, 0.02305345, 
    0.02570633, 0.03158995, 0.03797583, 0.04012007, 0.04075195, 0.04167982, 
    0.04410574, 0.04566501, 0.04625212, 0.04602392, 0.04500652, 0.04499717, 
    0.04460116, 0.04382543, 0.04298698, 0.04231602, 0.04275035, 0.04247812, 
    0.04188722, 0.0404474, 0.03977852, 0.03978972, 0.03913878, 0.03816434, 
    0.03751048, 0.03703305, 0.03646916, 0.03698964, 0.03707077, 0.03809562, 
    0.03908878, 0.03905139, 0.0384812, 0.03904901, 0.04001343, 0.04027605, 
    0.03939904, 0.03884761, 0.03979616, 0.04149957, 0.042618, 0.0425391, 
    0.04239728, 0.04295286, 0.04245597, 0.04210874, 0.04120596, 0.03986002, 
    0.03805458, 0.03601154, 0.03189158, 0.02762704, 0.02351773, 0.02041936, 
    0.01829983, 0.01661205, 0.0154638, 0.01660306, 0.01832638, 0.01976022, 
    0.02046684, 0.02118146, 0.02185098, 0.02150654, 0.02152883, 0.02116729, 
    0.02207598, 0.02311792, 0.02421118, 0.02540991, 0.02561928, 0.02543656, 
    0.02457922, 0.02345804, 0.022874, 0.0228874, 0.02367638, 0.02506924, 
    0.02763859, 0.03047154, 0.03338404, 0.03674917, 0.03828327, 0.04113702, 
    0.0447215, 0.04549435, 0.05097078, 0.051483, 0.04801818, 0.04280981, 
    0.04159031, 0.04157276, 0.04204204, 0.04234241, 0.04210711, 0.04139553, 
    0.04190632, 0.04313765, 0.04454526, 0.04639598, 0.04850403, 0.04961375, 
    0.05182867, 0.0536722, 0.05630877, 0.05822663, 0.05943311, 0.06066926, 
    0.06208022, 0.06248297, 0.06301212, 0.06381489, 0.06636697, 0.06855692, 
    0.0693512, 0.07047845, 0.07113522, 0.07178667, 0.07317575, 0.0751397, 
    0.07690898, 0.07940179, 0.08088185, 0.08028308, 0.07917225, 0.08016894, 
    0.08067675, 0.0813913, 0.08203259, 0.0815295, 0.08147067, 0.08231277, 
    0.08044263, 0.07828084, 0.07614668, 0.07471662, 0.07321749, 0.07258758, 
    0.07440677, 0.07333076, 0.07293589, 0.07281289, 0.07446589, 0.07589195, 
    0.0749955, 0.0748831, 0.07318562, 0.07062708, 0.06651312, 0.06380832, 
    0.06177296, 0.06047083, 0.0577311, 0.05589325, 0.05506251, 0.05292292, 
    0.0511197, 0.04987766, 0.04798136, 0.04509214, 0.04352095, 0.04316309, 
    0.04386979, 0.04289539, 0.04137246, 0.03973521, 0.03840071, 0.03680331, 
    0.03591794, 0.03506666, 0.03512555, 0.03674206, 0.03713009, 0.03695589, 
    0.03708171, 0.03736354, 0.03754037, 0.03704602, 0.03674684, 0.03719572, 
    0.03705858, 0.03736975, 0.0377099, 0.03792165, 0.03669368, 0.03528694, 
    0.03366947, 0.03117129, 0.02837028, 0.02521441, 0.0223154, 0.02016958, 
    0.01777822, 0.01541657, 0.01217414, 0.01179791, 0.004777961, 0.00628328, 
    0.010424, 0.03090131, 0.07573604, 0.06591199, 0.05393819, 0.05756689, 
    0.05987201, 0.06031356, 0.06189371, 0.06340681, 0.06175753, 0.06246753, 
    0.06138725, 0.06954543, 0.09130528, 0.1204408, 0.09068461, 0.06385652, 
    0.05767597, 0.05817661, 0.05928103, 0.06181669, 0.06333274, 0.06284567, 
    0.06080143, 0.05820772, 0.05610896, 0.05416416, 0.05059475, 0.04638224, 
    0.04376536, 0.04262724, 0.0407913, 0.03851717, 0.03729388, 0.03647433, 
    0.03523621, 0.0348346, 0.03369462, 0.03406364, 0.03454223, 0.03440248, 
    0.0337606, 0.0333319, 0.03240811, 0.03177606, 0.03185175, 0.03188721, 
    0.03230264, 0.03338056, 0.03499518, 0.03581178, 0.03565155, 0.03577984, 
    0.03560084,
  0.03558154, 0.03488076, 0.03358192, 0.03111119, 0.02733549, 0.02332893, 
    0.01905792, 0.01460956, 0.01085647, 0.008841584, 0.007937008, 
    0.008086857, 0.009182272, 0.01627027, 0.01761532, 0.01654336, 0.01841502, 
    0.02206286, 0.02587363, 0.02881414, 0.03542686, 0.04350714, 0.04940569, 
    0.05176781, 0.07292183, 0.06837657, 0.05440993, 0.04148966, 0.0320981, 
    0.02743282, 0.02533627, 0.02484295, 0.02345164, 0.02083196, 0.01923905, 
    0.02335198, 0.03619158, 0.04276586, 0.04322449, 0.04190343, 0.04160034, 
    0.04220885, 0.04298314, 0.04310053, 0.04310882, 0.04234978, 0.04244211, 
    0.04225248, 0.04216668, 0.04213675, 0.04168108, 0.04123785, 0.03982323, 
    0.03910709, 0.03816355, 0.03801468, 0.03725572, 0.03576051, 0.03542472, 
    0.03558217, 0.0348735, 0.03510118, 0.0356442, 0.03587621, 0.03771058, 
    0.0396671, 0.03969909, 0.03906544, 0.03844436, 0.03910193, 0.03916896, 
    0.03893303, 0.03850943, 0.03905877, 0.04067251, 0.04202942, 0.04230472, 
    0.04228706, 0.04234417, 0.0420115, 0.04155526, 0.04044804, 0.03909078, 
    0.03715088, 0.03461162, 0.03054341, 0.02670201, 0.02243219, 0.01926347, 
    0.01703096, 0.01501029, 0.01464694, 0.01598404, 0.01832532, 0.01990249, 
    0.02092683, 0.02179827, 0.02298348, 0.02270221, 0.02212188, 0.02192651, 
    0.02310994, 0.02372397, 0.02519413, 0.02798401, 0.02795354, 0.0273648, 
    0.02689658, 0.02592593, 0.02492367, 0.02484542, 0.02546208, 0.02662771, 
    0.02898123, 0.03250099, 0.03685423, 0.03991603, 0.04057499, 0.04554465, 
    0.05006269, 0.0493397, 0.05219673, 0.05048316, 0.04636265, 0.04292481, 
    0.04196671, 0.04121812, 0.04163632, 0.04222786, 0.04270436, 0.04205488, 
    0.04359479, 0.04530986, 0.04577846, 0.04664819, 0.04897879, 0.05096344, 
    0.05319334, 0.05441479, 0.05610786, 0.05806148, 0.05950466, 0.06180892, 
    0.06412925, 0.064914, 0.06581875, 0.06795441, 0.07096719, 0.07281654, 
    0.07400217, 0.07512346, 0.07593931, 0.07665633, 0.07739225, 0.0774144, 
    0.07804448, 0.07811908, 0.07763387, 0.07753102, 0.07743918, 0.07831211, 
    0.07846291, 0.07894453, 0.07994729, 0.08066389, 0.08009083, 0.07884135, 
    0.07637465, 0.07353712, 0.07215352, 0.07159439, 0.07070173, 0.07184777, 
    0.07329945, 0.07281225, 0.07252177, 0.07272138, 0.07358514, 0.07347745, 
    0.07247715, 0.07093536, 0.06791981, 0.06513877, 0.06208213, 0.05892645, 
    0.0564326, 0.05437497, 0.05229034, 0.05112859, 0.04933969, 0.04768731, 
    0.04563612, 0.04373178, 0.04247221, 0.04046054, 0.03925088, 0.03908675, 
    0.0393232, 0.03867966, 0.03724254, 0.03577599, 0.03457525, 0.03321953, 
    0.03206468, 0.03210272, 0.03272031, 0.0333771, 0.03354099, 0.03442132, 
    0.03563227, 0.03626871, 0.0357551, 0.03573145, 0.03604301, 0.03696651, 
    0.03768202, 0.03831411, 0.03895354, 0.03920119, 0.0380979, 0.03651739, 
    0.03465786, 0.03270736, 0.02992461, 0.02675663, 0.02406333, 0.02217263, 
    0.02001272, 0.01739822, 0.01398686, 0.01480752, 0.004242166, 0.004564054, 
    0.008012953, 0.02419527, 0.07062174, 0.07173765, 0.05476138, 0.0566819, 
    0.05965099, 0.05995691, 0.05847014, 0.05816573, 0.05756883, 0.05758441, 
    0.05662184, 0.06295866, 0.07714127, 0.1203882, 0.1015889, 0.07162353, 
    0.06303205, 0.05864671, 0.05714599, 0.05861101, 0.05844821, 0.05672165, 
    0.05505235, 0.05292417, 0.05038758, 0.04652529, 0.04340162, 0.0411401, 
    0.0394123, 0.03875333, 0.03686011, 0.03470916, 0.03402134, 0.03320495, 
    0.03193418, 0.03122469, 0.03142591, 0.03288196, 0.03345177, 0.03269525, 
    0.03209829, 0.03217029, 0.03219197, 0.03204974, 0.03146764, 0.03147818, 
    0.03198072, 0.03324131, 0.03462049, 0.03509431, 0.03564085, 0.03565482, 
    0.03562481,
  0.03661818, 0.03610699, 0.03464264, 0.03152805, 0.02718258, 0.02257165, 
    0.01783468, 0.01365247, 0.01081194, 0.009435712, 0.008701481, 
    0.008816324, 0.01016351, 0.01712661, 0.0187149, 0.01807991, 0.01944946, 
    0.02230396, 0.02523553, 0.02743341, 0.03386659, 0.03836412, 0.04214765, 
    0.04750035, 0.05776094, 0.05786961, 0.04872606, 0.0403328, 0.03274025, 
    0.02680272, 0.02384955, 0.02304696, 0.02180673, 0.01869916, 0.01840731, 
    0.02914157, 0.04501292, 0.06628891, 0.04841316, 0.04325769, 0.03976252, 
    0.03839215, 0.03876303, 0.03878652, 0.03934674, 0.03973638, 0.03975606, 
    0.03910443, 0.0392371, 0.04028152, 0.04019758, 0.03948566, 0.03781865, 
    0.03684208, 0.03595424, 0.0353304, 0.03400358, 0.03328775, 0.03329848, 
    0.03305791, 0.03342054, 0.03453164, 0.03539313, 0.03573446, 0.03736733, 
    0.03862512, 0.03837952, 0.03835443, 0.03886097, 0.03864519, 0.03835129, 
    0.03842896, 0.03907085, 0.03984156, 0.04075452, 0.04112814, 0.04164611, 
    0.04196738, 0.0425215, 0.0415156, 0.04003797, 0.03873553, 0.03751634, 
    0.03609946, 0.0336501, 0.02995694, 0.02636629, 0.02167919, 0.01877888, 
    0.01606914, 0.01385945, 0.01426285, 0.01654022, 0.01947238, 0.02053629, 
    0.0218094, 0.02266402, 0.02369889, 0.02334332, 0.02238454, 0.02268946, 
    0.02349312, 0.02439695, 0.02691068, 0.02832233, 0.0289965, 0.02992582, 
    0.03009332, 0.0292216, 0.02761761, 0.02752206, 0.02736507, 0.0279431, 
    0.03043793, 0.03419522, 0.03868062, 0.04066115, 0.04436246, 0.04999089, 
    0.05138075, 0.05220305, 0.05236077, 0.04851396, 0.0450956, 0.04329681, 
    0.04299818, 0.04254793, 0.04261206, 0.04226303, 0.04176564, 0.04108965, 
    0.04371313, 0.04544603, 0.04620255, 0.04769906, 0.04988381, 0.05211025, 
    0.0536872, 0.05491089, 0.0567494, 0.05859331, 0.0593341, 0.06217356, 
    0.06565176, 0.06738631, 0.06924583, 0.07174928, 0.07510361, 0.07680914, 
    0.07748327, 0.07840085, 0.08025114, 0.08057831, 0.07974413, 0.07916972, 
    0.07853581, 0.07643383, 0.07485916, 0.07544513, 0.07692547, 0.0778577, 
    0.07720363, 0.07670978, 0.07742328, 0.07795426, 0.07614138, 0.07364187, 
    0.07154679, 0.07000848, 0.06955331, 0.06973027, 0.06926797, 0.07120857, 
    0.072364, 0.07200016, 0.0713691, 0.07068215, 0.0698545, 0.06892207, 
    0.06737833, 0.06441624, 0.0608211, 0.05842441, 0.05627393, 0.0534979, 
    0.0508341, 0.04906655, 0.04714153, 0.0446506, 0.04169104, 0.04046738, 
    0.03957225, 0.03804595, 0.03677464, 0.03567936, 0.03474913, 0.034469, 
    0.03411343, 0.0332316, 0.03200389, 0.03100551, 0.03086245, 0.03064436, 
    0.03032404, 0.03063304, 0.03140629, 0.03213818, 0.03331046, 0.03456629, 
    0.03466548, 0.03481216, 0.0351854, 0.03593265, 0.03679639, 0.03823601, 
    0.03968722, 0.04054468, 0.04151723, 0.04191847, 0.04105761, 0.03931274, 
    0.03688706, 0.03498523, 0.03211927, 0.02883828, 0.02635863, 0.02460518, 
    0.02207961, 0.01902525, 0.01557068, 0.01240066, 0.002992814, 0.003332006, 
    0.005936498, 0.01444095, 0.06969758, 0.07839755, 0.05820132, 0.05648871, 
    0.05920576, 0.05789169, 0.05545053, 0.0555388, 0.05363466, 0.05441976, 
    0.0545994, 0.05719116, 0.06474774, 0.1000613, 0.1098802, 0.09432685, 
    0.08176807, 0.06923286, 0.05969993, 0.05712594, 0.05431402, 0.05202195, 
    0.05121934, 0.04936983, 0.04523481, 0.04145259, 0.03881222, 0.03687833, 
    0.03588938, 0.03493378, 0.03308297, 0.03084722, 0.03060886, 0.03078493, 
    0.02974828, 0.02908435, 0.02998382, 0.03112876, 0.03052526, 0.02974213, 
    0.03067171, 0.03101251, 0.03074351, 0.03087068, 0.03076956, 0.03108648, 
    0.03177088, 0.03278818, 0.03396202, 0.03520599, 0.03607091, 0.03674975, 
    0.03662799,
  0.03848476, 0.03743365, 0.03521763, 0.03183668, 0.02751298, 0.02237192, 
    0.01765375, 0.01401923, 0.01193771, 0.01113136, 0.01143246, 0.01152168, 
    0.01331884, 0.019068, 0.02146517, 0.02142563, 0.0221157, 0.02410303, 
    0.02707832, 0.02803737, 0.03010341, 0.03564378, 0.03658324, 0.04579053, 
    0.05395563, 0.05159913, 0.04455269, 0.03752987, 0.03311162, 0.02703949, 
    0.02430612, 0.02259479, 0.02081708, 0.01776644, 0.02035602, 0.03265831, 
    0.05227916, 0.09559172, 0.05358304, 0.04366489, 0.03723012, 0.03507854, 
    0.03478602, 0.03405685, 0.0354635, 0.03661876, 0.03649798, 0.03548026, 
    0.03553632, 0.03672716, 0.03803676, 0.03832223, 0.03714371, 0.03577981, 
    0.03399964, 0.03315005, 0.03253773, 0.03303493, 0.03299546, 0.03261981, 
    0.03298745, 0.03382845, 0.03475017, 0.03512706, 0.03575888, 0.03705524, 
    0.03668379, 0.03732322, 0.03919735, 0.03931496, 0.03890013, 0.03984365, 
    0.04086878, 0.04140911, 0.04126583, 0.04137847, 0.04211497, 0.04271875, 
    0.04205639, 0.04091892, 0.03991571, 0.03848622, 0.03715368, 0.03589042, 
    0.03356339, 0.03038515, 0.02651163, 0.02224129, 0.01818046, 0.01449793, 
    0.01269895, 0.01391825, 0.01717727, 0.02027287, 0.02157065, 0.02258207, 
    0.02322681, 0.02352848, 0.02302357, 0.02203046, 0.02283399, 0.02359234, 
    0.02526238, 0.02765633, 0.02874865, 0.03092813, 0.03170231, 0.03211265, 
    0.03226686, 0.0309223, 0.03035911, 0.03027856, 0.03098243, 0.03243114, 
    0.03481818, 0.0386407, 0.04214195, 0.0479878, 0.05207578, 0.05242042, 
    0.05075089, 0.04995792, 0.04664798, 0.04437511, 0.04404495, 0.04439596, 
    0.04329746, 0.04225313, 0.04150037, 0.04082229, 0.04016254, 0.042145, 
    0.04487952, 0.04756685, 0.04936912, 0.05154349, 0.0540096, 0.05612905, 
    0.05776589, 0.0590869, 0.06046819, 0.06122251, 0.0637373, 0.06755657, 
    0.07103612, 0.073978, 0.07561496, 0.07716762, 0.07755505, 0.078334, 
    0.07969206, 0.08089703, 0.08096327, 0.07958168, 0.0788052, 0.07725927, 
    0.07505217, 0.07352918, 0.07411428, 0.07507401, 0.07497679, 0.07353851, 
    0.07296859, 0.07312634, 0.07265177, 0.07101311, 0.06882647, 0.06646891, 
    0.06604084, 0.06703737, 0.06723642, 0.06699532, 0.07014745, 0.07180004, 
    0.07083962, 0.06858716, 0.06623965, 0.06373652, 0.06233124, 0.06049686, 
    0.05713922, 0.05404563, 0.052192, 0.04951218, 0.04673528, 0.0444504, 
    0.0424157, 0.04029383, 0.03738466, 0.03540229, 0.03493252, 0.03397374, 
    0.03258585, 0.03140558, 0.0313695, 0.03126789, 0.03075457, 0.03010555, 
    0.02961488, 0.02873375, 0.02812612, 0.02805133, 0.02842501, 0.0290192, 
    0.02984835, 0.0307408, 0.03169374, 0.03346449, 0.0344987, 0.03440674, 
    0.03423441, 0.0353127, 0.03714433, 0.03919871, 0.04154006, 0.04350676, 
    0.0445788, 0.0456443, 0.0454872, 0.04445527, 0.04270328, 0.04031278, 
    0.0380937, 0.03500924, 0.03178976, 0.02910227, 0.02707295, 0.02444829, 
    0.02115893, 0.01724496, 0.01403852, 0.004365588, 0.002598457, 
    0.004766081, 0.009797481, 0.05630038, 0.09270681, 0.06119815, 0.05776504, 
    0.05768934, 0.05548152, 0.05373901, 0.05272517, 0.04943731, 0.05119179, 
    0.05195929, 0.05235254, 0.05806495, 0.0694306, 0.08612703, 0.09940236, 
    0.1010736, 0.09328756, 0.07448779, 0.06222474, 0.05351101, 0.04911202, 
    0.04732018, 0.04474406, 0.04098004, 0.03776434, 0.03490607, 0.03249191, 
    0.03157476, 0.03034907, 0.02888872, 0.02773374, 0.02790911, 0.02802465, 
    0.02768004, 0.02724499, 0.02760468, 0.02798922, 0.0280863, 0.02824942, 
    0.02931247, 0.02964188, 0.02949443, 0.02945401, 0.02992775, 0.0310078, 
    0.03210905, 0.03401067, 0.03536615, 0.03691806, 0.03766481, 0.03864904, 
    0.03873218,
  0.04028976, 0.038646, 0.03621881, 0.03259465, 0.02776799, 0.0226165, 
    0.01842918, 0.01514432, 0.01357067, 0.01386704, 0.01527764, 0.01505473, 
    0.01697842, 0.0229812, 0.02634753, 0.02539769, 0.02479811, 0.02596377, 
    0.02944238, 0.02915762, 0.02937145, 0.03959797, 0.04191358, 0.04316095, 
    0.05315269, 0.05506762, 0.04489816, 0.03704993, 0.03196188, 0.02696973, 
    0.02468247, 0.0230367, 0.02079199, 0.01862499, 0.02240949, 0.03456271, 
    0.05019665, 0.09864617, 0.06123163, 0.04453077, 0.03509985, 0.03261838, 
    0.03104546, 0.03118475, 0.03281805, 0.0340697, 0.03428435, 0.03330547, 
    0.0334132, 0.03430296, 0.03566382, 0.03684237, 0.03662015, 0.03543936, 
    0.03376326, 0.03325166, 0.03364448, 0.03385044, 0.03377163, 0.03320186, 
    0.03332165, 0.03403426, 0.03438438, 0.03390907, 0.03425327, 0.03529169, 
    0.03542462, 0.03635954, 0.03859567, 0.03953825, 0.03931488, 0.04082987, 
    0.04187851, 0.04183038, 0.04202016, 0.04262282, 0.04315021, 0.04289394, 
    0.04215268, 0.04186522, 0.04105186, 0.03952451, 0.03783966, 0.03620952, 
    0.03368371, 0.03076205, 0.02615115, 0.02132738, 0.01688299, 0.01299473, 
    0.01132745, 0.01314061, 0.01650456, 0.01969431, 0.02176372, 0.02301378, 
    0.02280582, 0.02209545, 0.02203447, 0.02190957, 0.02320325, 0.02459593, 
    0.02719169, 0.02906372, 0.03075623, 0.03297628, 0.03383196, 0.03389376, 
    0.03326019, 0.03220251, 0.03242361, 0.03184157, 0.032187, 0.0333683, 
    0.03527654, 0.0390116, 0.04440171, 0.04984995, 0.05198995, 0.0524097, 
    0.05018027, 0.04730217, 0.04426716, 0.04341671, 0.04324597, 0.04338042, 
    0.04128829, 0.04049144, 0.04040397, 0.03970491, 0.03922709, 0.0417542, 
    0.04476995, 0.05029973, 0.05221424, 0.05367384, 0.05646154, 0.05855903, 
    0.06024832, 0.06236652, 0.06378359, 0.06463248, 0.06762025, 0.07189824, 
    0.07491825, 0.07645696, 0.07719115, 0.07721315, 0.07586969, 0.076345, 
    0.07797502, 0.07866675, 0.07903242, 0.07826058, 0.07774161, 0.07692449, 
    0.07528166, 0.0735027, 0.07258578, 0.07177079, 0.0698377, 0.06841808, 
    0.06797775, 0.0677414, 0.06761204, 0.06549062, 0.06309641, 0.06165051, 
    0.06243519, 0.06347894, 0.06314573, 0.06367501, 0.06716342, 0.06776683, 
    0.06524077, 0.06160669, 0.0587987, 0.05680491, 0.05427681, 0.05234139, 
    0.05014987, 0.0478134, 0.04508337, 0.04260444, 0.0405644, 0.03856136, 
    0.0369474, 0.03495636, 0.03240768, 0.03143027, 0.03112718, 0.0300461, 
    0.02866858, 0.02812207, 0.0284035, 0.02816357, 0.02778154, 0.02798572, 
    0.02764904, 0.0270492, 0.02630621, 0.0261385, 0.02706923, 0.02847386, 
    0.02931699, 0.03071713, 0.03231655, 0.03367521, 0.03472668, 0.03585567, 
    0.03715253, 0.03869382, 0.04081872, 0.04338728, 0.04561589, 0.04761343, 
    0.04931894, 0.04993666, 0.0492166, 0.04802803, 0.04612179, 0.04367947, 
    0.04101725, 0.03759952, 0.03468793, 0.03200628, 0.02951538, 0.0267453, 
    0.02382556, 0.01929851, 0.01507323, 0.007193554, 0.003293367, 
    0.006602765, 0.01435018, 0.05108481, 0.09294926, 0.06582335, 0.05734075, 
    0.05552851, 0.05300759, 0.050044, 0.04816326, 0.04615257, 0.04963334, 
    0.04989501, 0.04960303, 0.05139494, 0.05536118, 0.06074752, 0.06503028, 
    0.08315442, 0.1014807, 0.09263853, 0.07615501, 0.05889408, 0.04824818, 
    0.04342103, 0.04002608, 0.03680445, 0.03397757, 0.03117981, 0.02883738, 
    0.02776285, 0.02617534, 0.02513342, 0.02480072, 0.02453503, 0.02488074, 
    0.02541814, 0.02489298, 0.02518198, 0.02556166, 0.02631113, 0.02760179, 
    0.02852197, 0.0289121, 0.02854528, 0.02884011, 0.03010722, 0.03209128, 
    0.03402897, 0.03595295, 0.03761375, 0.03910172, 0.03974963, 0.04087928, 
    0.04126241,
  0.04155755, 0.03963783, 0.03676788, 0.03246231, 0.02755335, 0.02290317, 
    0.01892925, 0.01614955, 0.0153475, 0.0168688, 0.01769772, 0.01662633, 
    0.01961027, 0.02591334, 0.02804535, 0.02719978, 0.0271625, 0.02848984, 
    0.02985434, 0.0295117, 0.02853999, 0.03542211, 0.04521818, 0.05373802, 
    0.05981304, 0.05871317, 0.04984849, 0.03851438, 0.0307772, 0.02615522, 
    0.0236186, 0.02233323, 0.02076735, 0.01912225, 0.02217539, 0.03435904, 
    0.04267579, 0.1054762, 0.07803337, 0.04637302, 0.03424248, 0.03082314, 
    0.02881458, 0.0281226, 0.03083628, 0.03263747, 0.03281035, 0.03182388, 
    0.03223705, 0.03313947, 0.03354222, 0.03460943, 0.03547946, 0.03479402, 
    0.03374644, 0.03413063, 0.03462465, 0.03398942, 0.03399271, 0.03415924, 
    0.03438707, 0.03411851, 0.03381561, 0.03311484, 0.03344589, 0.0346565, 
    0.03528598, 0.03631052, 0.03790696, 0.03881345, 0.03984272, 0.04069249, 
    0.04131096, 0.0417341, 0.04295086, 0.04310378, 0.04263612, 0.04210968, 
    0.04172464, 0.04204646, 0.04138012, 0.03997834, 0.03826456, 0.036473, 
    0.03410667, 0.03053459, 0.02566634, 0.02027483, 0.01572796, 0.01245111, 
    0.01119644, 0.01189834, 0.01477886, 0.01767004, 0.01940405, 0.01984067, 
    0.01981487, 0.02020857, 0.02152472, 0.02305696, 0.02429327, 0.02644335, 
    0.02842029, 0.03010392, 0.03263312, 0.03377982, 0.03467181, 0.03378592, 
    0.03325905, 0.03321126, 0.0329779, 0.03127689, 0.03310031, 0.03472836, 
    0.03664081, 0.04096853, 0.04796053, 0.04870837, 0.0519194, 0.05127279, 
    0.04441672, 0.04149514, 0.04098314, 0.04124954, 0.04118371, 0.04086084, 
    0.03973563, 0.03986507, 0.04102153, 0.03999643, 0.04000472, 0.03960148, 
    0.04431047, 0.05355876, 0.05451285, 0.05534474, 0.05769902, 0.05990212, 
    0.06244895, 0.06453353, 0.06693432, 0.06993095, 0.07433824, 0.07688506, 
    0.07646511, 0.07525246, 0.07578892, 0.07629051, 0.07540859, 0.07542592, 
    0.07561097, 0.07603493, 0.07718431, 0.07728845, 0.07633819, 0.07537752, 
    0.07418618, 0.07186028, 0.06940091, 0.06738647, 0.06580456, 0.06445061, 
    0.06349698, 0.06262477, 0.06244396, 0.06069013, 0.05812285, 0.05757632, 
    0.05860009, 0.05917966, 0.05935371, 0.05995999, 0.0616174, 0.05974993, 
    0.05570116, 0.05264859, 0.05085234, 0.04872511, 0.04614759, 0.0450407, 
    0.04361912, 0.04123917, 0.03929344, 0.03723221, 0.03479517, 0.03344643, 
    0.03222003, 0.03048799, 0.02899776, 0.02858825, 0.02806287, 0.02674763, 
    0.02585599, 0.02564203, 0.02574769, 0.02595549, 0.02571911, 0.02588855, 
    0.0250362, 0.02480355, 0.02508421, 0.02580362, 0.02681372, 0.02832215, 
    0.02931329, 0.03117938, 0.03322739, 0.03502941, 0.03654204, 0.03833428, 
    0.04051844, 0.04289852, 0.04505702, 0.04783924, 0.04986884, 0.0514797, 
    0.05299488, 0.05324303, 0.05227294, 0.0512764, 0.04949561, 0.04653801, 
    0.04313298, 0.03967862, 0.03672488, 0.03422141, 0.03147369, 0.02854064, 
    0.02526513, 0.02038726, 0.01341081, 0.009903434, 0.004027471, 0.0106778, 
    0.01920674, 0.05279155, 0.084212, 0.06601435, 0.05526597, 0.05292657, 
    0.04991566, 0.04604028, 0.04476362, 0.04376495, 0.04778125, 0.04885961, 
    0.04905611, 0.04883939, 0.05003735, 0.0538695, 0.05548009, 0.06643351, 
    0.08635531, 0.09104959, 0.08267605, 0.06281079, 0.04780118, 0.03974854, 
    0.0359909, 0.03284637, 0.0298658, 0.02775005, 0.02594682, 0.02455248, 
    0.0231775, 0.02239563, 0.02192679, 0.0217841, 0.02246992, 0.02280786, 
    0.02281955, 0.02349836, 0.02448757, 0.02610885, 0.02723401, 0.02828491, 
    0.02837634, 0.02875873, 0.03014969, 0.03236313, 0.03424551, 0.03596223, 
    0.03755056, 0.03941764, 0.040874, 0.04205302, 0.04234504, 0.04227832,
  0.04216661, 0.04020581, 0.03634609, 0.03182127, 0.02732747, 0.0229917, 
    0.01934733, 0.017107, 0.0161265, 0.01768064, 0.01566215, 0.01695147, 
    0.02144136, 0.02663409, 0.02784944, 0.02705043, 0.02808168, 0.02936803, 
    0.03048057, 0.03028696, 0.03055059, 0.03283902, 0.04096051, 0.05458817, 
    0.06584486, 0.06504653, 0.06183807, 0.04370331, 0.03235639, 0.02688975, 
    0.0230163, 0.02090239, 0.01942638, 0.01740691, 0.02009662, 0.03582814, 
    0.0506283, 0.09828635, 0.1151878, 0.05281657, 0.03717807, 0.03063773, 
    0.02825263, 0.02520582, 0.02957463, 0.0313153, 0.0318794, 0.03102575, 
    0.03185653, 0.03233961, 0.0323418, 0.03254761, 0.0341011, 0.03453701, 
    0.03399521, 0.03360668, 0.03460462, 0.03474669, 0.03483608, 0.03563214, 
    0.03505635, 0.03358199, 0.03321274, 0.03353332, 0.03421601, 0.03522299, 
    0.03587227, 0.03670598, 0.03818079, 0.03901846, 0.03974996, 0.04033501, 
    0.04132147, 0.04186361, 0.04261445, 0.04228172, 0.04143681, 0.04128836, 
    0.04199928, 0.04192444, 0.04146271, 0.04056047, 0.03931369, 0.0370624, 
    0.03446442, 0.03021439, 0.02495596, 0.01985374, 0.01598517, 0.01346284, 
    0.01247358, 0.01201194, 0.01284966, 0.01485333, 0.01580286, 0.01588091, 
    0.01672291, 0.01845331, 0.02087268, 0.02303533, 0.02520124, 0.02743479, 
    0.02900012, 0.030958, 0.03291653, 0.03300916, 0.03352081, 0.03307303, 
    0.03389448, 0.03436151, 0.03375865, 0.03262619, 0.03412317, 0.03651707, 
    0.03697648, 0.04378682, 0.05231166, 0.05018347, 0.04989341, 0.04425039, 
    0.0407141, 0.03719612, 0.03740126, 0.03840427, 0.0387141, 0.03797661, 
    0.03812515, 0.03976738, 0.0417299, 0.04190538, 0.04121084, 0.04211729, 
    0.04954287, 0.05290252, 0.05402748, 0.05513133, 0.0568944, 0.06019673, 
    0.06400271, 0.06587535, 0.06907455, 0.07305945, 0.07659078, 0.0771058, 
    0.07442943, 0.07276041, 0.07393634, 0.07518421, 0.0744395, 0.07300154, 
    0.07265868, 0.07341288, 0.07495794, 0.0735574, 0.07201894, 0.07079641, 
    0.06934506, 0.06782095, 0.06654724, 0.06555276, 0.06357843, 0.06296413, 
    0.06151862, 0.06026734, 0.06018997, 0.05891904, 0.05618813, 0.05579792, 
    0.05619105, 0.05575038, 0.05613059, 0.05591631, 0.05464568, 0.05134986, 
    0.04765517, 0.04489631, 0.04267754, 0.04053786, 0.03958898, 0.03990055, 
    0.038598, 0.03651334, 0.03429711, 0.03173801, 0.03009669, 0.02962176, 
    0.02862615, 0.02730895, 0.02638271, 0.02585349, 0.02468498, 0.02340001, 
    0.02312918, 0.02351848, 0.02419589, 0.02412321, 0.02351749, 0.02342073, 
    0.02355894, 0.02395938, 0.0243246, 0.02574962, 0.02715274, 0.02853757, 
    0.02961561, 0.03143691, 0.03376797, 0.03655721, 0.0388452, 0.04136422, 
    0.04348985, 0.04587892, 0.04875981, 0.05181467, 0.05426519, 0.05599007, 
    0.05714191, 0.0565359, 0.0553298, 0.05424415, 0.05223805, 0.04870724, 
    0.04529761, 0.04200178, 0.03902503, 0.03630628, 0.03263576, 0.02919688, 
    0.02524982, 0.01948361, 0.01090508, 0.01037967, 0.006787633, 0.01365321, 
    0.01749688, 0.04187559, 0.07892479, 0.06413097, 0.05459251, 0.05132018, 
    0.0474399, 0.04418001, 0.04339489, 0.04346685, 0.04530154, 0.04897012, 
    0.05034319, 0.04889548, 0.0489109, 0.04998813, 0.0554516, 0.06299075, 
    0.07870051, 0.08674092, 0.09110413, 0.07751197, 0.04782173, 0.03700595, 
    0.03244402, 0.02901903, 0.02618299, 0.02422575, 0.02272582, 0.02207524, 
    0.02124491, 0.02036124, 0.01968801, 0.02002906, 0.02086822, 0.02139003, 
    0.02179507, 0.02316024, 0.02467102, 0.02580122, 0.02652885, 0.02813269, 
    0.02888783, 0.03046819, 0.03220164, 0.03453689, 0.03628084, 0.03794455, 
    0.03969404, 0.04180532, 0.04308701, 0.04379598, 0.04349544, 0.04313323,
  0.04299619, 0.04046569, 0.03595032, 0.03155327, 0.02679152, 0.02270715, 
    0.01933294, 0.01702348, 0.01592638, 0.01462514, 0.01499515, 0.01800529, 
    0.02391857, 0.02780724, 0.0280081, 0.02770762, 0.02892473, 0.03083539, 
    0.03224066, 0.03025328, 0.03175506, 0.03393847, 0.03679339, 0.04555036, 
    0.05576823, 0.06340671, 0.06522184, 0.04982583, 0.03674006, 0.02852702, 
    0.02401878, 0.0211426, 0.01974157, 0.01770893, 0.02133846, 0.04426489, 
    0.06670037, 0.08425589, 0.1368112, 0.06463555, 0.04347079, 0.03313056, 
    0.0297527, 0.02881162, 0.02934136, 0.03104293, 0.03126782, 0.03087722, 
    0.0312757, 0.03138644, 0.03160488, 0.03190243, 0.03329065, 0.03408207, 
    0.03420864, 0.034328, 0.03452777, 0.0352686, 0.03575455, 0.03614166, 
    0.0350758, 0.0340414, 0.03444733, 0.03496031, 0.03517469, 0.03575435, 
    0.03630284, 0.03679458, 0.03801546, 0.03997122, 0.04005531, 0.03955656, 
    0.03990714, 0.04070783, 0.04157228, 0.04199039, 0.04196958, 0.04209173, 
    0.04269627, 0.04271311, 0.04182439, 0.04089555, 0.03935581, 0.03673515, 
    0.03402108, 0.03043997, 0.02571412, 0.02095897, 0.01768775, 0.01548755, 
    0.01433755, 0.01322557, 0.01180003, 0.01195003, 0.0134536, 0.01335678, 
    0.01476588, 0.01686249, 0.01963797, 0.02286626, 0.02629939, 0.02852443, 
    0.03012799, 0.03129534, 0.03311356, 0.0337152, 0.03314454, 0.03260394, 
    0.03283203, 0.03339878, 0.03335463, 0.03382769, 0.03553708, 0.03861059, 
    0.04028288, 0.0484623, 0.06068283, 0.05440753, 0.04446974, 0.04207205, 
    0.03800037, 0.03533138, 0.03600015, 0.03705501, 0.03780264, 0.03780405, 
    0.0388079, 0.04088144, 0.04278272, 0.04394069, 0.04544021, 0.04647521, 
    0.05076092, 0.05320083, 0.05289754, 0.0540847, 0.05671911, 0.06031314, 
    0.06369644, 0.06555177, 0.06915063, 0.07320867, 0.07561161, 0.07384203, 
    0.07060695, 0.07077528, 0.07261758, 0.072463, 0.07096796, 0.06933644, 
    0.06911149, 0.07011735, 0.0705747, 0.06954268, 0.06800662, 0.065808, 
    0.0642744, 0.06354409, 0.06399719, 0.06471869, 0.06281945, 0.06103101, 
    0.05977151, 0.05811082, 0.05750418, 0.05550166, 0.05353658, 0.05358909, 
    0.05402653, 0.05343645, 0.05155057, 0.04915756, 0.04655074, 0.04299505, 
    0.03928615, 0.03699965, 0.03587903, 0.03529871, 0.03510327, 0.03534982, 
    0.03413093, 0.03262589, 0.03027541, 0.02791906, 0.02675869, 0.02627483, 
    0.02597089, 0.02483772, 0.02369543, 0.02290456, 0.02206892, 0.02159348, 
    0.02154334, 0.02204191, 0.02255537, 0.02225446, 0.02217358, 0.02237245, 
    0.02287953, 0.02328394, 0.02412557, 0.02551493, 0.02696547, 0.02825712, 
    0.02955289, 0.03224272, 0.03521082, 0.03824577, 0.04106702, 0.04372681, 
    0.04621296, 0.04895772, 0.05228245, 0.05556944, 0.05774397, 0.05956873, 
    0.06062847, 0.05994581, 0.05815795, 0.05655166, 0.0536874, 0.05024719, 
    0.04709954, 0.04362834, 0.04046646, 0.0368569, 0.0331995, 0.03006218, 
    0.0242169, 0.01611128, 0.007925609, 0.009655903, 0.01388041, 0.0181629, 
    0.02290377, 0.04681217, 0.07788865, 0.06623655, 0.05281707, 0.04955507, 
    0.04647796, 0.04345243, 0.04206785, 0.04379883, 0.04588091, 0.04952642, 
    0.05181029, 0.04952125, 0.04690299, 0.04694742, 0.05807507, 0.06276032, 
    0.06594647, 0.07605503, 0.07775799, 0.06916562, 0.0461049, 0.0348544, 
    0.02914186, 0.02600485, 0.02348928, 0.02157265, 0.02071496, 0.02038358, 
    0.01968517, 0.01889827, 0.0188628, 0.01963305, 0.02031436, 0.02070723, 
    0.02177501, 0.02329386, 0.02446716, 0.02521872, 0.02638271, 0.02822183, 
    0.02999086, 0.03245983, 0.0344477, 0.03658201, 0.03829025, 0.04032321, 
    0.04232977, 0.04476046, 0.04584832, 0.04566597, 0.04481791, 0.04442688,
  0.0438526, 0.04017429, 0.03556862, 0.03105348, 0.02627701, 0.02218474, 
    0.0187603, 0.01588864, 0.01372137, 0.0125213, 0.01670001, 0.0215173, 
    0.02612065, 0.02730876, 0.02714253, 0.02868257, 0.03068309, 0.03289949, 
    0.03381572, 0.03279519, 0.03288619, 0.03745565, 0.04369016, 0.04413052, 
    0.04689696, 0.05900144, 0.06201784, 0.05171086, 0.04548139, 0.03370902, 
    0.02688744, 0.02266541, 0.02126013, 0.02021242, 0.02622248, 0.05357946, 
    0.07544371, 0.08383951, 0.1197556, 0.08723862, 0.05121953, 0.03608569, 
    0.03188279, 0.03190073, 0.03228259, 0.03180504, 0.03153743, 0.03100622, 
    0.03103903, 0.03118718, 0.03140141, 0.03246156, 0.03362906, 0.03398958, 
    0.03391154, 0.03489592, 0.03539196, 0.03598131, 0.03630692, 0.0356042, 
    0.03473719, 0.03485343, 0.03530362, 0.0352762, 0.03514651, 0.03524602, 
    0.03594837, 0.03629936, 0.03736674, 0.03918044, 0.03879015, 0.03874275, 
    0.03934421, 0.04048342, 0.04159568, 0.04280999, 0.04344952, 0.04368071, 
    0.04382924, 0.04324847, 0.04195044, 0.04012496, 0.03828613, 0.03592164, 
    0.03381414, 0.03052397, 0.02626755, 0.02213668, 0.01893648, 0.01653146, 
    0.0148859, 0.01343015, 0.01196604, 0.0113471, 0.01104931, 0.01150517, 
    0.01329471, 0.01564633, 0.01902914, 0.02389062, 0.02867076, 0.03096062, 
    0.03197128, 0.03168355, 0.03327134, 0.03443199, 0.03339319, 0.03223993, 
    0.0326294, 0.03258887, 0.03322108, 0.03401827, 0.03624274, 0.04198333, 
    0.04605861, 0.04973472, 0.07270985, 0.0555191, 0.04557023, 0.04056946, 
    0.03732274, 0.03661832, 0.03799067, 0.03949851, 0.04104676, 0.04232741, 
    0.04306458, 0.04406103, 0.04452318, 0.04539291, 0.0465259, 0.04850939, 
    0.05031109, 0.05143594, 0.05233437, 0.05464555, 0.05731357, 0.05986365, 
    0.06177469, 0.06383494, 0.06803336, 0.0674677, 0.07242548, 0.07321045, 
    0.06874581, 0.0688331, 0.06986261, 0.06879231, 0.06658968, 0.06502623, 
    0.06455863, 0.06552148, 0.06593485, 0.06695178, 0.06563552, 0.06378717, 
    0.06199325, 0.06090527, 0.06186051, 0.06268932, 0.06106901, 0.05765215, 
    0.05443807, 0.05331505, 0.05271551, 0.05032908, 0.04874403, 0.04921388, 
    0.05053068, 0.04965336, 0.04641106, 0.04205368, 0.03881139, 0.03566756, 
    0.03265436, 0.03076101, 0.031022, 0.03078975, 0.03078995, 0.0311792, 
    0.03053983, 0.02904621, 0.02653274, 0.02467087, 0.02374399, 0.02308293, 
    0.02277796, 0.02197107, 0.02124229, 0.02119966, 0.02057861, 0.02027214, 
    0.02044329, 0.02047615, 0.02059363, 0.02101628, 0.02159561, 0.02211644, 
    0.02228736, 0.02306141, 0.02414324, 0.02511211, 0.02663281, 0.02879246, 
    0.03064672, 0.03360442, 0.03668704, 0.03987625, 0.04281673, 0.04543984, 
    0.04815377, 0.05169893, 0.05551193, 0.05911129, 0.0609998, 0.06232661, 
    0.06303822, 0.06217998, 0.05980429, 0.05717183, 0.05410192, 0.05076969, 
    0.04753764, 0.04396423, 0.04056324, 0.03678329, 0.03371868, 0.02756237, 
    0.01852737, 0.009719438, 0.01272843, 0.01634443, 0.02528441, 0.02523177, 
    0.03237272, 0.06694693, 0.08603094, 0.06301083, 0.05191104, 0.04695589, 
    0.04472154, 0.04215419, 0.04186198, 0.04461322, 0.04650064, 0.05006362, 
    0.05260324, 0.04914908, 0.04710566, 0.04676029, 0.05392382, 0.05613862, 
    0.05574117, 0.07567748, 0.07538401, 0.06690407, 0.04422141, 0.03237831, 
    0.02595668, 0.02310805, 0.02102509, 0.01957367, 0.01941929, 0.01905757, 
    0.01835135, 0.01824097, 0.01884322, 0.01924951, 0.01988084, 0.02066882, 
    0.02209419, 0.02340509, 0.02430952, 0.02514465, 0.027049, 0.02915192, 
    0.03173371, 0.03455109, 0.03661806, 0.03863632, 0.04102369, 0.043362, 
    0.04538382, 0.04724773, 0.04783748, 0.04755057, 0.04677325, 0.04585015,
  0.04372694, 0.03944189, 0.03492884, 0.03046212, 0.02570527, 0.02138029, 
    0.01826363, 0.01476855, 0.01170743, 0.01363416, 0.01966455, 0.02647003, 
    0.02895427, 0.02845836, 0.02920924, 0.03077395, 0.03283221, 0.03471357, 
    0.03495165, 0.03504256, 0.03410416, 0.04064623, 0.0456502, 0.04378717, 
    0.04191379, 0.04582771, 0.04858925, 0.05034202, 0.05349689, 0.04629545, 
    0.03443468, 0.02768509, 0.02559459, 0.02378613, 0.02991574, 0.05309578, 
    0.07468498, 0.07227303, 0.09987955, 0.1014256, 0.05836045, 0.04126669, 
    0.03436972, 0.03362927, 0.03380646, 0.03302662, 0.03260177, 0.03278142, 
    0.03214593, 0.03191883, 0.03175738, 0.03235656, 0.03368475, 0.03363681, 
    0.03339776, 0.03425755, 0.03571158, 0.03660661, 0.03669801, 0.03487508, 
    0.03479921, 0.03481994, 0.03473664, 0.03461182, 0.03498819, 0.03503728, 
    0.03604198, 0.03657696, 0.03720909, 0.03829285, 0.03829341, 0.03868871, 
    0.03934934, 0.04038218, 0.04102352, 0.04254564, 0.04379037, 0.04392882, 
    0.04354156, 0.04224923, 0.04063745, 0.03946017, 0.03742046, 0.03530335, 
    0.03348726, 0.03053409, 0.02698481, 0.02349564, 0.02019383, 0.01718689, 
    0.01467426, 0.0133032, 0.01261034, 0.01157182, 0.01048997, 0.01066793, 
    0.01210298, 0.0153386, 0.01909552, 0.02570804, 0.03295988, 0.03424773, 
    0.03399948, 0.03093428, 0.03302766, 0.03527831, 0.03505846, 0.03461272, 
    0.03565494, 0.03412964, 0.03323594, 0.0326906, 0.03535325, 0.04656459, 
    0.05249583, 0.05022857, 0.0790225, 0.05332664, 0.04408431, 0.03947807, 
    0.03830298, 0.03961573, 0.04140298, 0.04283235, 0.04552295, 0.04753767, 
    0.04636366, 0.04541756, 0.04483952, 0.04549576, 0.04708743, 0.04854121, 
    0.05076983, 0.05247863, 0.05450677, 0.05776904, 0.05924198, 0.06068392, 
    0.06078382, 0.06202624, 0.06426524, 0.05846934, 0.06632078, 0.07113531, 
    0.06815088, 0.06682927, 0.06523218, 0.06452254, 0.064033, 0.06221639, 
    0.06115323, 0.06095116, 0.06071622, 0.06181515, 0.06177664, 0.06084292, 
    0.05918142, 0.05761976, 0.05745764, 0.05658662, 0.05622137, 0.05400445, 
    0.05138407, 0.0489617, 0.04758181, 0.04621971, 0.04530085, 0.04473442, 
    0.0461167, 0.04512714, 0.04244014, 0.03756046, 0.03432648, 0.03082876, 
    0.02842413, 0.02734056, 0.02733945, 0.02735904, 0.02762375, 0.0271511, 
    0.02736499, 0.0264716, 0.02404844, 0.02245202, 0.0216526, 0.02094864, 
    0.02011472, 0.01946782, 0.01933558, 0.02011568, 0.02008649, 0.01940355, 
    0.01904011, 0.01900782, 0.01961632, 0.02065708, 0.02112338, 0.02122797, 
    0.02157535, 0.02233048, 0.02370135, 0.0250081, 0.02670619, 0.0287108, 
    0.03147346, 0.03448039, 0.03743424, 0.04092763, 0.0441213, 0.04685247, 
    0.04992304, 0.05396781, 0.05797727, 0.06104624, 0.06288786, 0.06419312, 
    0.06454305, 0.06266545, 0.05995233, 0.05703053, 0.05383236, 0.05042915, 
    0.04671544, 0.04254725, 0.03885854, 0.03489786, 0.02855926, 0.02265458, 
    0.02089814, 0.0159143, 0.01803419, 0.02369787, 0.02925832, 0.04431651, 
    0.07934052, 0.1055891, 0.101804, 0.06580637, 0.0504301, 0.04626942, 
    0.04312824, 0.04187994, 0.04277578, 0.04465055, 0.04679776, 0.04833857, 
    0.05014431, 0.05032055, 0.04690008, 0.04791697, 0.05305535, 0.05209569, 
    0.04667891, 0.06235106, 0.07125892, 0.06803547, 0.04695853, 0.03033884, 
    0.02324784, 0.02082735, 0.01957036, 0.01880782, 0.01847765, 0.0178809, 
    0.01765883, 0.0182228, 0.01876299, 0.01912465, 0.01998798, 0.02111909, 
    0.0224523, 0.02353086, 0.02456865, 0.02624884, 0.02841286, 0.03067891, 
    0.03363465, 0.03623569, 0.03851372, 0.0409611, 0.0436741, 0.0457488, 
    0.04741954, 0.04834727, 0.04884798, 0.04811301, 0.04766045, 0.04643441,
  0.0423949, 0.03856331, 0.03421891, 0.02990185, 0.02512141, 0.02119477, 
    0.01821075, 0.01475818, 0.01219589, 0.01574056, 0.02226985, 0.0292813, 
    0.03261842, 0.03055008, 0.03156164, 0.03353705, 0.03505921, 0.03651413, 
    0.03606935, 0.03779737, 0.03660414, 0.03966139, 0.04450943, 0.04259096, 
    0.04047976, 0.04355882, 0.04611431, 0.05309533, 0.06590915, 0.06194624, 
    0.04852507, 0.03728782, 0.03035218, 0.02720808, 0.03062593, 0.04420776, 
    0.06084031, 0.06483798, 0.0694019, 0.08895489, 0.06210097, 0.04633205, 
    0.03663347, 0.03391965, 0.03323886, 0.03338155, 0.03364369, 0.03397766, 
    0.03330067, 0.03268604, 0.03305941, 0.03327546, 0.03309934, 0.03248401, 
    0.03261665, 0.03433501, 0.03660735, 0.03746996, 0.03669937, 0.03536653, 
    0.0354795, 0.03549141, 0.0354714, 0.035191, 0.03548574, 0.03570432, 
    0.03648338, 0.03710609, 0.03748785, 0.03790559, 0.03845489, 0.03884868, 
    0.03987444, 0.04034669, 0.04074914, 0.04216696, 0.04330424, 0.04329067, 
    0.04232334, 0.04067639, 0.03919495, 0.03772219, 0.03587474, 0.03386695, 
    0.03279931, 0.03076672, 0.02781128, 0.02490882, 0.0216952, 0.01851279, 
    0.01614048, 0.01516884, 0.01387933, 0.01245862, 0.01110858, 0.01084151, 
    0.01240851, 0.01519109, 0.01900224, 0.02695726, 0.03597397, 0.03670685, 
    0.03211699, 0.02908001, 0.03216954, 0.03594033, 0.03709366, 0.03600565, 
    0.03561295, 0.03321263, 0.03240282, 0.03353531, 0.03728151, 0.04927275, 
    0.05366713, 0.04559201, 0.06007801, 0.04903309, 0.0442246, 0.04107937, 
    0.0407376, 0.04300776, 0.04483647, 0.04559296, 0.04831963, 0.05074701, 
    0.04781984, 0.04681242, 0.04694786, 0.04744564, 0.04901708, 0.05044056, 
    0.05246776, 0.05446525, 0.05676081, 0.05963834, 0.06136656, 0.06207142, 
    0.06107199, 0.06090267, 0.06088246, 0.05812981, 0.05698504, 0.06354034, 
    0.06587187, 0.06499133, 0.06373025, 0.062833, 0.06298885, 0.06071918, 
    0.05913566, 0.05804224, 0.05588056, 0.05534394, 0.05514839, 0.05502402, 
    0.05529966, 0.05416299, 0.05282305, 0.05124819, 0.05065544, 0.04867977, 
    0.04720569, 0.04503676, 0.04323735, 0.04327734, 0.04232058, 0.042113, 
    0.04103119, 0.04078171, 0.03788549, 0.03411185, 0.03160734, 0.02862064, 
    0.02601809, 0.02422785, 0.02382262, 0.0246033, 0.02498772, 0.02461247, 
    0.02525831, 0.02485637, 0.0223107, 0.02039269, 0.01942692, 0.01871275, 
    0.018215, 0.01777463, 0.01799039, 0.01875514, 0.01898772, 0.01802482, 
    0.01774975, 0.01829854, 0.01883074, 0.01947946, 0.01956977, 0.01948165, 
    0.02032898, 0.02197524, 0.02326285, 0.02480912, 0.02656201, 0.02850087, 
    0.03133273, 0.03457382, 0.03757948, 0.04120052, 0.0448335, 0.04825151, 
    0.05189013, 0.05516703, 0.05862549, 0.06150848, 0.06349091, 0.06445613, 
    0.06427598, 0.06185449, 0.05898437, 0.05614277, 0.05233178, 0.04827186, 
    0.04420245, 0.04016254, 0.03642736, 0.03091875, 0.02557761, 0.02291697, 
    0.0181032, 0.02232335, 0.02369202, 0.02659, 0.05140363, 0.1065519, 
    0.1462363, 0.1086347, 0.07796828, 0.05558821, 0.0471767, 0.04633998, 
    0.04575913, 0.04572587, 0.04505551, 0.04466271, 0.04479125, 0.04540203, 
    0.05014691, 0.05030254, 0.04741082, 0.0493385, 0.0511089, 0.05098052, 
    0.044441, 0.04888824, 0.06196655, 0.06941041, 0.05146205, 0.02938227, 
    0.02149954, 0.01982455, 0.01924172, 0.018562, 0.01786986, 0.01694527, 
    0.01728759, 0.01818483, 0.01865406, 0.0195828, 0.02073389, 0.02187862, 
    0.02300319, 0.02413843, 0.02553338, 0.02767143, 0.03031901, 0.03258086, 
    0.03491087, 0.0374235, 0.04051651, 0.0431995, 0.04550757, 0.04694874, 
    0.04817284, 0.04866418, 0.0486232, 0.04784316, 0.04718381, 0.04563356,
  0.04050653, 0.03661808, 0.03316415, 0.02921615, 0.02476963, 0.02154741, 
    0.01891518, 0.01659021, 0.01520508, 0.01977461, 0.02581844, 0.03088743, 
    0.03596399, 0.03499757, 0.03575072, 0.03806856, 0.03887907, 0.0394092, 
    0.03965051, 0.03959093, 0.0409591, 0.04057135, 0.04416884, 0.04835761, 
    0.04388713, 0.04853316, 0.05509684, 0.06448945, 0.06235783, 0.06240244, 
    0.05474456, 0.04537286, 0.03483298, 0.02928142, 0.0281132, 0.03136106, 
    0.03994293, 0.05551067, 0.06290723, 0.09365547, 0.06765097, 0.04991401, 
    0.03841304, 0.0343981, 0.03281315, 0.03329922, 0.0349794, 0.03582134, 
    0.0354066, 0.03339516, 0.03343681, 0.03416229, 0.03317022, 0.0325169, 
    0.03304029, 0.03420899, 0.03656944, 0.0376826, 0.03668908, 0.03525547, 
    0.03458036, 0.03532722, 0.03623234, 0.03653434, 0.03731915, 0.03733536, 
    0.03688402, 0.03703085, 0.03723086, 0.0375601, 0.03814457, 0.03759909, 
    0.03851705, 0.03922637, 0.03981932, 0.0413799, 0.04289924, 0.04350807, 
    0.04255586, 0.04058793, 0.03868502, 0.0368694, 0.03523763, 0.03404868, 
    0.0326296, 0.02974375, 0.02729351, 0.02461172, 0.02209649, 0.01977246, 
    0.01792642, 0.01779787, 0.01573359, 0.01407812, 0.01233706, 0.01181114, 
    0.01303789, 0.01496265, 0.01741374, 0.02465165, 0.03261919, 0.03150361, 
    0.02784272, 0.02657806, 0.03142634, 0.03741539, 0.0382749, 0.03331175, 
    0.03098175, 0.0300375, 0.03158044, 0.03563758, 0.04045684, 0.0491795, 
    0.04959489, 0.04166645, 0.04517756, 0.04602648, 0.04331268, 0.04169086, 
    0.04209011, 0.04466268, 0.04681282, 0.04818467, 0.05040513, 0.05300961, 
    0.05088897, 0.05051056, 0.05098573, 0.05030406, 0.05058, 0.05276914, 
    0.05313672, 0.05511943, 0.05802134, 0.06004245, 0.06220571, 0.06289529, 
    0.06152394, 0.06015876, 0.05906887, 0.05949437, 0.06082168, 0.06044924, 
    0.05920873, 0.061891, 0.06260938, 0.059829, 0.0582189, 0.05691197, 
    0.05689246, 0.05510455, 0.05252872, 0.05113339, 0.05092624, 0.05087198, 
    0.05062775, 0.04853333, 0.0464734, 0.04608842, 0.04572261, 0.04279872, 
    0.04071469, 0.03889536, 0.03866828, 0.03941374, 0.03835178, 0.03816426, 
    0.03702658, 0.03750522, 0.03351784, 0.03054725, 0.02929246, 0.02646149, 
    0.02404354, 0.0225214, 0.02208837, 0.02244057, 0.02317571, 0.02322556, 
    0.02365432, 0.02319926, 0.02097494, 0.01888145, 0.01757783, 0.01657392, 
    0.0161033, 0.01603166, 0.01645806, 0.01689385, 0.01717219, 0.01708503, 
    0.01731521, 0.01768837, 0.01786532, 0.01818875, 0.01839059, 0.01839181, 
    0.01933372, 0.02065714, 0.02206651, 0.02364392, 0.02560746, 0.02788349, 
    0.03073349, 0.03400457, 0.03715068, 0.04063113, 0.04416993, 0.0478645, 
    0.05148387, 0.05429765, 0.05738654, 0.06007865, 0.06193878, 0.06269704, 
    0.06238955, 0.06051991, 0.05724955, 0.05374532, 0.04969157, 0.04533629, 
    0.0410517, 0.03700485, 0.032291, 0.02405378, 0.01692557, 0.01113079, 
    0.01447757, 0.02740481, 0.03856573, 0.04782503, 0.08921872, 0.1605405, 
    0.1226006, 0.07535321, 0.06340627, 0.05053923, 0.04452368, 0.04575381, 
    0.04654424, 0.0479566, 0.04794954, 0.04451418, 0.0425236, 0.04369676, 
    0.04942588, 0.05159236, 0.0505666, 0.04764144, 0.04594873, 0.04605681, 
    0.04634189, 0.04310733, 0.05476864, 0.07279998, 0.05451851, 0.02832363, 
    0.02090216, 0.01920757, 0.01818561, 0.01753137, 0.01695056, 0.01636301, 
    0.01702121, 0.01774183, 0.01830944, 0.0193414, 0.0204946, 0.02169838, 
    0.02322596, 0.02488628, 0.02609788, 0.02836271, 0.03094267, 0.03361933, 
    0.03615672, 0.0389691, 0.04183476, 0.04397804, 0.04562122, 0.04678354, 
    0.04787558, 0.04877107, 0.04871219, 0.04785758, 0.04601702, 0.04334622,
  0.03912099, 0.03560761, 0.03192582, 0.02881582, 0.02538509, 0.02265582, 
    0.02051756, 0.01924281, 0.01917386, 0.025306, 0.02911218, 0.03517016, 
    0.04021771, 0.04017081, 0.04063577, 0.04296523, 0.04158752, 0.04349092, 
    0.04564485, 0.0445949, 0.04644999, 0.04743167, 0.04770497, 0.05426038, 
    0.05146442, 0.05102421, 0.0474655, 0.0550837, 0.05296158, 0.05303105, 
    0.04821289, 0.0425736, 0.03551565, 0.02927175, 0.02637043, 0.02565384, 
    0.0296233, 0.0491663, 0.06395064, 0.09607846, 0.06601256, 0.05038868, 
    0.03966537, 0.03547928, 0.03433359, 0.03457078, 0.03554283, 0.03501182, 
    0.03472545, 0.0333191, 0.03319709, 0.03334275, 0.03276109, 0.03249565, 
    0.0329184, 0.03301679, 0.03471864, 0.03651986, 0.03630247, 0.03547251, 
    0.03395424, 0.03440218, 0.03571664, 0.03656793, 0.03826575, 0.03862574, 
    0.03735876, 0.03677277, 0.03674496, 0.03728814, 0.03828515, 0.0366209, 
    0.03598523, 0.03705488, 0.03828762, 0.04012987, 0.04227782, 0.04322559, 
    0.04198967, 0.03969487, 0.03681069, 0.03449487, 0.03395031, 0.03331894, 
    0.03133061, 0.02886097, 0.02614449, 0.02305413, 0.02078336, 0.01958788, 
    0.01900994, 0.01944815, 0.01700542, 0.01530346, 0.01416587, 0.01419279, 
    0.01474376, 0.01465048, 0.01520631, 0.01989563, 0.02434973, 0.02394375, 
    0.02391214, 0.02583561, 0.03421036, 0.04050468, 0.03850719, 0.03142729, 
    0.02931735, 0.02921637, 0.03027405, 0.03311987, 0.03835684, 0.04485234, 
    0.04105033, 0.03765632, 0.04071658, 0.0406828, 0.03988202, 0.03950992, 
    0.04164362, 0.04414833, 0.04663981, 0.0488672, 0.05201446, 0.05527632, 
    0.05450232, 0.0555859, 0.05635344, 0.05489212, 0.0539741, 0.05550429, 
    0.0546939, 0.05721994, 0.05973494, 0.0612287, 0.06290676, 0.06357452, 
    0.06195489, 0.06020622, 0.06082327, 0.06027309, 0.05941769, 0.05839914, 
    0.05725694, 0.05719089, 0.05808048, 0.05619975, 0.05499083, 0.05349671, 
    0.05319118, 0.05066816, 0.04819098, 0.04709313, 0.04631614, 0.045531, 
    0.04355615, 0.04227877, 0.04112504, 0.04159252, 0.04138544, 0.03870272, 
    0.03580738, 0.03402898, 0.0342709, 0.03349264, 0.03293268, 0.03343574, 
    0.03263597, 0.03381223, 0.02964286, 0.02657222, 0.02568323, 0.02344706, 
    0.02255517, 0.02156384, 0.02051706, 0.0209663, 0.02205626, 0.02181734, 
    0.02166425, 0.02104607, 0.01963766, 0.01779085, 0.01645398, 0.01530559, 
    0.01488408, 0.01502836, 0.01554226, 0.01589447, 0.0162187, 0.01668832, 
    0.01686288, 0.01675743, 0.01708334, 0.01734545, 0.01750509, 0.01770705, 
    0.0182754, 0.01892399, 0.02035211, 0.02238189, 0.02449338, 0.02655024, 
    0.02963885, 0.03266433, 0.03601581, 0.03918953, 0.04198304, 0.04517559, 
    0.04840641, 0.05104105, 0.05418834, 0.05698632, 0.05845216, 0.05882981, 
    0.05833581, 0.05585507, 0.05322711, 0.05000649, 0.04605918, 0.0413142, 
    0.03730951, 0.03290447, 0.02513211, 0.01400885, 0.008650097, 0.009522755, 
    0.0218685, 0.05844008, 0.07474729, 0.1021618, 0.1461661, 0.1255836, 
    0.07980169, 0.06199441, 0.05293473, 0.04830332, 0.04699446, 0.04824562, 
    0.04696181, 0.04694797, 0.0465351, 0.04428196, 0.04288042, 0.04300329, 
    0.04746458, 0.0497242, 0.04857172, 0.04404603, 0.03979084, 0.04360088, 
    0.04921331, 0.04268617, 0.04582225, 0.06604269, 0.05727803, 0.02818624, 
    0.02022443, 0.01778742, 0.01682038, 0.0160357, 0.01574039, 0.01591924, 
    0.01680895, 0.01755313, 0.01820654, 0.01892653, 0.01986574, 0.0212488, 
    0.02305979, 0.02477727, 0.02661039, 0.02877467, 0.03138195, 0.03414688, 
    0.03676705, 0.03940123, 0.0412425, 0.0430281, 0.04481013, 0.04582468, 
    0.04721179, 0.04794342, 0.04791381, 0.04683756, 0.04488129, 0.04199958,
  0.03878085, 0.03493361, 0.03116632, 0.0283684, 0.0259635, 0.0238595, 
    0.02227317, 0.02141577, 0.02155914, 0.02793596, 0.03471843, 0.03922781, 
    0.04527927, 0.04413455, 0.04349053, 0.04483127, 0.0434676, 0.04538088, 
    0.04864746, 0.05023402, 0.05258783, 0.05248149, 0.04954701, 0.05474991, 
    0.06184628, 0.04645648, 0.03770771, 0.0417677, 0.05267588, 0.05132286, 
    0.04616842, 0.03943922, 0.03315541, 0.02877627, 0.02601336, 0.02472, 
    0.02849909, 0.04323968, 0.05290506, 0.04586206, 0.0489108, 0.04668191, 
    0.04011345, 0.0376744, 0.03688094, 0.0354933, 0.03446247, 0.0326597, 
    0.03244914, 0.0326809, 0.03296896, 0.03305622, 0.03268243, 0.03202596, 
    0.03132515, 0.03131866, 0.03263611, 0.03468373, 0.03570719, 0.03664817, 
    0.03540096, 0.03484475, 0.03509146, 0.0356786, 0.03690333, 0.03723141, 
    0.03644469, 0.03649453, 0.03674761, 0.03708041, 0.03804761, 0.03722012, 
    0.03575785, 0.03553746, 0.03652783, 0.03852418, 0.04050336, 0.04147696, 
    0.04011032, 0.03736756, 0.03453764, 0.03216493, 0.03207855, 0.03132529, 
    0.0298953, 0.02770014, 0.02499495, 0.02230939, 0.02022534, 0.01936158, 
    0.01868671, 0.01757617, 0.01577503, 0.01491465, 0.01445526, 0.01513542, 
    0.01626406, 0.01553464, 0.01471401, 0.01644974, 0.01785066, 0.01807032, 
    0.02033385, 0.02603271, 0.03799345, 0.04498928, 0.04140437, 0.03156256, 
    0.02880847, 0.02819709, 0.02825789, 0.02963898, 0.0346373, 0.03958044, 
    0.03658553, 0.03647683, 0.03774714, 0.035698, 0.0355549, 0.03649278, 
    0.03932595, 0.0420409, 0.04461055, 0.05004323, 0.05600702, 0.05896175, 
    0.05937911, 0.05982292, 0.05933544, 0.05918918, 0.05885854, 0.05810567, 
    0.0565308, 0.05794821, 0.05998507, 0.06274399, 0.06456778, 0.06519686, 
    0.06379513, 0.0628669, 0.06363327, 0.06046359, 0.05760123, 0.05573648, 
    0.05566748, 0.05521052, 0.05456784, 0.05468443, 0.05481305, 0.05230077, 
    0.05012597, 0.04678284, 0.04407182, 0.04163373, 0.0396789, 0.03694971, 
    0.03473293, 0.03531466, 0.0362841, 0.03733348, 0.03663687, 0.03325815, 
    0.03075614, 0.03032563, 0.02991121, 0.02961962, 0.02932382, 0.02932427, 
    0.02847865, 0.02688079, 0.02531276, 0.02307246, 0.02265938, 0.02068112, 
    0.01997314, 0.01975786, 0.01960775, 0.02021036, 0.02031359, 0.01943975, 
    0.01909351, 0.01893092, 0.01787219, 0.01661292, 0.01565404, 0.01488902, 
    0.01462238, 0.01491126, 0.01538988, 0.01558018, 0.01569333, 0.01615386, 
    0.0161876, 0.0161152, 0.01644004, 0.01639955, 0.01639025, 0.01677394, 
    0.01735643, 0.01799057, 0.01917037, 0.02089945, 0.02307057, 0.02511485, 
    0.02777869, 0.03042985, 0.03346079, 0.03647517, 0.0389626, 0.04230043, 
    0.04555852, 0.04806136, 0.05054454, 0.05228535, 0.05345275, 0.05361055, 
    0.05264177, 0.05074747, 0.04846155, 0.04499923, 0.04123559, 0.03768196, 
    0.03364699, 0.02733271, 0.01586093, 0.007166484, 0.01190725, 0.02169514, 
    0.07672745, 0.1117368, 0.1296194, 0.1650919, 0.1548588, 0.07555573, 
    0.06277859, 0.05269743, 0.04849338, 0.04791363, 0.04879242, 0.04950685, 
    0.04850142, 0.04938689, 0.04695013, 0.04470184, 0.04472522, 0.04477263, 
    0.04487383, 0.04407359, 0.04483669, 0.04307286, 0.04017419, 0.04216865, 
    0.04930147, 0.04297352, 0.04721652, 0.06110052, 0.05606444, 0.02775775, 
    0.01957101, 0.01622926, 0.01544013, 0.01482289, 0.01494272, 0.01566069, 
    0.0166517, 0.01725021, 0.01744118, 0.01815502, 0.01928981, 0.02069979, 
    0.02241441, 0.02446781, 0.02640421, 0.02820377, 0.03020827, 0.03244908, 
    0.03537826, 0.03790539, 0.03952328, 0.04127985, 0.04352053, 0.04458643, 
    0.04577079, 0.04671418, 0.04640473, 0.04563091, 0.04358928, 0.04155273,
  0.03755791, 0.03453217, 0.03110169, 0.02857629, 0.02655727, 0.02480066, 
    0.02324592, 0.02246073, 0.02306661, 0.02733148, 0.04047787, 0.04432981, 
    0.04661399, 0.04791588, 0.04515084, 0.04347184, 0.04337459, 0.04687808, 
    0.04986137, 0.05353642, 0.05402862, 0.0550168, 0.05192055, 0.04525053, 
    0.0587681, 0.05483134, 0.04128827, 0.04605203, 0.05021961, 0.04935754, 
    0.04427588, 0.03745947, 0.03265255, 0.02888366, 0.0250452, 0.02321386, 
    0.02525277, 0.0305248, 0.03428219, 0.03402434, 0.04200177, 0.04391901, 
    0.04099589, 0.03982061, 0.04032899, 0.03697019, 0.0348414, 0.03397675, 
    0.03421101, 0.03372591, 0.0335333, 0.03483243, 0.03535217, 0.03446578, 
    0.03266518, 0.03226313, 0.03295735, 0.03448261, 0.03508064, 0.03590327, 
    0.03605485, 0.03542838, 0.03454923, 0.03523528, 0.03606075, 0.03585393, 
    0.03560141, 0.03579247, 0.03636716, 0.03695549, 0.03724914, 0.03715829, 
    0.03597762, 0.0343926, 0.0339866, 0.03526365, 0.03632166, 0.03735054, 
    0.03692093, 0.03486785, 0.0327706, 0.03087467, 0.03029644, 0.02960366, 
    0.02902932, 0.0264547, 0.02333231, 0.02099488, 0.01944427, 0.0186229, 
    0.01759944, 0.01588944, 0.01491218, 0.01458966, 0.01430759, 0.01467675, 
    0.01578909, 0.01552078, 0.01528092, 0.01637919, 0.01667332, 0.01703017, 
    0.01914839, 0.0258155, 0.03726483, 0.03857512, 0.0343484, 0.02779124, 
    0.02659863, 0.02694428, 0.02531859, 0.02655356, 0.03085515, 0.03451673, 
    0.03449631, 0.03474632, 0.03388328, 0.03352865, 0.03471323, 0.03850687, 
    0.04030824, 0.04149914, 0.04405287, 0.05030148, 0.05927445, 0.06238917, 
    0.06425201, 0.06326766, 0.06091328, 0.06200593, 0.06291165, 0.06039861, 
    0.05807103, 0.05908972, 0.06071087, 0.06519275, 0.0682502, 0.06929122, 
    0.06851462, 0.06596784, 0.06447748, 0.05990601, 0.05635721, 0.05467459, 
    0.05530366, 0.05490793, 0.05379457, 0.05329983, 0.05276116, 0.0498955, 
    0.04721371, 0.04390439, 0.04075155, 0.03702822, 0.03444942, 0.03142879, 
    0.03040328, 0.03164926, 0.03251958, 0.03260054, 0.03098698, 0.02826064, 
    0.02691194, 0.02740375, 0.02772141, 0.02801431, 0.02763579, 0.02715388, 
    0.02521108, 0.0229317, 0.02115203, 0.0206257, 0.01970084, 0.01843995, 
    0.01822589, 0.01897147, 0.01972371, 0.02003251, 0.01916178, 0.01747431, 
    0.01655077, 0.01659509, 0.01592219, 0.01506782, 0.0145585, 0.01457911, 
    0.01456423, 0.0146723, 0.01468074, 0.01454196, 0.0145699, 0.01528181, 
    0.01559289, 0.01564625, 0.01588702, 0.01564512, 0.0156416, 0.01582589, 
    0.01630411, 0.01703884, 0.01813046, 0.01962958, 0.0215009, 0.02383166, 
    0.02601825, 0.02808663, 0.03065029, 0.03366201, 0.03645767, 0.03990391, 
    0.04321113, 0.04562029, 0.04700408, 0.04807216, 0.04850055, 0.04848348, 
    0.04758359, 0.04589523, 0.04335354, 0.04071581, 0.03759969, 0.0342448, 
    0.02984516, 0.02061823, 0.008921111, 0.009628393, 0.02479095, 0.06223937, 
    0.1306416, 0.1443544, 0.1314225, 0.1190315, 0.0785855, 0.06013626, 
    0.05305789, 0.04984933, 0.04884085, 0.04974245, 0.04948071, 0.04893238, 
    0.05226706, 0.05415189, 0.05053717, 0.04611492, 0.04724663, 0.04572117, 
    0.0415817, 0.03992937, 0.04272679, 0.04444754, 0.04178867, 0.04340576, 
    0.05103402, 0.04369699, 0.04330924, 0.05252602, 0.05086487, 0.03355493, 
    0.02028083, 0.01606001, 0.01473622, 0.01437518, 0.01459162, 0.01558172, 
    0.01650751, 0.01689865, 0.01712145, 0.01779589, 0.0186984, 0.01986994, 
    0.02147211, 0.02303925, 0.02476423, 0.02641311, 0.02800153, 0.03044235, 
    0.03311912, 0.0352614, 0.03717154, 0.03936204, 0.0413268, 0.04261477, 
    0.04380403, 0.04499237, 0.04507411, 0.04424183, 0.04254121, 0.04047656,
  0.0375273, 0.03478645, 0.0313192, 0.02889857, 0.02702646, 0.02528637, 
    0.02336341, 0.02293937, 0.02448793, 0.02580344, 0.04026657, 0.04393364, 
    0.04595832, 0.04875669, 0.04698424, 0.04140012, 0.04283667, 0.04994723, 
    0.05373645, 0.0541933, 0.05181693, 0.05206366, 0.05250445, 0.04660169, 
    0.04784034, 0.05639151, 0.04661103, 0.05231894, 0.05045853, 0.05265594, 
    0.04489746, 0.0382296, 0.03316589, 0.03006677, 0.02658789, 0.02380733, 
    0.02381619, 0.02513765, 0.02852767, 0.03414698, 0.03918673, 0.04227448, 
    0.03939676, 0.03840461, 0.03907568, 0.03673568, 0.03480998, 0.03470937, 
    0.03496395, 0.03445977, 0.03459429, 0.0354242, 0.03548143, 0.03505443, 
    0.03389635, 0.03372924, 0.03514265, 0.03582091, 0.03463382, 0.03460807, 
    0.03585596, 0.03542955, 0.03464552, 0.0354372, 0.03613609, 0.03601567, 
    0.03559125, 0.03514643, 0.03565881, 0.03581578, 0.036117, 0.0356904, 
    0.03419676, 0.03282375, 0.03240491, 0.03254771, 0.03283582, 0.03283292, 
    0.03349663, 0.0327368, 0.03150272, 0.0300147, 0.02837239, 0.02717944, 
    0.02622234, 0.02410895, 0.02167139, 0.01950659, 0.01790858, 0.01694287, 
    0.01563257, 0.01463163, 0.0140835, 0.01385517, 0.013848, 0.01410267, 
    0.01520819, 0.01565583, 0.01594574, 0.01696886, 0.01698174, 0.01806221, 
    0.01939, 0.02215276, 0.02517012, 0.02420475, 0.0227703, 0.02187122, 
    0.02389186, 0.0273647, 0.02477834, 0.02444545, 0.02579702, 0.02864379, 
    0.03226549, 0.03242822, 0.03203248, 0.03581398, 0.04074254, 0.04414979, 
    0.04447621, 0.04272175, 0.04468, 0.05171378, 0.05738278, 0.0613086, 
    0.06473036, 0.06519751, 0.06242186, 0.06219086, 0.06329142, 0.06313763, 
    0.06231892, 0.06349438, 0.06516349, 0.06847908, 0.06960304, 0.07051796, 
    0.06928223, 0.06433726, 0.06196488, 0.05848365, 0.0556428, 0.05411381, 
    0.0529337, 0.05258017, 0.05209548, 0.05055955, 0.04817487, 0.04609483, 
    0.04388502, 0.04027086, 0.03724275, 0.03352833, 0.03109461, 0.02898942, 
    0.0293651, 0.03010395, 0.0301163, 0.02945765, 0.02724379, 0.02619186, 
    0.02600022, 0.02574001, 0.02656102, 0.02649644, 0.02510114, 0.0239107, 
    0.02175576, 0.02010511, 0.01905269, 0.01857656, 0.01704, 0.01681199, 
    0.01741019, 0.01805185, 0.01882, 0.01905757, 0.01800277, 0.01602688, 
    0.01511192, 0.01545242, 0.01498704, 0.01455343, 0.0139479, 0.01390586, 
    0.01387007, 0.01375331, 0.0136371, 0.01358793, 0.01385676, 0.01483403, 
    0.01519065, 0.01515983, 0.01541116, 0.0153916, 0.01543604, 0.01535234, 
    0.01528917, 0.0158514, 0.01725403, 0.01854656, 0.02014624, 0.02247693, 
    0.02480256, 0.02652115, 0.02915661, 0.03218944, 0.03505009, 0.03799124, 
    0.0407143, 0.04243866, 0.04395159, 0.04444959, 0.04468349, 0.04484234, 
    0.04399522, 0.04240048, 0.04016038, 0.0377843, 0.03494764, 0.03170665, 
    0.02577673, 0.01450374, 0.007603481, 0.02004693, 0.05443425, 0.1163759, 
    0.1328436, 0.09967396, 0.08183423, 0.07126284, 0.06148378, 0.05119469, 
    0.04801753, 0.04837068, 0.04961465, 0.0521558, 0.05289544, 0.05410042, 
    0.05522531, 0.05451911, 0.0526971, 0.04891959, 0.04855297, 0.04582565, 
    0.04171047, 0.04103832, 0.04449187, 0.0467032, 0.04254233, 0.04390001, 
    0.04917857, 0.04068715, 0.03514274, 0.04392091, 0.04461459, 0.0407213, 
    0.02532224, 0.01814705, 0.01572924, 0.01479603, 0.01477379, 0.01565087, 
    0.01631418, 0.01684083, 0.01687329, 0.01737081, 0.01804993, 0.01905049, 
    0.02016493, 0.02119663, 0.02280483, 0.02445067, 0.02596925, 0.02827203, 
    0.03027036, 0.03238663, 0.0347597, 0.03701727, 0.03891977, 0.04041893, 
    0.04187569, 0.04334076, 0.04376047, 0.042658, 0.04119175, 0.03962855,
  0.03777961, 0.03486234, 0.03180903, 0.02920298, 0.02693239, 0.02547367, 
    0.02390613, 0.02356504, 0.02511982, 0.0254573, 0.03801426, 0.04528654, 
    0.04376829, 0.04831244, 0.04900077, 0.04289374, 0.0448246, 0.05219474, 
    0.05473434, 0.05320421, 0.0502604, 0.0497435, 0.05339919, 0.05275194, 
    0.04794987, 0.05392912, 0.04496509, 0.04701335, 0.05422916, 0.05530155, 
    0.04559386, 0.03979766, 0.03409839, 0.03194332, 0.02952582, 0.02642136, 
    0.02576542, 0.02622986, 0.02850889, 0.03298267, 0.03744656, 0.03876941, 
    0.0371616, 0.03675393, 0.03729251, 0.03604449, 0.03426803, 0.03441014, 
    0.03493753, 0.03489649, 0.03411481, 0.03383804, 0.034059, 0.03383894, 
    0.03392791, 0.03463673, 0.03670856, 0.03666013, 0.03514324, 0.03506121, 
    0.03603133, 0.03466595, 0.03379807, 0.03469584, 0.03451895, 0.03407198, 
    0.03382417, 0.03391797, 0.03447868, 0.03465868, 0.03535163, 0.03429162, 
    0.03201566, 0.03054162, 0.0302716, 0.02981649, 0.02969145, 0.02906433, 
    0.02854467, 0.02896794, 0.02832506, 0.0272354, 0.0255966, 0.02447683, 
    0.0241112, 0.02269953, 0.02106795, 0.01881708, 0.01749783, 0.01630295, 
    0.01495729, 0.0137419, 0.01296198, 0.01312511, 0.01345743, 0.0140027, 
    0.01531211, 0.01553972, 0.01508815, 0.01642262, 0.01813946, 0.01923143, 
    0.01922236, 0.01963933, 0.01903941, 0.01907692, 0.01888556, 0.02066012, 
    0.0240244, 0.02610185, 0.02514808, 0.02379328, 0.02401371, 0.02602442, 
    0.03056453, 0.0308183, 0.03477234, 0.04250447, 0.04707152, 0.05763844, 
    0.05244981, 0.04557348, 0.04426701, 0.04914695, 0.05566271, 0.06025765, 
    0.06336274, 0.06283993, 0.06234228, 0.06340435, 0.06388797, 0.06597619, 
    0.06648238, 0.06648047, 0.06692347, 0.0686885, 0.067453, 0.06725949, 
    0.06515297, 0.06087463, 0.05878754, 0.05617794, 0.05251748, 0.05035304, 
    0.04822376, 0.04712398, 0.04810939, 0.0475623, 0.04380496, 0.04185569, 
    0.04070746, 0.03764618, 0.03461853, 0.03149075, 0.02936226, 0.02791338, 
    0.02798594, 0.02812934, 0.02775287, 0.02692284, 0.02582229, 0.02505983, 
    0.02454288, 0.02425071, 0.02456437, 0.02330591, 0.02135629, 0.01979584, 
    0.01810198, 0.01708025, 0.01686206, 0.0166746, 0.01554406, 0.01622989, 
    0.01787189, 0.01750463, 0.01758474, 0.01793554, 0.01652435, 0.01499279, 
    0.01484172, 0.0152144, 0.0154632, 0.01555644, 0.01432041, 0.01325481, 
    0.01270338, 0.0129405, 0.01317874, 0.01333216, 0.01356876, 0.01416126, 
    0.01420177, 0.01446043, 0.01490989, 0.01480342, 0.01471888, 0.01438133, 
    0.01461432, 0.0153415, 0.01650225, 0.01800954, 0.01954149, 0.02164695, 
    0.02359565, 0.02554495, 0.02836846, 0.03162023, 0.0342262, 0.03716632, 
    0.03921502, 0.04072463, 0.04209796, 0.04212775, 0.04248287, 0.04277281, 
    0.04194127, 0.04009737, 0.03786587, 0.03581696, 0.03228882, 0.02890689, 
    0.02049924, 0.01062863, 0.01107613, 0.03533061, 0.09462909, 0.1437356, 
    0.0968252, 0.08041043, 0.06534827, 0.05841433, 0.05222129, 0.04905873, 
    0.0472631, 0.04905039, 0.05114717, 0.05367472, 0.0565888, 0.05814872, 
    0.05680412, 0.05530395, 0.05597663, 0.05199485, 0.04877963, 0.0457839, 
    0.0435193, 0.04431358, 0.04673971, 0.04739689, 0.04215307, 0.04093539, 
    0.04405599, 0.03895662, 0.03294208, 0.03825974, 0.03699326, 0.03854879, 
    0.03246901, 0.02239986, 0.01890182, 0.01616873, 0.01546504, 0.01591303, 
    0.01670205, 0.01703082, 0.016592, 0.016796, 0.01713291, 0.01773032, 
    0.01881089, 0.01995606, 0.02132274, 0.0227087, 0.02418352, 0.02600167, 
    0.0277062, 0.02973564, 0.03196495, 0.03407931, 0.03659906, 0.03836817, 
    0.0403255, 0.0422106, 0.04239566, 0.04091593, 0.03979975, 0.03922258,
  0.03697853, 0.03456987, 0.03191122, 0.02920529, 0.02686938, 0.02548641, 
    0.02437004, 0.02416392, 0.02571667, 0.02624517, 0.03641636, 0.04569927, 
    0.0445573, 0.04883794, 0.04916116, 0.0453894, 0.04912983, 0.05253093, 
    0.050449, 0.04963802, 0.05274182, 0.05018884, 0.05154691, 0.05461045, 
    0.05227516, 0.0535803, 0.04482502, 0.04920565, 0.0728175, 0.0510009, 
    0.04391587, 0.03526955, 0.0329565, 0.03202536, 0.03185679, 0.02890828, 
    0.02807294, 0.02847214, 0.02884901, 0.03109895, 0.03445924, 0.03482472, 
    0.03364362, 0.0342303, 0.03650662, 0.03630437, 0.03496158, 0.03530335, 
    0.03495738, 0.03524891, 0.03471504, 0.03387226, 0.0338706, 0.03432399, 
    0.03558401, 0.03674855, 0.03840862, 0.0375266, 0.03603273, 0.03607021, 
    0.03608341, 0.03501831, 0.03370511, 0.0334604, 0.03319582, 0.03293982, 
    0.03230911, 0.03286073, 0.03405083, 0.03470229, 0.03493397, 0.03453876, 
    0.03198826, 0.02929078, 0.0281457, 0.02700272, 0.02624554, 0.02480494, 
    0.02381014, 0.0238817, 0.02418053, 0.02393166, 0.02278677, 0.02239741, 
    0.0224512, 0.0216712, 0.02103486, 0.02051673, 0.02105043, 0.01929684, 
    0.0171233, 0.0157749, 0.01491005, 0.01513545, 0.01442006, 0.01582921, 
    0.01660431, 0.01488306, 0.01539728, 0.01756791, 0.02082138, 0.01961485, 
    0.01896674, 0.01950208, 0.02024074, 0.02110215, 0.02106671, 0.02262437, 
    0.02355037, 0.02467697, 0.0252788, 0.02569774, 0.02747091, 0.03357383, 
    0.03950573, 0.03698409, 0.04558649, 0.05915711, 0.06382871, 0.05819725, 
    0.05333719, 0.04974179, 0.04826624, 0.04996998, 0.05642509, 0.06022453, 
    0.06036006, 0.05990446, 0.06326409, 0.06714997, 0.06778838, 0.06692493, 
    0.0658428, 0.06620675, 0.06589423, 0.06632616, 0.0647992, 0.06421018, 
    0.06267314, 0.06064869, 0.05764574, 0.0532908, 0.04850749, 0.04667449, 
    0.04544551, 0.04385008, 0.04383137, 0.04308023, 0.04102849, 0.03976013, 
    0.03788407, 0.03599711, 0.03370637, 0.03080785, 0.02832955, 0.0267712, 
    0.02632935, 0.02569236, 0.0246508, 0.02357626, 0.02329684, 0.02278866, 
    0.02270122, 0.02238283, 0.02113774, 0.01986933, 0.01900226, 0.0171787, 
    0.0156196, 0.01509567, 0.01492111, 0.01512397, 0.01559587, 0.01660634, 
    0.01750071, 0.01672197, 0.0173646, 0.01885034, 0.01690089, 0.01500419, 
    0.01451937, 0.01456973, 0.01584945, 0.01784375, 0.01650087, 0.01435958, 
    0.01362053, 0.01328941, 0.01321824, 0.01314494, 0.01335024, 0.01401529, 
    0.01411155, 0.01409062, 0.01444759, 0.01448921, 0.01423246, 0.01414614, 
    0.01439356, 0.01512372, 0.01636038, 0.01789152, 0.01959292, 0.02119602, 
    0.02275569, 0.02497626, 0.02749934, 0.03044192, 0.03304298, 0.03637274, 
    0.03833374, 0.03977513, 0.04071159, 0.04103138, 0.04115548, 0.04120607, 
    0.0398761, 0.0383542, 0.0365867, 0.03376108, 0.03019565, 0.02535902, 
    0.0163019, 0.01017105, 0.02091132, 0.06449201, 0.1239362, 0.1297764, 
    0.09042368, 0.06441171, 0.05366633, 0.05273742, 0.05037632, 0.0490426, 
    0.04824718, 0.04998954, 0.05195786, 0.0543428, 0.05736521, 0.058082, 
    0.05844673, 0.0593911, 0.05946308, 0.05400675, 0.0505902, 0.04806706, 
    0.04528432, 0.04630939, 0.04676368, 0.04651559, 0.04192406, 0.03952511, 
    0.03979502, 0.04062006, 0.03797964, 0.03686409, 0.03272602, 0.0339308, 
    0.04632644, 0.03546029, 0.02374596, 0.01894371, 0.0168745, 0.01676147, 
    0.01758571, 0.01778712, 0.01752821, 0.01777392, 0.01787838, 0.01789591, 
    0.01822112, 0.01900579, 0.01969181, 0.02094365, 0.02234739, 0.02418323, 
    0.0255738, 0.02735695, 0.02929956, 0.03181129, 0.03440712, 0.03655051, 
    0.03836079, 0.04054476, 0.04072788, 0.0396611, 0.03899707, 0.0382298,
  0.03575835, 0.03413881, 0.03216938, 0.02984145, 0.02800251, 0.02650119, 
    0.02572676, 0.0258378, 0.02716212, 0.02901812, 0.03931527, 0.04955111, 
    0.05014, 0.05501343, 0.05439851, 0.04981045, 0.05159785, 0.05196014, 
    0.04870563, 0.04804659, 0.05311194, 0.05534385, 0.05327202, 0.05011186, 
    0.04766705, 0.05054717, 0.04024673, 0.04513488, 0.066043, 0.05477131, 
    0.04270754, 0.03494619, 0.03151435, 0.02974711, 0.02998375, 0.02871585, 
    0.02864033, 0.02821196, 0.02809829, 0.02932597, 0.03013499, 0.03037677, 
    0.03003029, 0.03221425, 0.03416963, 0.03518101, 0.03640698, 0.03915675, 
    0.0362438, 0.03521639, 0.03566374, 0.03598532, 0.03653882, 0.03661779, 
    0.03865495, 0.03990853, 0.03997116, 0.0388999, 0.03637256, 0.03586983, 
    0.0349818, 0.03475578, 0.03455165, 0.03425289, 0.03490955, 0.03518183, 
    0.03406494, 0.03436986, 0.03569054, 0.03523428, 0.03509163, 0.0350305, 
    0.03269659, 0.03016896, 0.02814018, 0.02648168, 0.02511238, 0.02380635, 
    0.02272938, 0.02201472, 0.02227384, 0.02282915, 0.02203686, 0.02179626, 
    0.02320519, 0.02418994, 0.02598251, 0.02624421, 0.0286418, 0.028459, 
    0.02918109, 0.02511222, 0.0173969, 0.01990318, 0.01966733, 0.01870301, 
    0.01816644, 0.01635201, 0.01785457, 0.02065515, 0.02026069, 0.02053527, 
    0.01980125, 0.02133047, 0.02198005, 0.02188816, 0.02351615, 0.02425047, 
    0.02409187, 0.02429742, 0.02627332, 0.0312271, 0.04010949, 0.05026059, 
    0.05882866, 0.05726496, 0.06663499, 0.09143805, 0.07986571, 0.06465331, 
    0.059789, 0.05915273, 0.05667485, 0.05618672, 0.06042207, 0.06330228, 
    0.06315535, 0.06494334, 0.06650286, 0.07097001, 0.07005565, 0.06503442, 
    0.06337252, 0.06334437, 0.06313179, 0.06325285, 0.06206425, 0.06154634, 
    0.06036821, 0.05931552, 0.05582445, 0.04880048, 0.04463495, 0.04573625, 
    0.04513161, 0.04115888, 0.03907697, 0.03820544, 0.03786253, 0.0361715, 
    0.034247, 0.03287963, 0.03138348, 0.02872968, 0.02645679, 0.02491311, 
    0.02431953, 0.02253385, 0.02050804, 0.0199612, 0.02061497, 0.02066999, 
    0.02110657, 0.02076631, 0.0197417, 0.01841168, 0.01683638, 0.01506877, 
    0.01440546, 0.01406285, 0.01359493, 0.0134783, 0.01418535, 0.01556902, 
    0.01601452, 0.01697931, 0.01739426, 0.01852529, 0.01679613, 0.0160167, 
    0.01478655, 0.01429679, 0.01497322, 0.01631514, 0.01615474, 0.01589925, 
    0.0155347, 0.01462744, 0.01420166, 0.01345656, 0.01366905, 0.01489876, 
    0.01544693, 0.01519534, 0.01503881, 0.01493437, 0.01423872, 0.01416158, 
    0.01479399, 0.01556159, 0.01673284, 0.01779098, 0.01894037, 0.02037848, 
    0.02216421, 0.02432476, 0.02665528, 0.02923393, 0.03251302, 0.03557765, 
    0.03790896, 0.03976705, 0.0405101, 0.04077842, 0.0409787, 0.04081795, 
    0.03934493, 0.03728923, 0.03525003, 0.03281274, 0.0287335, 0.02183601, 
    0.01416848, 0.01354077, 0.03804784, 0.0802568, 0.1368025, 0.1049095, 
    0.07957564, 0.05738157, 0.05183366, 0.05180987, 0.04979891, 0.04966881, 
    0.05139569, 0.0526316, 0.05310005, 0.05508714, 0.0571074, 0.05813513, 
    0.06066922, 0.06473007, 0.06323055, 0.05825516, 0.05641387, 0.05349156, 
    0.04988715, 0.04857394, 0.04790016, 0.04755756, 0.0432948, 0.0402364, 
    0.04098668, 0.04568169, 0.04816903, 0.04716994, 0.04514906, 0.04059403, 
    0.04927631, 0.04835478, 0.02657236, 0.02166523, 0.01867981, 0.01827248, 
    0.01847384, 0.01812644, 0.01807705, 0.01842414, 0.01821884, 0.01844677, 
    0.0187638, 0.01913003, 0.01934765, 0.02031433, 0.02113963, 0.02227025, 
    0.02330441, 0.02469217, 0.02673046, 0.02923539, 0.03183549, 0.03396333, 
    0.03588527, 0.03815001, 0.03885647, 0.03828182, 0.03813324, 0.03721977,
  0.03493152, 0.0339125, 0.03243966, 0.03056847, 0.02926255, 0.02816563, 
    0.02770035, 0.02829272, 0.02979407, 0.03390556, 0.04468679, 0.0562759, 
    0.05959613, 0.06719816, 0.06284668, 0.05212026, 0.05346792, 0.05202274, 
    0.04976676, 0.04800522, 0.05033496, 0.05770066, 0.05463898, 0.05050221, 
    0.04733623, 0.05024038, 0.04259187, 0.0380149, 0.05293625, 0.05399632, 
    0.04428679, 0.03724948, 0.03174035, 0.02860681, 0.02799018, 0.02748857, 
    0.02749402, 0.02720486, 0.02605573, 0.02602153, 0.02644871, 0.02665981, 
    0.02784117, 0.03035853, 0.03109873, 0.03231356, 0.03567149, 0.03726162, 
    0.03597855, 0.03588514, 0.03614109, 0.03718022, 0.03741917, 0.0384098, 
    0.04067836, 0.041081, 0.03924544, 0.03784383, 0.03619791, 0.03608525, 
    0.03550641, 0.03520196, 0.03589756, 0.03565565, 0.03643304, 0.03701982, 
    0.03638188, 0.03805325, 0.039202, 0.03689273, 0.0369991, 0.03697493, 
    0.03376215, 0.03039855, 0.02833113, 0.02634603, 0.02485699, 0.02369907, 
    0.02382063, 0.02352091, 0.02339613, 0.02356297, 0.02310884, 0.02412574, 
    0.02824794, 0.03905322, 0.04111297, 0.03999716, 0.0494557, 0.04221318, 
    0.03153486, 0.02393954, 0.01770869, 0.01818828, 0.01893118, 0.01814026, 
    0.0170902, 0.01738512, 0.01755231, 0.01937926, 0.02065542, 0.02202342, 
    0.02184104, 0.0224511, 0.02184977, 0.02370824, 0.02679701, 0.02734007, 
    0.02804626, 0.03030602, 0.03582665, 0.05020423, 0.0628721, 0.07672398, 
    0.103355, 0.1152726, 0.110388, 0.09728608, 0.08856943, 0.07259589, 
    0.06914875, 0.07026814, 0.06753159, 0.06533447, 0.06566404, 0.06798816, 
    0.06833789, 0.07156541, 0.07049105, 0.07064754, 0.06895746, 0.06470983, 
    0.06365329, 0.06215328, 0.06096834, 0.06173521, 0.06130951, 0.05990684, 
    0.0578942, 0.05607929, 0.05282942, 0.04755462, 0.04422181, 0.04485912, 
    0.04289237, 0.03895188, 0.03643923, 0.03456806, 0.03371397, 0.03250587, 
    0.02969907, 0.028361, 0.02752875, 0.02676223, 0.02441551, 0.02265649, 
    0.02166023, 0.02024226, 0.01917412, 0.01933206, 0.01973186, 0.01971976, 
    0.02003523, 0.01914733, 0.0184361, 0.01698028, 0.01574348, 0.0147803, 
    0.0141435, 0.01334189, 0.01243552, 0.0123557, 0.01265133, 0.01430221, 
    0.01547412, 0.01575837, 0.01500107, 0.01441762, 0.01543356, 0.01635884, 
    0.01581654, 0.01516131, 0.01491368, 0.0150248, 0.01547577, 0.01609395, 
    0.01597195, 0.01609499, 0.01557237, 0.01463644, 0.01464608, 0.01565245, 
    0.01696924, 0.01684707, 0.01682534, 0.01671659, 0.01625962, 0.01594235, 
    0.01547082, 0.01618499, 0.01738572, 0.01797414, 0.01897347, 0.02042574, 
    0.02191854, 0.02370558, 0.02596023, 0.0289987, 0.03286117, 0.0356982, 
    0.03809317, 0.04058481, 0.0411041, 0.04179611, 0.04187233, 0.04085206, 
    0.03909859, 0.03685381, 0.03465833, 0.03219711, 0.02792686, 0.0207914, 
    0.01614321, 0.02872266, 0.07100279, 0.09287656, 0.1134454, 0.08367833, 
    0.06754008, 0.05433488, 0.05297858, 0.05325281, 0.05315908, 0.05443067, 
    0.05656248, 0.05688726, 0.05608822, 0.05734748, 0.05976924, 0.06240494, 
    0.06634746, 0.0705715, 0.06858398, 0.06656303, 0.06494103, 0.06089393, 
    0.05671112, 0.05180652, 0.05151025, 0.05125643, 0.04666752, 0.04436903, 
    0.04801123, 0.05690412, 0.05950789, 0.05779184, 0.06166842, 0.05099192, 
    0.03715068, 0.03964629, 0.02717237, 0.02377256, 0.02103703, 0.02054937, 
    0.01980546, 0.01888639, 0.01835096, 0.01832205, 0.01829815, 0.0182753, 
    0.01840095, 0.01878531, 0.01890441, 0.01966614, 0.02040765, 0.02102954, 
    0.02217968, 0.02345667, 0.0254486, 0.0270722, 0.02933916, 0.03142175, 
    0.03322164, 0.03507682, 0.03616505, 0.03642191, 0.03598673, 0.03557087,
  0.03487334, 0.03424211, 0.03311295, 0.03227409, 0.03138405, 0.03076926, 
    0.0304852, 0.03256394, 0.03515086, 0.042187, 0.05248145, 0.06300046, 
    0.06876102, 0.07448072, 0.06578833, 0.05440881, 0.05430818, 0.05164987, 
    0.05080842, 0.04991474, 0.04823094, 0.05461124, 0.05464148, 0.04603402, 
    0.0500218, 0.05302415, 0.04500199, 0.04603022, 0.03903724, 0.05164977, 
    0.04667848, 0.03852282, 0.03232459, 0.02718713, 0.02582045, 0.02640964, 
    0.02735149, 0.0273841, 0.02530195, 0.0243631, 0.02558751, 0.02505798, 
    0.0251744, 0.02618715, 0.02733668, 0.02849779, 0.03087328, 0.03299877, 
    0.03414128, 0.03453249, 0.03448509, 0.0360889, 0.03679821, 0.03863684, 
    0.04108057, 0.03925335, 0.03761694, 0.03659048, 0.03597129, 0.03667458, 
    0.03730236, 0.03659585, 0.036339, 0.03566639, 0.03736146, 0.03786367, 
    0.03708976, 0.03882173, 0.03946749, 0.03850199, 0.03887163, 0.04000615, 
    0.03672893, 0.03217656, 0.03038064, 0.02817372, 0.02535013, 0.02416148, 
    0.0249149, 0.02568357, 0.02512293, 0.0262567, 0.02935095, 0.03097467, 
    0.03646186, 0.050191, 0.04661267, 0.03871201, 0.04066421, 0.03631268, 
    0.02834515, 0.0240422, 0.02079649, 0.02009708, 0.01966602, 0.01810832, 
    0.01761162, 0.01769995, 0.01814478, 0.01932398, 0.0211284, 0.02251904, 
    0.0229095, 0.02293628, 0.02406421, 0.0262876, 0.02870896, 0.03194033, 
    0.03131299, 0.03686193, 0.053661, 0.08165934, 0.1055818, 0.1324933, 
    0.1564011, 0.1670117, 0.1388515, 0.1285713, 0.09041059, 0.07510005, 
    0.07858011, 0.0842769, 0.08273396, 0.07324641, 0.07179131, 0.07495324, 
    0.07704569, 0.07498824, 0.07230563, 0.06799788, 0.06382636, 0.06265096, 
    0.06263042, 0.05909826, 0.05758693, 0.05855808, 0.05987466, 0.05798012, 
    0.05530112, 0.05296357, 0.04947794, 0.04612261, 0.04318207, 0.04225147, 
    0.04027566, 0.03685948, 0.03302168, 0.03079154, 0.02971289, 0.02778285, 
    0.0255493, 0.02490872, 0.02526244, 0.02490434, 0.02214367, 0.02052785, 
    0.01962346, 0.01893835, 0.01831631, 0.01821481, 0.01842061, 0.01789454, 
    0.0167248, 0.01612725, 0.01589778, 0.01546905, 0.01497783, 0.01487104, 
    0.0145294, 0.01443165, 0.01334547, 0.01320374, 0.01355123, 0.01369258, 
    0.01405852, 0.01410829, 0.01389337, 0.01404078, 0.01494752, 0.01489522, 
    0.01535952, 0.01522835, 0.01544028, 0.01573941, 0.01661685, 0.01688481, 
    0.01706063, 0.01762425, 0.01744497, 0.0171039, 0.01695431, 0.01742186, 
    0.01846762, 0.0187093, 0.01881083, 0.01880432, 0.018681, 0.01879579, 
    0.01852379, 0.01865177, 0.0195336, 0.01981211, 0.02024075, 0.02165488, 
    0.02347797, 0.02464296, 0.0263227, 0.02938317, 0.03232143, 0.03486868, 
    0.03684926, 0.03938115, 0.04097284, 0.04225944, 0.04216857, 0.04086305, 
    0.038932, 0.03742337, 0.03517096, 0.03217719, 0.02738623, 0.02272283, 
    0.02238781, 0.05124058, 0.07930399, 0.09891617, 0.08294417, 0.07408072, 
    0.06286363, 0.05565285, 0.0565678, 0.05882927, 0.06157094, 0.06243389, 
    0.06237647, 0.06151182, 0.06238007, 0.06369664, 0.06452898, 0.06754201, 
    0.07202365, 0.07425182, 0.0741992, 0.07383427, 0.06961948, 0.06531996, 
    0.06003425, 0.05519921, 0.0561984, 0.0558068, 0.05100444, 0.05193954, 
    0.0606801, 0.07178632, 0.06727889, 0.06072675, 0.0644676, 0.05117049, 
    0.02991548, 0.03262377, 0.02934365, 0.02707523, 0.02493127, 0.02376842, 
    0.02252438, 0.0213567, 0.01981815, 0.01908465, 0.01892136, 0.01830819, 
    0.01813469, 0.0185447, 0.01850833, 0.01912292, 0.02011804, 0.02100899, 
    0.02252097, 0.02394878, 0.02482075, 0.02580002, 0.02719607, 0.02889542, 
    0.0309225, 0.03290287, 0.03468833, 0.03492293, 0.03492472, 0.03473541,
  0.03564094, 0.03554423, 0.03477551, 0.03429584, 0.03385805, 0.03390836, 
    0.03424655, 0.03734693, 0.04327977, 0.05369688, 0.06632914, 0.07408176, 
    0.07401963, 0.07288881, 0.06446843, 0.05608709, 0.05515351, 0.05394955, 
    0.05426733, 0.05398351, 0.05148677, 0.05630549, 0.05586204, 0.05125744, 
    0.05784165, 0.05724708, 0.05053721, 0.04601223, 0.0415171, 0.05188767, 
    0.0477555, 0.03903967, 0.03228416, 0.02546328, 0.0241234, 0.0237765, 
    0.02419088, 0.02476695, 0.0241401, 0.02500097, 0.02590966, 0.02457557, 
    0.02319551, 0.02313597, 0.02442757, 0.02533401, 0.02644566, 0.02903861, 
    0.02969746, 0.02919638, 0.03003951, 0.03241001, 0.03402122, 0.03564642, 
    0.04027359, 0.0381077, 0.03562189, 0.03379896, 0.03329242, 0.03317888, 
    0.03394966, 0.03324625, 0.03333429, 0.03369116, 0.03680499, 0.03777702, 
    0.0382434, 0.03981276, 0.03887969, 0.0384066, 0.03796675, 0.04047117, 
    0.03876431, 0.0349406, 0.03304584, 0.0313651, 0.02854862, 0.02728002, 
    0.0284867, 0.02966142, 0.03048539, 0.03674082, 0.04400611, 0.05133343, 
    0.04815916, 0.03979129, 0.03272124, 0.03135058, 0.03139551, 0.0281516, 
    0.02645889, 0.02590639, 0.02399093, 0.02179175, 0.01946276, 0.02063217, 
    0.02089236, 0.0228906, 0.02292414, 0.02200288, 0.02160028, 0.02343845, 
    0.02415262, 0.02440519, 0.02612787, 0.0284633, 0.03213723, 0.03865615, 
    0.05149431, 0.0792221, 0.1115273, 0.129431, 0.1506341, 0.1881483, 
    0.1975873, 0.1739022, 0.1367363, 0.1071241, 0.07701308, 0.07110598, 
    0.08176082, 0.08904488, 0.08780589, 0.07918087, 0.07604201, 0.07994033, 
    0.07951773, 0.07660802, 0.07200847, 0.0649059, 0.05988119, 0.05879939, 
    0.05657474, 0.05219296, 0.05300033, 0.05396058, 0.05541798, 0.05317667, 
    0.05154993, 0.04970482, 0.04539604, 0.04078129, 0.03805178, 0.03786828, 
    0.03766446, 0.0360055, 0.03190207, 0.02861207, 0.02695393, 0.02562061, 
    0.02350109, 0.02339045, 0.02302819, 0.02246287, 0.02103089, 0.01979217, 
    0.0187241, 0.01759344, 0.01683951, 0.01671997, 0.01663326, 0.01563233, 
    0.01449376, 0.01389069, 0.01394355, 0.01399298, 0.01442469, 0.01515974, 
    0.01522974, 0.01566562, 0.01549112, 0.01509832, 0.0150978, 0.01427483, 
    0.01415207, 0.01412703, 0.01401612, 0.01413545, 0.01407283, 0.0140471, 
    0.01490198, 0.01509247, 0.01551452, 0.01624813, 0.01788719, 0.01815678, 
    0.01836339, 0.01904672, 0.01978737, 0.02008346, 0.02010948, 0.02076653, 
    0.02050852, 0.02027856, 0.02036118, 0.02090435, 0.02125556, 0.02141947, 
    0.02141156, 0.02145418, 0.02192584, 0.02214232, 0.02259781, 0.02353513, 
    0.0253821, 0.02585921, 0.02681415, 0.02917434, 0.03167664, 0.0339183, 
    0.0347746, 0.03618319, 0.03839235, 0.03990213, 0.03991544, 0.03946123, 
    0.03901706, 0.03828633, 0.03539785, 0.03197788, 0.0273182, 0.02768897, 
    0.03320754, 0.06885754, 0.07324846, 0.08948622, 0.07726973, 0.07676837, 
    0.06694998, 0.06323689, 0.06449677, 0.06791856, 0.07005854, 0.06990941, 
    0.06843717, 0.06709477, 0.06720167, 0.0684754, 0.06940895, 0.07197369, 
    0.07384783, 0.07387713, 0.07553254, 0.07458115, 0.07017479, 0.06622846, 
    0.06361435, 0.06152099, 0.06295392, 0.06051871, 0.05499098, 0.05980646, 
    0.07076139, 0.0799823, 0.0663214, 0.05127314, 0.04979815, 0.03876797, 
    0.0262391, 0.02821489, 0.03140304, 0.02913081, 0.02719777, 0.02561441, 
    0.0247818, 0.02411393, 0.02294516, 0.0210884, 0.02062686, 0.01977938, 
    0.01945723, 0.01944649, 0.01941584, 0.01982132, 0.02099012, 0.0220537, 
    0.02273585, 0.02366723, 0.02428519, 0.02468977, 0.02598112, 0.02722827, 
    0.02918248, 0.03143714, 0.03373698, 0.0345887, 0.03468323, 0.03503968,
  0.03694466, 0.0382422, 0.03795723, 0.03870073, 0.03923833, 0.03988134, 
    0.04144657, 0.04642914, 0.05566603, 0.07567552, 0.08328536, 0.08558458, 
    0.07961488, 0.07070976, 0.06410881, 0.0591481, 0.05789498, 0.05788683, 
    0.0591541, 0.05962382, 0.06244728, 0.07126341, 0.07064586, 0.06011312, 
    0.06909812, 0.06850331, 0.06375666, 0.04961316, 0.04420176, 0.04526794, 
    0.0439272, 0.03857789, 0.03166983, 0.02435919, 0.02257728, 0.02195682, 
    0.02143321, 0.02196993, 0.02332888, 0.02489093, 0.02504998, 0.02208346, 
    0.02044763, 0.02059447, 0.02144326, 0.02213634, 0.02391349, 0.02500308, 
    0.02490144, 0.02523256, 0.02557583, 0.0277306, 0.02879108, 0.02970371, 
    0.03175205, 0.03229538, 0.03000076, 0.02783139, 0.02766455, 0.02951054, 
    0.02954867, 0.02791546, 0.0285156, 0.02896202, 0.03198916, 0.03512764, 
    0.03745586, 0.03824089, 0.03726198, 0.03764084, 0.03675796, 0.03791739, 
    0.03713306, 0.03498738, 0.03499179, 0.033812, 0.0322038, 0.03432335, 
    0.03620872, 0.03793969, 0.04305101, 0.0571094, 0.06784124, 0.071651, 
    0.05405298, 0.0356577, 0.03091435, 0.02895311, 0.0279424, 0.02708209, 
    0.02693988, 0.02734493, 0.02559485, 0.02303627, 0.02339788, 0.02681139, 
    0.02952421, 0.03304961, 0.02959393, 0.02536377, 0.02543741, 0.02826388, 
    0.02824329, 0.02845673, 0.0295019, 0.03348583, 0.04121254, 0.05373334, 
    0.09844673, 0.1618935, 0.1876701, 0.1662115, 0.1508648, 0.1596777, 
    0.1591933, 0.1273834, 0.1003589, 0.08006404, 0.06472678, 0.06801056, 
    0.07889608, 0.08186914, 0.08113743, 0.07640966, 0.07682096, 0.07793424, 
    0.07453372, 0.07047578, 0.06773381, 0.06195152, 0.05584181, 0.05283869, 
    0.04894016, 0.04623357, 0.0467888, 0.04845846, 0.04860222, 0.04651154, 
    0.04542462, 0.04210504, 0.03800364, 0.03638228, 0.03473695, 0.0336863, 
    0.03212356, 0.02982416, 0.02696121, 0.02415709, 0.02255841, 0.02166355, 
    0.02026393, 0.01960226, 0.0192065, 0.01932775, 0.01951219, 0.0188668, 
    0.01762787, 0.01642963, 0.01585666, 0.01582276, 0.01548431, 0.01523542, 
    0.0147188, 0.01412731, 0.01368858, 0.01431117, 0.01583792, 0.01722993, 
    0.01779729, 0.01754242, 0.01663878, 0.01578317, 0.01594065, 0.01532904, 
    0.01530369, 0.01433366, 0.0139006, 0.0138479, 0.01353279, 0.01369191, 
    0.01412251, 0.01408967, 0.01459097, 0.01592986, 0.01731918, 0.01811192, 
    0.0191055, 0.02018061, 0.02083416, 0.02093315, 0.02129865, 0.0223824, 
    0.0223666, 0.02190669, 0.02110348, 0.02231758, 0.02328908, 0.02286435, 
    0.02260336, 0.02245151, 0.02359861, 0.02444608, 0.02479326, 0.02572529, 
    0.02689889, 0.02708943, 0.02729824, 0.02849843, 0.03019892, 0.03212212, 
    0.03249557, 0.03240925, 0.0340084, 0.03539319, 0.03633656, 0.03734212, 
    0.03810608, 0.03780213, 0.03551304, 0.03170596, 0.02832934, 0.03627906, 
    0.0471838, 0.09346407, 0.1274338, 0.1067394, 0.1147661, 0.09068668, 
    0.07078975, 0.07233475, 0.07647525, 0.07898542, 0.07784031, 0.07554247, 
    0.07426099, 0.07188267, 0.07088097, 0.07103427, 0.07323387, 0.07321987, 
    0.07318419, 0.07369054, 0.0743476, 0.07192336, 0.07009003, 0.06878358, 
    0.0708608, 0.0724678, 0.07028605, 0.06246411, 0.05576202, 0.06118865, 
    0.06960724, 0.07457945, 0.05706327, 0.03756782, 0.03025248, 0.02615468, 
    0.02502132, 0.02913899, 0.03101897, 0.02871715, 0.02768494, 0.02648357, 
    0.02609829, 0.02632029, 0.02541187, 0.023906, 0.02257684, 0.02115989, 
    0.02044637, 0.0203755, 0.02080154, 0.02155632, 0.02275574, 0.02366046, 
    0.02456659, 0.02521414, 0.02471081, 0.02483477, 0.02625975, 0.02759182, 
    0.02925317, 0.03105704, 0.0328341, 0.03400045, 0.03523461, 0.0357913,
  0.0382762, 0.04038275, 0.04230547, 0.04440977, 0.0470889, 0.04978958, 
    0.05368901, 0.060885, 0.07908836, 0.1005865, 0.1034366, 0.09433055, 
    0.08146201, 0.07184997, 0.06755377, 0.06434916, 0.0624712, 0.06224139, 
    0.06528851, 0.07022974, 0.08291967, 0.1020621, 0.09276504, 0.0688585, 
    0.07485193, 0.07760081, 0.07638754, 0.05772716, 0.04748695, 0.04741462, 
    0.04240557, 0.03845928, 0.02999533, 0.02263326, 0.02080789, 0.02027641, 
    0.02019605, 0.02079702, 0.02246584, 0.02272595, 0.02086761, 0.01857929, 
    0.01809125, 0.0186678, 0.01873546, 0.01963213, 0.02127696, 0.02248179, 
    0.0227478, 0.02364595, 0.02515753, 0.0286979, 0.02869077, 0.02786159, 
    0.02800424, 0.02864554, 0.02671114, 0.02516153, 0.02475309, 0.0255043, 
    0.02688787, 0.02583218, 0.02514235, 0.02605193, 0.02830887, 0.03038382, 
    0.03089566, 0.03252708, 0.0340513, 0.03616768, 0.03565325, 0.03564529, 
    0.03482841, 0.03429612, 0.0364255, 0.03734102, 0.03638995, 0.03933481, 
    0.04279965, 0.04806173, 0.06245995, 0.0788668, 0.08825094, 0.07656065, 
    0.05346042, 0.03360535, 0.02976752, 0.02858766, 0.03026194, 0.03369871, 
    0.03470335, 0.03593819, 0.03176574, 0.02809714, 0.03534209, 0.05908957, 
    0.062336, 0.06213625, 0.03500351, 0.02937021, 0.0314314, 0.03473974, 
    0.03388861, 0.03325353, 0.03355686, 0.03959068, 0.05417973, 0.06721823, 
    0.1247521, 0.1934718, 0.2045083, 0.1593876, 0.1289631, 0.1054529, 
    0.08464123, 0.06854398, 0.05827199, 0.05473001, 0.05678838, 0.06281763, 
    0.07131384, 0.07405102, 0.07237827, 0.07131662, 0.06935518, 0.06890437, 
    0.06919795, 0.06591197, 0.06120654, 0.05731682, 0.05231298, 0.04860625, 
    0.04421, 0.04202429, 0.04188424, 0.04173386, 0.04018677, 0.03846913, 
    0.0369063, 0.03386238, 0.03108241, 0.02904116, 0.02788422, 0.02676966, 
    0.02486212, 0.02276846, 0.02170303, 0.02077538, 0.02003362, 0.01887663, 
    0.01772726, 0.01670622, 0.01628451, 0.01683177, 0.01776902, 0.01688593, 
    0.01576019, 0.01506844, 0.01485191, 0.01478402, 0.01497418, 0.0152421, 
    0.01511559, 0.01487513, 0.01481716, 0.01591709, 0.01718114, 0.0171161, 
    0.01681445, 0.01658092, 0.01605617, 0.01534694, 0.01541374, 0.01516416, 
    0.01480051, 0.01388963, 0.01369, 0.01388809, 0.01377963, 0.01351322, 
    0.01395474, 0.01416007, 0.01453501, 0.01528492, 0.01637552, 0.01819474, 
    0.0197282, 0.02008243, 0.02102265, 0.02133114, 0.02068937, 0.02122303, 
    0.02128052, 0.02084341, 0.02063075, 0.02161588, 0.02195239, 0.02114068, 
    0.02061942, 0.02138216, 0.02272294, 0.02361316, 0.02478532, 0.02520581, 
    0.02570741, 0.02648373, 0.02676949, 0.02655299, 0.02750396, 0.0292414, 
    0.02987393, 0.02876156, 0.02877189, 0.02995108, 0.0316228, 0.03353434, 
    0.03578214, 0.03659116, 0.03510501, 0.03184594, 0.0292524, 0.0399374, 
    0.05215508, 0.1243496, 0.1262044, 0.1446105, 0.1330147, 0.09994409, 
    0.07771534, 0.08124233, 0.08881675, 0.09007047, 0.08595379, 0.08214604, 
    0.08021207, 0.07855324, 0.07587928, 0.07463477, 0.07450414, 0.07204553, 
    0.07241935, 0.07529942, 0.07586963, 0.07509999, 0.07147085, 0.07242814, 
    0.07665791, 0.07928644, 0.07496459, 0.06251694, 0.05409707, 0.05461426, 
    0.05343571, 0.05162969, 0.03960741, 0.02613087, 0.02279702, 0.02492555, 
    0.02886153, 0.0310367, 0.03025473, 0.02890582, 0.02798066, 0.02686859, 
    0.02642918, 0.0264152, 0.02495337, 0.02362223, 0.02264654, 0.02174221, 
    0.02091755, 0.02117724, 0.02202699, 0.02280969, 0.02394927, 0.02545263, 
    0.02671127, 0.02634057, 0.02583692, 0.02613478, 0.02716606, 0.02787008, 
    0.02908796, 0.03055617, 0.03232203, 0.03385856, 0.03499023, 0.03627475,
  0.03969647, 0.04300163, 0.04598461, 0.04899006, 0.05370684, 0.05906362, 
    0.06607973, 0.08041007, 0.1078989, 0.121472, 0.1103801, 0.0954961, 
    0.07900711, 0.07176669, 0.0681003, 0.06648468, 0.06417209, 0.06483824, 
    0.06993862, 0.07673551, 0.09584796, 0.1225855, 0.1111212, 0.07212044, 
    0.07000728, 0.0784074, 0.0788694, 0.06438176, 0.05069111, 0.0498029, 
    0.04326764, 0.03372537, 0.02911233, 0.02116129, 0.01940667, 0.01928019, 
    0.01920581, 0.01909841, 0.01913005, 0.01888848, 0.01848438, 0.01764763, 
    0.01712427, 0.01745606, 0.01782916, 0.01777396, 0.01881128, 0.02016427, 
    0.02093821, 0.02275091, 0.02375939, 0.02485129, 0.0257363, 0.02691507, 
    0.02665357, 0.02650443, 0.02497029, 0.02367982, 0.02306764, 0.02350031, 
    0.02406562, 0.02352435, 0.0238109, 0.02453317, 0.02518549, 0.02563316, 
    0.02561466, 0.0269421, 0.02802363, 0.03052412, 0.03200809, 0.03358148, 
    0.03472307, 0.03445196, 0.03616092, 0.03683957, 0.03661733, 0.03941902, 
    0.045752, 0.05783081, 0.07757754, 0.1010161, 0.0918774, 0.06672993, 
    0.04505426, 0.03340741, 0.03203329, 0.03531049, 0.04606872, 0.05321857, 
    0.05862848, 0.05794941, 0.04449917, 0.03525521, 0.05606708, 0.098839, 
    0.08558085, 0.06317693, 0.03889162, 0.02816742, 0.02702859, 0.02905538, 
    0.0318694, 0.03378383, 0.03824168, 0.05611363, 0.07280658, 0.06495827, 
    0.06824373, 0.1031076, 0.1187458, 0.09545632, 0.07639904, 0.05911249, 
    0.04990678, 0.04928797, 0.05221164, 0.05348872, 0.05440559, 0.05635818, 
    0.06017836, 0.06302513, 0.0639153, 0.06122038, 0.05935182, 0.05977867, 
    0.059579, 0.0557877, 0.05252327, 0.04863932, 0.0448553, 0.04093298, 
    0.03662878, 0.03439616, 0.0341361, 0.0343569, 0.03392533, 0.03242612, 
    0.03084905, 0.02772167, 0.02520586, 0.02328862, 0.02195253, 0.02036838, 
    0.01922374, 0.01838417, 0.01804298, 0.01868402, 0.01986801, 0.01976522, 
    0.01712549, 0.0163218, 0.01597828, 0.01651341, 0.01661594, 0.01540738, 
    0.01405189, 0.01378787, 0.01392943, 0.01434485, 0.01523853, 0.01570166, 
    0.01606811, 0.0159227, 0.01595492, 0.01665711, 0.01735057, 0.01675392, 
    0.01596538, 0.0154631, 0.01473786, 0.01425848, 0.01381014, 0.01349495, 
    0.01400091, 0.01339934, 0.01340003, 0.0141691, 0.01429802, 0.01424013, 
    0.01475164, 0.01512155, 0.01510218, 0.01484898, 0.01553614, 0.01739405, 
    0.01754456, 0.01723458, 0.01820416, 0.01872339, 0.01867154, 0.01833866, 
    0.01805578, 0.01829282, 0.01862051, 0.01900429, 0.01902505, 0.01867086, 
    0.01858402, 0.02015099, 0.02195568, 0.0229558, 0.02375579, 0.02405254, 
    0.02371852, 0.02378784, 0.02393793, 0.02397927, 0.02455298, 0.02567758, 
    0.02638943, 0.02584417, 0.02506922, 0.02480566, 0.02683792, 0.02982995, 
    0.0326406, 0.03486012, 0.03407186, 0.03284597, 0.03133163, 0.04167135, 
    0.05367817, 0.1363705, 0.1397548, 0.1489866, 0.1349803, 0.1127423, 
    0.09083549, 0.09261881, 0.09997908, 0.1018746, 0.09514752, 0.0885658, 
    0.08591256, 0.08476973, 0.08292019, 0.07988731, 0.07983439, 0.07767636, 
    0.07944898, 0.08239561, 0.08041541, 0.07738365, 0.07198235, 0.07143985, 
    0.07115945, 0.07021865, 0.0669812, 0.05598596, 0.04611669, 0.04056394, 
    0.03374138, 0.02939977, 0.02455612, 0.02207817, 0.02434047, 0.02787849, 
    0.03067746, 0.03209776, 0.03138878, 0.02962541, 0.02727909, 0.02512528, 
    0.02422692, 0.02336476, 0.02215017, 0.02092221, 0.02036701, 0.0196173, 
    0.01966608, 0.02047997, 0.02103655, 0.02116642, 0.02197916, 0.02390949, 
    0.0256444, 0.02541129, 0.02538793, 0.02530269, 0.026218, 0.02734682, 
    0.02913164, 0.03090546, 0.03245188, 0.0336664, 0.03474759, 0.03679678,
  0.04144642, 0.04484772, 0.04820599, 0.052476, 0.05819209, 0.06512067, 
    0.07459297, 0.1007296, 0.1336126, 0.1252988, 0.1087815, 0.09019716, 
    0.07499489, 0.06938522, 0.06646585, 0.06554845, 0.06384842, 0.06671029, 
    0.07355291, 0.08033129, 0.09998533, 0.1302446, 0.1207896, 0.07580983, 
    0.07402187, 0.08750512, 0.09711254, 0.087062, 0.06046377, 0.06652912, 
    0.04955833, 0.03313785, 0.02803948, 0.02093872, 0.01912349, 0.01989314, 
    0.02046379, 0.01992582, 0.01795106, 0.01796254, 0.01928642, 0.01877195, 
    0.01764657, 0.01750071, 0.01775583, 0.01776295, 0.01824349, 0.01887596, 
    0.01982504, 0.02143069, 0.02190795, 0.02194994, 0.02267791, 0.02411639, 
    0.02525095, 0.02642547, 0.02513007, 0.02446212, 0.02443341, 0.02408451, 
    0.02335065, 0.02269253, 0.0223841, 0.02151701, 0.02153927, 0.02232429, 
    0.02398749, 0.02487861, 0.02432167, 0.02436733, 0.02544423, 0.02828979, 
    0.03108463, 0.03259779, 0.03355171, 0.03618953, 0.03800479, 0.04118764, 
    0.05019063, 0.07084948, 0.08679076, 0.09772561, 0.0801959, 0.05051129, 
    0.03567563, 0.03392106, 0.03706853, 0.05023299, 0.07234931, 0.08004351, 
    0.08292133, 0.07677828, 0.05407217, 0.03780816, 0.05543747, 0.08648252, 
    0.07076576, 0.05333718, 0.03584851, 0.02707452, 0.02466282, 0.02586936, 
    0.02910698, 0.03496124, 0.04853847, 0.08359783, 0.1015244, 0.06138967, 
    0.04265099, 0.04338343, 0.04539152, 0.04165837, 0.0403536, 0.04159333, 
    0.04475991, 0.04771409, 0.04753188, 0.04855396, 0.0518789, 0.05377995, 
    0.05530237, 0.05392912, 0.05211226, 0.05008589, 0.04740098, 0.0470636, 
    0.0469915, 0.04490169, 0.04320828, 0.03997047, 0.04009936, 0.03568359, 
    0.03378323, 0.03286403, 0.03216245, 0.03216631, 0.03100266, 0.02893059, 
    0.02772518, 0.02597152, 0.02359286, 0.02135772, 0.01981591, 0.01852509, 
    0.01793329, 0.01722978, 0.0167395, 0.0172369, 0.01883266, 0.01895672, 
    0.01725189, 0.01749753, 0.01681095, 0.01610511, 0.01611912, 0.01583332, 
    0.01451226, 0.0150244, 0.01574774, 0.01605296, 0.01652514, 0.01695841, 
    0.01704675, 0.01623666, 0.0159428, 0.01704171, 0.01710473, 0.01622909, 
    0.01507252, 0.01410608, 0.01310973, 0.01298436, 0.01311646, 0.01306518, 
    0.01396699, 0.01422056, 0.0149971, 0.01493378, 0.01481531, 0.01519904, 
    0.01527138, 0.01490547, 0.01509906, 0.01465931, 0.01502973, 0.01589638, 
    0.01447621, 0.01361362, 0.01394444, 0.01433926, 0.01525372, 0.01587846, 
    0.01606386, 0.01759716, 0.01759078, 0.01652554, 0.01628949, 0.01658328, 
    0.01736523, 0.01867829, 0.01965293, 0.0205171, 0.02103869, 0.02137961, 
    0.02139548, 0.02148897, 0.02132894, 0.02162126, 0.0225843, 0.02322379, 
    0.02381823, 0.02449298, 0.02439211, 0.02438069, 0.02734307, 0.03160863, 
    0.03361268, 0.03477323, 0.03579187, 0.03675916, 0.03835237, 0.04939943, 
    0.06260584, 0.1473858, 0.1404598, 0.1984071, 0.1309234, 0.1336459, 
    0.1022716, 0.1043097, 0.1099899, 0.1126668, 0.1066467, 0.09825425, 
    0.09269796, 0.08868723, 0.08609302, 0.08356307, 0.08635841, 0.08955904, 
    0.09141212, 0.09373733, 0.08978576, 0.0773825, 0.06579293, 0.06193459, 
    0.06030207, 0.05732282, 0.0531189, 0.04513808, 0.03811883, 0.02972463, 
    0.02350077, 0.02168236, 0.0225363, 0.02391019, 0.02664515, 0.02868378, 
    0.02971901, 0.02923629, 0.02693867, 0.02462146, 0.02276845, 0.02131262, 
    0.01987867, 0.01908451, 0.01854781, 0.01886341, 0.01873495, 0.01778505, 
    0.0177622, 0.01799675, 0.01887252, 0.01972198, 0.02067358, 0.02178462, 
    0.02344709, 0.02357928, 0.02427968, 0.02480804, 0.02583479, 0.0283238, 
    0.03119552, 0.0328052, 0.03405284, 0.03457751, 0.03630761, 0.03856224,
  0.04564964, 0.04918648, 0.05344176, 0.05804072, 0.06382769, 0.07146662, 
    0.0796456, 0.1124855, 0.1453766, 0.1348253, 0.1134031, 0.0899772, 
    0.07366952, 0.06982324, 0.06609782, 0.06577051, 0.06575765, 0.06798378, 
    0.07191719, 0.08002506, 0.09585802, 0.1165006, 0.1152688, 0.07781619, 
    0.07627635, 0.09342211, 0.1151978, 0.1093577, 0.06995356, 0.0790842, 
    0.05299069, 0.03429923, 0.02777172, 0.02295635, 0.01978443, 0.02198051, 
    0.02249807, 0.02233846, 0.0217632, 0.02166845, 0.02273641, 0.02203057, 
    0.02044136, 0.01954997, 0.0187867, 0.01826475, 0.01809487, 0.01804989, 
    0.01884593, 0.01968232, 0.02029406, 0.02192587, 0.02340688, 0.02447821, 
    0.02557222, 0.02724179, 0.02747227, 0.02773753, 0.02813471, 0.02446154, 
    0.02414753, 0.02537229, 0.02483331, 0.02274387, 0.02079632, 0.02042781, 
    0.02170007, 0.02316828, 0.02243237, 0.02162332, 0.02185623, 0.02366399, 
    0.02629584, 0.02913469, 0.03117591, 0.03378513, 0.03736194, 0.04167927, 
    0.05277132, 0.07041078, 0.08518031, 0.08919548, 0.06725462, 0.03995897, 
    0.03365217, 0.03595219, 0.04206599, 0.06496944, 0.09696753, 0.1042428, 
    0.09851641, 0.09083464, 0.06892003, 0.04537698, 0.03707092, 0.04459516, 
    0.03816796, 0.03409632, 0.02832889, 0.02671107, 0.02450652, 0.02494191, 
    0.03013858, 0.0336157, 0.04169093, 0.05680138, 0.05748445, 0.04390349, 
    0.03158543, 0.02866537, 0.02939491, 0.03122962, 0.03192151, 0.03485339, 
    0.04126359, 0.04607936, 0.04884477, 0.05005344, 0.05046749, 0.04967235, 
    0.04934575, 0.04814013, 0.0479771, 0.04644149, 0.04390257, 0.04194877, 
    0.04025572, 0.03952574, 0.03839376, 0.03676733, 0.03778385, 0.0355649, 
    0.03499463, 0.03465552, 0.03247054, 0.0318761, 0.03069559, 0.02901737, 
    0.0275086, 0.02678503, 0.02427576, 0.02130729, 0.0199945, 0.01924322, 
    0.01855667, 0.01769974, 0.01728109, 0.01745064, 0.01752051, 0.01766785, 
    0.01848378, 0.01944344, 0.01827111, 0.01731056, 0.01790139, 0.01696019, 
    0.01684439, 0.01867269, 0.01877235, 0.01772859, 0.01807476, 0.01859893, 
    0.0186564, 0.01839924, 0.01863758, 0.01864603, 0.01744018, 0.01684268, 
    0.01614195, 0.01485893, 0.01411418, 0.01452143, 0.01523729, 0.01484755, 
    0.01559213, 0.01576696, 0.01547562, 0.0146574, 0.01482117, 0.01579634, 
    0.01544265, 0.01514752, 0.01488409, 0.01416514, 0.01440819, 0.01452968, 
    0.01292885, 0.01250047, 0.01303127, 0.01393875, 0.01479696, 0.01471797, 
    0.01506804, 0.01552029, 0.01519842, 0.01495381, 0.01535452, 0.01620945, 
    0.01731378, 0.01821378, 0.01915822, 0.01968677, 0.01983934, 0.0204213, 
    0.02102952, 0.02180574, 0.02244465, 0.02284802, 0.02293463, 0.02323283, 
    0.02448813, 0.02607032, 0.02614081, 0.02636035, 0.02714727, 0.02990422, 
    0.03432838, 0.03713189, 0.03906231, 0.04164972, 0.04702779, 0.05611863, 
    0.07522336, 0.1623715, 0.1809311, 0.1778388, 0.1529607, 0.1613728, 
    0.1172286, 0.1100199, 0.1152917, 0.1175998, 0.1146548, 0.1109925, 
    0.1029816, 0.09138937, 0.0886348, 0.08981584, 0.09307755, 0.1003316, 
    0.1021986, 0.1026041, 0.09784792, 0.07820296, 0.06309605, 0.0544925, 
    0.05136295, 0.04976251, 0.04329831, 0.03511009, 0.03072517, 0.0266341, 
    0.0239425, 0.02326826, 0.02438705, 0.02468398, 0.02519523, 0.02580579, 
    0.02568693, 0.02405693, 0.02183514, 0.02014718, 0.01854483, 0.01798542, 
    0.01748005, 0.01717737, 0.01708054, 0.0175447, 0.01770257, 0.0175636, 
    0.01755503, 0.01804996, 0.01899214, 0.01996569, 0.02163424, 0.02258541, 
    0.02327332, 0.02438207, 0.02597382, 0.02682121, 0.0273907, 0.0299175, 
    0.03321686, 0.03475304, 0.03628001, 0.03777347, 0.04068837, 0.04349675,
  0.04986641, 0.05250838, 0.0578535, 0.06325568, 0.06961139, 0.07571922, 
    0.0836582, 0.1214588, 0.1475727, 0.1349078, 0.1128942, 0.08370227, 
    0.07291131, 0.07031843, 0.06747958, 0.06702866, 0.06657697, 0.06654649, 
    0.06878867, 0.0761376, 0.08548865, 0.09672415, 0.1046744, 0.08914529, 
    0.07931412, 0.08542266, 0.1040794, 0.09937237, 0.0784643, 0.05909843, 
    0.04026609, 0.03847471, 0.03260865, 0.02794892, 0.02369966, 0.02334933, 
    0.02432884, 0.0255366, 0.02618611, 0.02623522, 0.02580932, 0.02422889, 
    0.02261715, 0.02087159, 0.01930872, 0.01847786, 0.01841001, 0.01896793, 
    0.01960123, 0.02006363, 0.02079988, 0.02264374, 0.02540141, 0.0261703, 
    0.02732331, 0.02879318, 0.03051184, 0.0321148, 0.03070435, 0.02922055, 
    0.02917485, 0.02902232, 0.02802, 0.02539031, 0.02380629, 0.02245311, 
    0.02224929, 0.02251834, 0.02202991, 0.02196065, 0.02205356, 0.02229265, 
    0.02349075, 0.026244, 0.02900013, 0.0337813, 0.03829216, 0.0457903, 
    0.05972428, 0.07402333, 0.08192742, 0.07627591, 0.05606763, 0.03682502, 
    0.03267089, 0.03534758, 0.04422747, 0.07499411, 0.1052454, 0.1230207, 
    0.1202913, 0.1096966, 0.08955316, 0.0596628, 0.03409068, 0.03096375, 
    0.03006517, 0.02806548, 0.02625393, 0.02593587, 0.02454463, 0.02659701, 
    0.03061546, 0.02742809, 0.02712231, 0.02950217, 0.03198462, 0.02757056, 
    0.0240135, 0.02463272, 0.02501951, 0.02648623, 0.02920306, 0.03365777, 
    0.04048881, 0.04418516, 0.04614387, 0.04796452, 0.04686943, 0.04542331, 
    0.04686569, 0.04655413, 0.04647433, 0.04683776, 0.04628544, 0.04382055, 
    0.04098234, 0.03984062, 0.03832961, 0.03691808, 0.03761068, 0.03714723, 
    0.03514845, 0.03408166, 0.03341963, 0.03303269, 0.03256755, 0.03054819, 
    0.02895771, 0.02831364, 0.02637961, 0.02340868, 0.02122947, 0.020465, 
    0.02085959, 0.02000273, 0.01948805, 0.01994014, 0.01920858, 0.01882501, 
    0.01903498, 0.01959538, 0.01994213, 0.01998699, 0.02091383, 0.02113875, 
    0.02025143, 0.01946691, 0.01876058, 0.01835893, 0.02006911, 0.02111643, 
    0.02035845, 0.02092565, 0.02202035, 0.02210996, 0.02088757, 0.02023904, 
    0.01951499, 0.02049798, 0.01929159, 0.01913104, 0.01930414, 0.01885005, 
    0.01864226, 0.01864866, 0.01731954, 0.0165975, 0.01699436, 0.01739988, 
    0.01622744, 0.01612895, 0.0156996, 0.01487574, 0.0154013, 0.01396028, 
    0.0136697, 0.01401149, 0.01383958, 0.01437888, 0.01566895, 0.01572165, 
    0.01515434, 0.01490873, 0.01463513, 0.0151213, 0.01628646, 0.01755709, 
    0.01842, 0.01939281, 0.02075398, 0.02154955, 0.02229657, 0.02346654, 
    0.02428624, 0.02598541, 0.02757626, 0.02794338, 0.02787872, 0.02863023, 
    0.03028448, 0.03137179, 0.03165954, 0.03265331, 0.03006847, 0.03297586, 
    0.04124347, 0.04451757, 0.04681375, 0.04960691, 0.05668755, 0.06345232, 
    0.0802638, 0.1412204, 0.1989398, 0.1368316, 0.1731685, 0.1618586, 
    0.1398883, 0.1125651, 0.1122657, 0.1157179, 0.1186229, 0.1233425, 
    0.1170517, 0.09325142, 0.08801771, 0.09429511, 0.09934294, 0.1058316, 
    0.1038702, 0.1024153, 0.09583161, 0.07564175, 0.06321659, 0.05523722, 
    0.05163421, 0.05386793, 0.04407772, 0.03833924, 0.03398187, 0.02981362, 
    0.02690833, 0.02610506, 0.02621646, 0.02600565, 0.02525775, 0.02454406, 
    0.02457901, 0.02379547, 0.02301147, 0.02287964, 0.02096757, 0.02002626, 
    0.01944628, 0.01897758, 0.0187995, 0.01929435, 0.01916927, 0.01902577, 
    0.01993129, 0.02099839, 0.02160992, 0.02226663, 0.02416926, 0.02510426, 
    0.02535264, 0.02696589, 0.02931349, 0.03135295, 0.03221764, 0.03298968, 
    0.03483218, 0.03744278, 0.03999544, 0.04254351, 0.0456947, 0.04793811,
  0.05229943, 0.05357234, 0.05819419, 0.06290362, 0.06827145, 0.07483136, 
    0.08609691, 0.1184235, 0.1309348, 0.1201339, 0.1088458, 0.0862074, 
    0.0734887, 0.06875373, 0.06557295, 0.06598467, 0.06580473, 0.06593693, 
    0.065853, 0.07097982, 0.07657026, 0.0807339, 0.08798672, 0.08101064, 
    0.06994822, 0.07706167, 0.08597628, 0.07899498, 0.07985171, 0.05007197, 
    0.0401657, 0.04496102, 0.04095409, 0.03504317, 0.02950704, 0.02560217, 
    0.02537163, 0.02691182, 0.02836986, 0.02920709, 0.02807115, 0.02668603, 
    0.02574917, 0.02404128, 0.02345044, 0.02281377, 0.02264042, 0.02280862, 
    0.02328165, 0.02342708, 0.02355334, 0.02455767, 0.02571525, 0.02606276, 
    0.02748615, 0.02846558, 0.03022716, 0.03230684, 0.03359711, 0.03404871, 
    0.03354619, 0.03090414, 0.02766794, 0.0248694, 0.02313944, 0.02200054, 
    0.02173867, 0.0222494, 0.02234067, 0.02182334, 0.02192638, 0.02165036, 
    0.02311962, 0.02601673, 0.0287889, 0.03337736, 0.03966104, 0.05528697, 
    0.06689974, 0.06609202, 0.07284351, 0.06130292, 0.04515888, 0.03502545, 
    0.0326853, 0.03334016, 0.03974072, 0.06185333, 0.08674236, 0.1175975, 
    0.1374136, 0.1247973, 0.1040512, 0.07430073, 0.04216116, 0.02944004, 
    0.02759772, 0.02546934, 0.02502669, 0.02638138, 0.02451529, 0.02591522, 
    0.0285333, 0.02452369, 0.02391472, 0.02382727, 0.02350976, 0.02250996, 
    0.02339371, 0.02518848, 0.02580319, 0.02671865, 0.02942351, 0.03385334, 
    0.03821384, 0.04215182, 0.04596968, 0.04880125, 0.04757516, 0.04627372, 
    0.04658451, 0.04805026, 0.04992319, 0.0515697, 0.05050924, 0.04721128, 
    0.04644659, 0.04666764, 0.04581078, 0.04444991, 0.04379598, 0.0403644, 
    0.03759375, 0.03961641, 0.03905955, 0.03850272, 0.03782439, 0.03554578, 
    0.03521479, 0.03404951, 0.03197655, 0.02871371, 0.02567578, 0.02466312, 
    0.02479726, 0.02413456, 0.02362987, 0.02335491, 0.0225041, 0.02129678, 
    0.02166044, 0.02273113, 0.02331744, 0.02485853, 0.0252875, 0.02474649, 
    0.02280181, 0.02122043, 0.02075997, 0.02065354, 0.02159375, 0.02233032, 
    0.022988, 0.02368848, 0.02354774, 0.02331976, 0.02383492, 0.02324636, 
    0.02301266, 0.02249191, 0.0222241, 0.02367183, 0.02351884, 0.02356571, 
    0.02356754, 0.0251518, 0.02460156, 0.02402717, 0.02341036, 0.02301211, 
    0.02159064, 0.02088142, 0.02010399, 0.02007314, 0.01938451, 0.01828404, 
    0.01728349, 0.01665409, 0.01646638, 0.01690709, 0.018192, 0.0192056, 
    0.01936119, 0.01920625, 0.01846243, 0.01874742, 0.01971387, 0.02100742, 
    0.02247307, 0.02393516, 0.02584661, 0.02731759, 0.02909592, 0.03040838, 
    0.03207435, 0.03488418, 0.03739217, 0.03974159, 0.04026159, 0.04133252, 
    0.04240828, 0.04295504, 0.04412303, 0.04557312, 0.04476215, 0.04940616, 
    0.05442471, 0.05600093, 0.05807179, 0.06254619, 0.07020036, 0.07574535, 
    0.08783913, 0.1157054, 0.2010647, 0.1755401, 0.1716934, 0.1621544, 
    0.1371242, 0.1243115, 0.1090929, 0.1125887, 0.1213785, 0.1336445, 
    0.1332411, 0.1050389, 0.08554439, 0.08832256, 0.0943388, 0.09827821, 
    0.09814787, 0.1014775, 0.09218153, 0.07246607, 0.06440153, 0.05953001, 
    0.06021297, 0.06056698, 0.04917613, 0.04259603, 0.03797711, 0.03496122, 
    0.03290766, 0.03265138, 0.03274468, 0.0319223, 0.03089156, 0.02979274, 
    0.02929613, 0.02849301, 0.02770463, 0.02785376, 0.02682653, 0.0257498, 
    0.02504284, 0.02415432, 0.02373921, 0.02508823, 0.0251289, 0.02421833, 
    0.02508114, 0.02597523, 0.02669863, 0.02755061, 0.02894411, 0.02988499, 
    0.03114431, 0.03327955, 0.0353252, 0.03727366, 0.03815947, 0.03878073, 
    0.0402206, 0.04156673, 0.04312441, 0.04561012, 0.04778424, 0.05075113,
  0.05179634, 0.05451632, 0.05708887, 0.06002564, 0.06493659, 0.07348485, 
    0.08615708, 0.108013, 0.1286253, 0.1141866, 0.1054193, 0.08962395, 
    0.07562353, 0.06885372, 0.06440905, 0.0628779, 0.06338336, 0.06413663, 
    0.06439903, 0.06756474, 0.0689643, 0.07001548, 0.0750255, 0.07154681, 
    0.06586843, 0.07386217, 0.06869753, 0.05825225, 0.0627449, 0.04160522, 
    0.03930461, 0.04873616, 0.0451591, 0.04054433, 0.03406364, 0.02907655, 
    0.02687808, 0.02792265, 0.03072871, 0.03233701, 0.03195917, 0.03138547, 
    0.03105298, 0.02916325, 0.02806829, 0.02681047, 0.02690853, 0.0279346, 
    0.02767514, 0.02733348, 0.02821402, 0.0281651, 0.02794807, 0.02788883, 
    0.02769732, 0.02923205, 0.03168881, 0.03309454, 0.03496552, 0.03729142, 
    0.03573319, 0.03160542, 0.02957223, 0.02816009, 0.02633095, 0.02535466, 
    0.02417951, 0.02363037, 0.02321573, 0.02199046, 0.02217423, 0.02309948, 
    0.02468709, 0.026126, 0.02913002, 0.03237063, 0.04546176, 0.06784577, 
    0.0720567, 0.07093643, 0.06817248, 0.05536269, 0.04674968, 0.03546417, 
    0.0317614, 0.03112123, 0.0336726, 0.03976326, 0.05241111, 0.08074851, 
    0.1156979, 0.1216318, 0.1071698, 0.08996606, 0.04836839, 0.02821214, 
    0.02431729, 0.0237328, 0.02461402, 0.02463896, 0.02413435, 0.02360757, 
    0.02460493, 0.02435243, 0.02389937, 0.02458107, 0.02371201, 0.02339938, 
    0.02431253, 0.02615457, 0.02745729, 0.02837377, 0.03101077, 0.03533801, 
    0.03888926, 0.04028147, 0.04416792, 0.04731575, 0.04815015, 0.0484316, 
    0.04871658, 0.05014458, 0.05168357, 0.05225987, 0.05145884, 0.05037756, 
    0.05117728, 0.05186155, 0.05142887, 0.05117663, 0.04944124, 0.04735002, 
    0.04648421, 0.04766786, 0.04599241, 0.04418365, 0.0426169, 0.04212745, 
    0.04284725, 0.04263914, 0.04109502, 0.03815038, 0.0351375, 0.0333699, 
    0.03198151, 0.03146535, 0.03053496, 0.02911511, 0.02786765, 0.02724672, 
    0.02808828, 0.02901429, 0.02938939, 0.03096159, 0.03114763, 0.02987807, 
    0.02909971, 0.02871905, 0.02856501, 0.02765215, 0.02664495, 0.02715771, 
    0.02823512, 0.0282695, 0.02735601, 0.0270615, 0.0275594, 0.0287574, 
    0.02900844, 0.02809591, 0.02752163, 0.02987361, 0.03008633, 0.03119655, 
    0.03324803, 0.03488878, 0.0349169, 0.03387226, 0.03316629, 0.03193708, 
    0.03028104, 0.02937988, 0.02872566, 0.02833983, 0.0276145, 0.0263796, 
    0.02544067, 0.02490757, 0.02490543, 0.02550521, 0.02678556, 0.02843541, 
    0.02873779, 0.02837603, 0.02756545, 0.02781266, 0.02865536, 0.02998594, 
    0.03157002, 0.03332013, 0.03586826, 0.03860395, 0.04074928, 0.04270023, 
    0.04561539, 0.04973901, 0.05298469, 0.0566787, 0.05787273, 0.05923574, 
    0.05957647, 0.06041395, 0.0627175, 0.06484255, 0.06505142, 0.06746313, 
    0.06954252, 0.07224782, 0.07722738, 0.08120805, 0.08482239, 0.09051513, 
    0.09882186, 0.1093226, 0.1543367, 0.2251481, 0.1696371, 0.1392592, 
    0.1278817, 0.1231363, 0.1121999, 0.1090877, 0.1237253, 0.1432736, 
    0.1532738, 0.1228534, 0.08058333, 0.08119396, 0.08517177, 0.08769926, 
    0.08816963, 0.09641781, 0.08604, 0.07192607, 0.063842, 0.06062502, 
    0.06377136, 0.05590926, 0.04859745, 0.04389085, 0.04166502, 0.0402115, 
    0.03997936, 0.04014896, 0.04058409, 0.04020153, 0.03851191, 0.03659303, 
    0.03584037, 0.03535854, 0.03471472, 0.03490839, 0.03475742, 0.03430277, 
    0.03311156, 0.03200661, 0.03173422, 0.03176932, 0.03150924, 0.03163839, 
    0.03353735, 0.03586274, 0.03750089, 0.03739775, 0.03852263, 0.03940742, 
    0.03930281, 0.0406975, 0.04197417, 0.04351396, 0.04404034, 0.04443109, 
    0.04439978, 0.04460325, 0.0457202, 0.04736349, 0.04888625, 0.05019845,
  0.04883888, 0.05207846, 0.0557684, 0.05899125, 0.06564034, 0.0774603, 
    0.09343915, 0.1128652, 0.1404617, 0.1116451, 0.09705063, 0.084846, 
    0.07715022, 0.06871299, 0.06298815, 0.06253467, 0.06129386, 0.06088484, 
    0.06213624, 0.06354686, 0.06298351, 0.06215923, 0.06596717, 0.06725674, 
    0.06589434, 0.07712184, 0.06232239, 0.05449207, 0.06130175, 0.04722662, 
    0.04390738, 0.0505407, 0.04854626, 0.04450474, 0.0382524, 0.03119005, 
    0.02783287, 0.02699283, 0.03040961, 0.03271791, 0.03347649, 0.03429069, 
    0.0345801, 0.03318458, 0.03036327, 0.02897567, 0.02879186, 0.02870567, 
    0.02790796, 0.02767961, 0.02928001, 0.02989681, 0.03032114, 0.03067068, 
    0.0302767, 0.03134691, 0.03277866, 0.03262723, 0.03286873, 0.03489966, 
    0.03425456, 0.03276259, 0.0337799, 0.03445676, 0.03024925, 0.02932792, 
    0.02776497, 0.02672202, 0.02652298, 0.02514144, 0.02402805, 0.02421146, 
    0.02467509, 0.02601925, 0.02906999, 0.03532917, 0.05477495, 0.06145175, 
    0.0697154, 0.06325381, 0.06436722, 0.05952332, 0.05349459, 0.03737344, 
    0.0316072, 0.03123541, 0.03281618, 0.03458112, 0.03762868, 0.04722734, 
    0.07387168, 0.1003562, 0.09717338, 0.09307718, 0.050696, 0.02832583, 
    0.02297624, 0.02208195, 0.02328471, 0.02484998, 0.02648141, 0.02488117, 
    0.02483638, 0.02504472, 0.02588945, 0.02732346, 0.02515432, 0.02471932, 
    0.02607164, 0.02793185, 0.02986871, 0.0312715, 0.03423305, 0.03739439, 
    0.03971124, 0.0407814, 0.04613769, 0.0492657, 0.05060571, 0.05165395, 
    0.05227783, 0.05382256, 0.05507325, 0.05351476, 0.05261897, 0.05337119, 
    0.05477208, 0.05469283, 0.05406009, 0.05389338, 0.05342441, 0.05325766, 
    0.05308734, 0.05442834, 0.05307288, 0.05130561, 0.05230546, 0.05217601, 
    0.05157642, 0.0512783, 0.0518851, 0.05042449, 0.04807186, 0.04689195, 
    0.04450653, 0.0418048, 0.03971557, 0.03883458, 0.03787918, 0.03745075, 
    0.03741636, 0.03796552, 0.03805178, 0.03890582, 0.03875898, 0.03804915, 
    0.03822937, 0.03810505, 0.03761837, 0.03600506, 0.03521143, 0.03543708, 
    0.03607991, 0.0365377, 0.0364548, 0.03711151, 0.03822165, 0.04041172, 
    0.04097278, 0.0400704, 0.04013021, 0.04331563, 0.04650907, 0.04877845, 
    0.05156443, 0.05160406, 0.05063362, 0.04922061, 0.0483287, 0.04684845, 
    0.04559768, 0.04504215, 0.04439674, 0.04438442, 0.04259121, 0.04051853, 
    0.03953658, 0.03893713, 0.03862131, 0.039554, 0.04086574, 0.0426972, 
    0.04380123, 0.04368706, 0.04311957, 0.04323966, 0.04413147, 0.04598963, 
    0.04725104, 0.04924154, 0.05193194, 0.05452498, 0.05827531, 0.06199812, 
    0.0662024, 0.07002578, 0.07206206, 0.07653134, 0.07773007, 0.07900678, 
    0.08208504, 0.08524244, 0.08758701, 0.08839321, 0.08762951, 0.08715571, 
    0.08772764, 0.09001775, 0.09340809, 0.09451589, 0.09529917, 0.09777389, 
    0.1023369, 0.1099159, 0.1228478, 0.2071744, 0.1782843, 0.1280806, 
    0.126758, 0.1145395, 0.1167193, 0.1075257, 0.1243438, 0.1483686, 
    0.1589983, 0.1190686, 0.08326109, 0.08435445, 0.07808921, 0.06791012, 
    0.06756666, 0.07929652, 0.07422719, 0.06724503, 0.05695672, 0.05779675, 
    0.06252621, 0.04967194, 0.04348904, 0.04175106, 0.04231432, 0.0428918, 
    0.04441659, 0.04543127, 0.04586346, 0.04630256, 0.0448552, 0.04317228, 
    0.04310319, 0.04308272, 0.04269306, 0.04341133, 0.04461282, 0.04531863, 
    0.04456108, 0.04373526, 0.04315275, 0.04223269, 0.04212509, 0.04232476, 
    0.04367933, 0.0451284, 0.04650279, 0.0470052, 0.04910181, 0.05027647, 
    0.04910763, 0.05059471, 0.05282351, 0.05300889, 0.05318496, 0.05237241, 
    0.04968585, 0.04613129, 0.0437906, 0.04404783, 0.04505183, 0.04622821,
  0.04589806, 0.04834366, 0.05292371, 0.05917929, 0.07104979, 0.08434532, 
    0.1036541, 0.1281839, 0.1312312, 0.1147722, 0.09885063, 0.08425944, 
    0.07742715, 0.06784906, 0.06163255, 0.0613455, 0.06025069, 0.05910351, 
    0.05998555, 0.05900616, 0.05861693, 0.05725485, 0.05817165, 0.05892462, 
    0.06239516, 0.07295182, 0.06492011, 0.06420512, 0.07677308, 0.06588352, 
    0.05202347, 0.05293332, 0.04825455, 0.04706685, 0.04148302, 0.0333258, 
    0.03071754, 0.02467944, 0.02611362, 0.03070828, 0.03226675, 0.03352658, 
    0.03384781, 0.03334852, 0.031458, 0.02978773, 0.0291572, 0.02931046, 
    0.02857089, 0.02812643, 0.02962439, 0.03056234, 0.03110812, 0.03257262, 
    0.03308641, 0.03228596, 0.03171023, 0.03157042, 0.0317435, 0.03277948, 
    0.03252235, 0.03229588, 0.03519554, 0.03665205, 0.03453123, 0.03160849, 
    0.02855498, 0.02756751, 0.0280889, 0.02685898, 0.0255363, 0.0250191, 
    0.02590718, 0.02627223, 0.02755795, 0.03415854, 0.04742798, 0.06755874, 
    0.05725481, 0.05554872, 0.05873578, 0.06067783, 0.05763929, 0.03958735, 
    0.03343518, 0.03266213, 0.03282337, 0.0320847, 0.03168993, 0.0342777, 
    0.04488577, 0.06878589, 0.07845326, 0.07719603, 0.05206931, 0.02960412, 
    0.02271289, 0.0221017, 0.0246885, 0.02868749, 0.03071656, 0.0291551, 
    0.02653991, 0.02642395, 0.02740264, 0.02874096, 0.02769181, 0.02794419, 
    0.02982902, 0.03098221, 0.03262771, 0.03486636, 0.03855042, 0.04168312, 
    0.04156403, 0.0429176, 0.04772613, 0.05056026, 0.05164365, 0.05185647, 
    0.05380339, 0.05696391, 0.05861051, 0.05828356, 0.05793695, 0.05902091, 
    0.05865157, 0.05864482, 0.05862342, 0.05791178, 0.05808692, 0.05742078, 
    0.05671876, 0.05823026, 0.05911991, 0.05893645, 0.05954497, 0.05921469, 
    0.05721171, 0.05737682, 0.05836525, 0.05800781, 0.05667484, 0.05663272, 
    0.05656931, 0.05483519, 0.05372664, 0.05235979, 0.05262083, 0.05239738, 
    0.05210334, 0.05284294, 0.05187751, 0.05055766, 0.0489516, 0.04757382, 
    0.04735276, 0.04782788, 0.04725866, 0.04625741, 0.04666347, 0.04825916, 
    0.04939736, 0.05037833, 0.0503078, 0.05117651, 0.05289491, 0.05534542, 
    0.05563162, 0.05675091, 0.0593378, 0.06323208, 0.06573076, 0.06648124, 
    0.06684333, 0.06731362, 0.06886741, 0.06854027, 0.06742227, 0.06676183, 
    0.06585046, 0.06528906, 0.06596967, 0.06634127, 0.06410767, 0.06116844, 
    0.05892134, 0.0576822, 0.05729831, 0.05815331, 0.05864356, 0.05987791, 
    0.06179534, 0.06320518, 0.06339034, 0.06389747, 0.06495681, 0.06635178, 
    0.06737942, 0.06994507, 0.07112075, 0.07241466, 0.07703286, 0.08283644, 
    0.08672891, 0.09004501, 0.09375018, 0.09844629, 0.09951411, 0.102338, 
    0.10826, 0.1114455, 0.1106761, 0.1058263, 0.1005445, 0.09812774, 
    0.09971543, 0.1017688, 0.1011941, 0.09647854, 0.09245783, 0.09518746, 
    0.09972955, 0.1054489, 0.1164774, 0.196929, 0.2321772, 0.1437634, 
    0.1300364, 0.1134284, 0.105139, 0.110228, 0.1169645, 0.1362031, 
    0.1308693, 0.0987137, 0.09161043, 0.09926193, 0.06929956, 0.04827131, 
    0.05213542, 0.06041135, 0.05590325, 0.05088041, 0.04701529, 0.051068, 
    0.04938715, 0.04221347, 0.04020627, 0.04091909, 0.04296901, 0.04454561, 
    0.04656802, 0.04816124, 0.04955246, 0.05048264, 0.04949328, 0.04777836, 
    0.04790648, 0.04872162, 0.04971419, 0.05034576, 0.05065368, 0.05206226, 
    0.05194512, 0.05131026, 0.0505615, 0.04936946, 0.04914546, 0.04980595, 
    0.04980806, 0.05175494, 0.05335218, 0.05305861, 0.0548066, 0.05601532, 
    0.05653772, 0.06032214, 0.06458553, 0.06657273, 0.06689629, 0.06431508, 
    0.05661671, 0.04942723, 0.04672094, 0.04545285, 0.0441326, 0.04445795,
  0.0457286, 0.0478846, 0.05155115, 0.05987031, 0.07853939, 0.09286968, 
    0.112978, 0.122041, 0.1034327, 0.09757135, 0.09835058, 0.08307677, 
    0.07197738, 0.06475214, 0.05894481, 0.05711766, 0.05768393, 0.05771187, 
    0.05603747, 0.05494858, 0.05456998, 0.05148897, 0.0523911, 0.05332775, 
    0.0581013, 0.06662201, 0.06972522, 0.08215453, 0.09602542, 0.0955858, 
    0.07598194, 0.0701125, 0.0542199, 0.04977514, 0.04481956, 0.04091912, 
    0.0355735, 0.02697895, 0.02411562, 0.02833537, 0.03045692, 0.03213936, 
    0.03298115, 0.0334084, 0.03330198, 0.03226626, 0.03063435, 0.02967102, 
    0.02908302, 0.02866756, 0.02833801, 0.02799061, 0.02801911, 0.02900825, 
    0.02959566, 0.03014884, 0.03015356, 0.03066458, 0.03066236, 0.03209119, 
    0.03215068, 0.03150955, 0.03503985, 0.0378005, 0.03333072, 0.03220377, 
    0.02972521, 0.02677956, 0.02706519, 0.02710952, 0.02655797, 0.02668952, 
    0.02789797, 0.02739757, 0.02668661, 0.02909667, 0.03149635, 0.03873442, 
    0.04261219, 0.04103664, 0.04897959, 0.05461355, 0.05053348, 0.03648377, 
    0.03315528, 0.03275239, 0.03243277, 0.03171181, 0.03005778, 0.03064525, 
    0.03360368, 0.04342002, 0.0548628, 0.06371824, 0.05088899, 0.0312306, 
    0.02463548, 0.02580291, 0.03076884, 0.03731127, 0.03963207, 0.03905732, 
    0.03323049, 0.03110332, 0.03133984, 0.03227173, 0.0328095, 0.03250253, 
    0.03279964, 0.0335844, 0.0351812, 0.03724592, 0.03986079, 0.04245454, 
    0.04281548, 0.04518891, 0.04945318, 0.05133661, 0.05112813, 0.04922695, 
    0.05180546, 0.05512983, 0.05686945, 0.05831607, 0.05941842, 0.05980465, 
    0.05921773, 0.05874623, 0.05964778, 0.05848455, 0.05728613, 0.05712925, 
    0.05614773, 0.05785547, 0.05965118, 0.06014472, 0.06049122, 0.0608254, 
    0.0605162, 0.06117262, 0.06139848, 0.06211004, 0.06207179, 0.06350145, 
    0.06503243, 0.06538725, 0.06528068, 0.06480274, 0.06268547, 0.06249857, 
    0.06401477, 0.0648397, 0.06370712, 0.06237927, 0.06108204, 0.05916771, 
    0.05969063, 0.06053837, 0.06004527, 0.05926127, 0.06054537, 0.06306778, 
    0.06486022, 0.06560118, 0.0661473, 0.06689603, 0.06855097, 0.07040298, 
    0.07167114, 0.07494978, 0.07818179, 0.08096636, 0.08186241, 0.08109967, 
    0.08072784, 0.08001984, 0.08099347, 0.08320327, 0.08480702, 0.08590253, 
    0.08477212, 0.08460677, 0.08675283, 0.08435401, 0.08145466, 0.07851275, 
    0.07569309, 0.07414995, 0.07378177, 0.07442726, 0.07545555, 0.07839615, 
    0.07956687, 0.08085965, 0.08118448, 0.08146254, 0.08283637, 0.08578791, 
    0.08923754, 0.0910614, 0.09029373, 0.08966035, 0.09338712, 0.09919361, 
    0.1027901, 0.1068233, 0.1117671, 0.1170486, 0.1183539, 0.1197786, 
    0.1227431, 0.1207513, 0.1140594, 0.1063389, 0.1000628, 0.09839185, 
    0.1005419, 0.1004474, 0.09674043, 0.08798659, 0.08419739, 0.08621107, 
    0.0879923, 0.09400932, 0.1115899, 0.1870288, 0.2298715, 0.1547712, 
    0.1386014, 0.1071124, 0.09156919, 0.1038265, 0.1067417, 0.1134217, 
    0.1002757, 0.08474399, 0.09993, 0.09515645, 0.06564442, 0.06707708, 
    0.05448309, 0.0454823, 0.03800407, 0.03645157, 0.03729429, 0.03865641, 
    0.03877585, 0.03898203, 0.04073184, 0.0438589, 0.04718714, 0.04898629, 
    0.0502359, 0.05081332, 0.05049293, 0.05003227, 0.04936592, 0.04855116, 
    0.04899113, 0.04993936, 0.0520372, 0.05276117, 0.0520832, 0.0523281, 
    0.05240058, 0.05169404, 0.05143316, 0.05219736, 0.05142377, 0.05265403, 
    0.05385877, 0.05608376, 0.0576265, 0.05810763, 0.05908216, 0.06180924, 
    0.06545754, 0.07064918, 0.07580774, 0.08045565, 0.08730312, 0.07979757, 
    0.0670667, 0.06050773, 0.05899139, 0.05950329, 0.05561388, 0.04908825,
  0.05243298, 0.05190288, 0.05825469, 0.0668688, 0.07729503, 0.08165443, 
    0.09571967, 0.0991933, 0.08175094, 0.07994569, 0.0815462, 0.07188552, 
    0.06112352, 0.0584593, 0.05512154, 0.05165155, 0.05314015, 0.05390555, 
    0.05339517, 0.05325707, 0.05087776, 0.04795932, 0.04874486, 0.05071012, 
    0.05494633, 0.0609672, 0.07168358, 0.09660362, 0.09958061, 0.1155266, 
    0.09289731, 0.08667054, 0.05922179, 0.05700114, 0.05247873, 0.04904858, 
    0.0425964, 0.03397981, 0.02704951, 0.02639638, 0.02792053, 0.02896164, 
    0.03002032, 0.03075467, 0.03188932, 0.03141463, 0.03013936, 0.02888803, 
    0.02837475, 0.02810218, 0.02723541, 0.02710635, 0.02673952, 0.02669797, 
    0.02666045, 0.02688713, 0.02747582, 0.02830817, 0.02870806, 0.0294848, 
    0.02978224, 0.03028359, 0.03427413, 0.03711968, 0.05006626, 0.03675403, 
    0.03369838, 0.02753047, 0.02665354, 0.0272968, 0.02808106, 0.02808431, 
    0.02807883, 0.02818427, 0.0269712, 0.02812876, 0.03074709, 0.03326106, 
    0.0331471, 0.0348983, 0.04010919, 0.03966983, 0.03876363, 0.03350795, 
    0.03321093, 0.03419041, 0.03529706, 0.0354298, 0.03310524, 0.03212805, 
    0.03249224, 0.03608013, 0.04135934, 0.04743697, 0.04107318, 0.03142054, 
    0.02980699, 0.03527032, 0.04586899, 0.06222319, 0.05358434, 0.04923726, 
    0.04189903, 0.03877736, 0.0379241, 0.03814414, 0.03798731, 0.03621383, 
    0.0360469, 0.03734984, 0.03932207, 0.03836565, 0.03937757, 0.04151199, 
    0.04339442, 0.04511584, 0.04818676, 0.0501184, 0.04932878, 0.04868222, 
    0.05129987, 0.05320757, 0.05508092, 0.05874679, 0.0595977, 0.05844279, 
    0.0585673, 0.05747877, 0.05597914, 0.05506203, 0.05366465, 0.05194024, 
    0.05179242, 0.05357135, 0.05593162, 0.05684721, 0.05806283, 0.05941026, 
    0.05923298, 0.0603048, 0.0616301, 0.06193368, 0.06277113, 0.06495329, 
    0.06544695, 0.0653372, 0.06590417, 0.06578053, 0.06616698, 0.0670898, 
    0.06650943, 0.06742966, 0.06806649, 0.06919316, 0.06947188, 0.06826963, 
    0.06865086, 0.06873808, 0.06823321, 0.06913048, 0.07159768, 0.07325273, 
    0.07509277, 0.07607956, 0.07863615, 0.08105278, 0.08218025, 0.08396509, 
    0.08612701, 0.0881194, 0.08897891, 0.08912562, 0.09114033, 0.09053434, 
    0.08951386, 0.08791916, 0.08711606, 0.08864114, 0.09130885, 0.09385484, 
    0.09464271, 0.09559885, 0.0949965, 0.09227613, 0.09014239, 0.08796883, 
    0.08524537, 0.08347917, 0.08183887, 0.08114079, 0.08185182, 0.08477782, 
    0.08628175, 0.08743861, 0.09003703, 0.0922745, 0.09459753, 0.09692322, 
    0.1028318, 0.1050522, 0.1022673, 0.10016, 0.1035568, 0.1075555, 
    0.1098181, 0.1120495, 0.1158748, 0.1203068, 0.1194732, 0.1190751, 
    0.117741, 0.1095231, 0.1004412, 0.09476339, 0.09115983, 0.0891711, 
    0.08771286, 0.0832878, 0.07958499, 0.07605355, 0.07396518, 0.07882128, 
    0.08335813, 0.08548491, 0.100047, 0.1551971, 0.1733794, 0.1461696, 
    0.1544292, 0.102448, 0.08154808, 0.08677424, 0.09392811, 0.08746134, 
    0.07987249, 0.0766984, 0.07436937, 0.05899989, 0.048177, 0.04783915, 
    0.04293912, 0.03306518, 0.02436708, 0.02569251, 0.0293389, 0.03341536, 
    0.03697374, 0.03816646, 0.04084089, 0.04415267, 0.0461293, 0.04752768, 
    0.04914623, 0.04842831, 0.04739136, 0.04633022, 0.04606566, 0.04670718, 
    0.04692335, 0.04731394, 0.04963287, 0.05117201, 0.05173125, 0.05237664, 
    0.05351228, 0.05284422, 0.05153544, 0.0529456, 0.05463774, 0.05662683, 
    0.05815332, 0.06085093, 0.06285218, 0.06458426, 0.06516053, 0.06792141, 
    0.07273137, 0.07962786, 0.08573261, 0.09811158, 0.0929506, 0.07969087, 
    0.06701776, 0.06190515, 0.06222123, 0.06280194, 0.05784311, 0.05367771,
  0.05608489, 0.06035349, 0.06983824, 0.0752639, 0.07158773, 0.07022344, 
    0.07633506, 0.07681914, 0.07034085, 0.06077309, 0.06052647, 0.05724704, 
    0.05161966, 0.05165395, 0.04831569, 0.0451626, 0.04818129, 0.0498985, 
    0.04839369, 0.04747771, 0.04574471, 0.04481749, 0.04471932, 0.04625067, 
    0.05032805, 0.05618039, 0.07285128, 0.1086147, 0.09979778, 0.1064707, 
    0.09111166, 0.07165086, 0.06068331, 0.06412558, 0.05457838, 0.04445785, 
    0.04262874, 0.03783755, 0.02762993, 0.02351683, 0.02579901, 0.02500321, 
    0.02521937, 0.02583379, 0.02699902, 0.02765316, 0.0275341, 0.02709636, 
    0.02760663, 0.0276922, 0.02794196, 0.02755237, 0.02637006, 0.02616483, 
    0.02630238, 0.02704532, 0.02783459, 0.02824612, 0.0281203, 0.02868137, 
    0.02977401, 0.02993452, 0.03349351, 0.03599915, 0.0460257, 0.03967113, 
    0.03581498, 0.02828522, 0.02669952, 0.02786978, 0.02958566, 0.02988895, 
    0.02857457, 0.02837807, 0.02823576, 0.02903237, 0.02946426, 0.02945283, 
    0.03321895, 0.03682951, 0.03706574, 0.03550012, 0.03415871, 0.03459586, 
    0.03592787, 0.03768745, 0.0401323, 0.04039932, 0.03883645, 0.03733677, 
    0.03636063, 0.0359125, 0.03517168, 0.03782834, 0.03687936, 0.03533482, 
    0.03567724, 0.0426144, 0.05813991, 0.07183065, 0.07188759, 0.05888205, 
    0.05045001, 0.04629659, 0.04419125, 0.04252151, 0.04075627, 0.03855356, 
    0.0378857, 0.03942829, 0.04014604, 0.03978512, 0.04003176, 0.04147349, 
    0.04354741, 0.0453558, 0.04817552, 0.05035514, 0.04856683, 0.04981893, 
    0.05264092, 0.05435606, 0.05620144, 0.05908739, 0.05965048, 0.05755793, 
    0.05571971, 0.05329654, 0.05067739, 0.05000177, 0.04964172, 0.04709496, 
    0.04677539, 0.04886495, 0.05117758, 0.05287857, 0.05454692, 0.05530584, 
    0.05528899, 0.05624204, 0.05588252, 0.05494918, 0.05631785, 0.05757856, 
    0.05718395, 0.05778811, 0.06074443, 0.06399892, 0.06659526, 0.06686927, 
    0.06610674, 0.0652755, 0.06537993, 0.06632292, 0.0664052, 0.06540778, 
    0.06505962, 0.06567322, 0.06703302, 0.0692331, 0.07211971, 0.07394871, 
    0.07613424, 0.07843073, 0.08059781, 0.08421196, 0.08588891, 0.08588605, 
    0.08666491, 0.08792265, 0.08847824, 0.09032013, 0.09343155, 0.09261366, 
    0.09229975, 0.09044863, 0.08830366, 0.08852063, 0.09035902, 0.09126785, 
    0.09133448, 0.09116547, 0.08962554, 0.08767184, 0.08462778, 0.08373934, 
    0.08232847, 0.08143999, 0.08075476, 0.07997023, 0.08072858, 0.08144248, 
    0.0810405, 0.082376, 0.08548304, 0.08992379, 0.09336365, 0.09386885, 
    0.09678318, 0.09912988, 0.09667598, 0.09685497, 0.09985622, 0.1020139, 
    0.1016094, 0.1017895, 0.1020401, 0.1033304, 0.1005784, 0.09630528, 
    0.09367199, 0.08686554, 0.07895774, 0.07551445, 0.07381663, 0.07044635, 
    0.06622453, 0.06240666, 0.06160411, 0.06389514, 0.07772423, 0.081821, 
    0.07199226, 0.07025368, 0.07769078, 0.1038164, 0.114978, 0.1158042, 
    0.1263518, 0.08495602, 0.05925608, 0.06265133, 0.0688597, 0.06859561, 
    0.06162036, 0.05763126, 0.04791713, 0.0327499, 0.03041994, 0.03477615, 
    0.03176697, 0.02437766, 0.02279621, 0.02562189, 0.02854234, 0.03121905, 
    0.03371095, 0.03572441, 0.03800306, 0.04063363, 0.04137972, 0.04243767, 
    0.04377886, 0.04300224, 0.041362, 0.04057363, 0.04081821, 0.04197293, 
    0.04203008, 0.04336404, 0.04655787, 0.04980263, 0.0516493, 0.05272131, 
    0.05433715, 0.05558387, 0.0535075, 0.05214072, 0.05345461, 0.05586325, 
    0.05739329, 0.05998403, 0.06195508, 0.06508944, 0.06855445, 0.07267126, 
    0.07998131, 0.09060573, 0.1012063, 0.1014438, 0.08749818, 0.0714274, 
    0.06243314, 0.05885784, 0.05945316, 0.05762782, 0.05303568, 0.0556884,
  0.05345307, 0.05534841, 0.06189281, 0.05813013, 0.05675507, 0.06503336, 
    0.06978922, 0.06420311, 0.05879938, 0.04805994, 0.04579399, 0.04464504, 
    0.04287574, 0.0421496, 0.03911906, 0.03802187, 0.04084135, 0.041625, 
    0.03897763, 0.03760995, 0.03764689, 0.03917056, 0.03975299, 0.04076402, 
    0.04483338, 0.0501019, 0.0679144, 0.09972058, 0.09845768, 0.1008841, 
    0.07762234, 0.06311834, 0.05698079, 0.06174193, 0.04660654, 0.0319481, 
    0.03821448, 0.03802304, 0.02706929, 0.02046681, 0.02291455, 0.0236023, 
    0.02222753, 0.02271531, 0.02409831, 0.02515203, 0.02573505, 0.026706, 
    0.02793199, 0.02811064, 0.02823283, 0.02772011, 0.02716054, 0.0270295, 
    0.02721304, 0.02873967, 0.02940103, 0.02946366, 0.02937698, 0.0312909, 
    0.03440816, 0.0352261, 0.03724235, 0.03756274, 0.03815816, 0.03775954, 
    0.03485266, 0.03006556, 0.02923672, 0.02991281, 0.03155061, 0.03229623, 
    0.03150147, 0.03097673, 0.03140908, 0.03128309, 0.03129585, 0.03338944, 
    0.03725153, 0.04056835, 0.03938277, 0.03729727, 0.03815563, 0.04072917, 
    0.04044873, 0.04129932, 0.04437134, 0.04595092, 0.04536551, 0.04416436, 
    0.04230801, 0.03876592, 0.03647415, 0.03881689, 0.04030626, 0.04065445, 
    0.04082426, 0.0444384, 0.05266613, 0.06005393, 0.07413203, 0.05924625, 
    0.05068444, 0.04581438, 0.04381552, 0.0432342, 0.04067446, 0.0386619, 
    0.03742732, 0.03804829, 0.03849375, 0.03880434, 0.03976521, 0.04017506, 
    0.04151643, 0.04357323, 0.04727805, 0.04921268, 0.04799205, 0.04915478, 
    0.0506803, 0.05266103, 0.05418409, 0.05593357, 0.05685601, 0.05485952, 
    0.05136911, 0.0488169, 0.04534718, 0.04513217, 0.04541991, 0.04404333, 
    0.04512629, 0.04743305, 0.04815789, 0.04854067, 0.04941194, 0.04921339, 
    0.04977734, 0.05032238, 0.04899475, 0.04796146, 0.04845577, 0.04791865, 
    0.04751949, 0.04858061, 0.05145791, 0.05411108, 0.05535315, 0.05570206, 
    0.05555427, 0.05476114, 0.0542864, 0.0544767, 0.05534462, 0.05572141, 
    0.05605181, 0.05745432, 0.05940767, 0.06112962, 0.06419643, 0.06741823, 
    0.07013489, 0.07325635, 0.07394109, 0.07587638, 0.07656052, 0.07605117, 
    0.07771453, 0.0791974, 0.08167154, 0.0843389, 0.08551206, 0.0838214, 
    0.08445282, 0.08327845, 0.0828858, 0.0831115, 0.08388694, 0.08384174, 
    0.08193242, 0.07981985, 0.07754851, 0.07701109, 0.07360408, 0.0721053, 
    0.07187159, 0.07194107, 0.07263621, 0.07230937, 0.07351188, 0.0729524, 
    0.07200362, 0.07287546, 0.07541426, 0.07860371, 0.08050186, 0.07896488, 
    0.07895987, 0.0793565, 0.07798538, 0.07997005, 0.08194105, 0.0827266, 
    0.08121189, 0.08040956, 0.07897906, 0.07900673, 0.07761682, 0.07281344, 
    0.07090311, 0.06743492, 0.06178792, 0.0580017, 0.05661423, 0.05312266, 
    0.05037297, 0.04912028, 0.05127877, 0.06386884, 0.07413544, 0.06856319, 
    0.0594278, 0.06077348, 0.05249545, 0.05704942, 0.0596463, 0.06932046, 
    0.07862999, 0.06018959, 0.05308184, 0.0498653, 0.04994573, 0.05523776, 
    0.04669126, 0.04395777, 0.03363037, 0.02474075, 0.02735636, 0.02684261, 
    0.02234831, 0.021146, 0.0215788, 0.02408512, 0.02648213, 0.02805969, 
    0.03014752, 0.03200868, 0.03380541, 0.03477873, 0.03515255, 0.03601885, 
    0.03634506, 0.03489209, 0.03388325, 0.03532391, 0.03596908, 0.03649924, 
    0.03749718, 0.03936746, 0.042439, 0.04501104, 0.04676861, 0.04797165, 
    0.04938341, 0.05118472, 0.05050617, 0.04894041, 0.04869412, 0.04948731, 
    0.05052535, 0.05263443, 0.05560961, 0.06076206, 0.06651087, 0.072826, 
    0.08337981, 0.09584143, 0.1013424, 0.09045696, 0.07071152, 0.05925229, 
    0.05560481, 0.05447879, 0.0534962, 0.04930124, 0.04853484, 0.05358144,
  0.04602036, 0.04658765, 0.04700706, 0.04709936, 0.05453397, 0.0657941, 
    0.06287082, 0.04787971, 0.04286979, 0.03910012, 0.0360431, 0.03325357, 
    0.03330067, 0.03361613, 0.03233024, 0.03102532, 0.03199643, 0.03330225, 
    0.0316394, 0.03011093, 0.03052714, 0.03171076, 0.03393304, 0.03610464, 
    0.03995963, 0.04375389, 0.05730303, 0.07636759, 0.09381768, 0.1026837, 
    0.07937243, 0.06679252, 0.05715704, 0.0493504, 0.03939172, 0.03818316, 
    0.03767071, 0.03351253, 0.02706805, 0.01943015, 0.02137843, 0.02278769, 
    0.02064488, 0.02109626, 0.02252604, 0.02391525, 0.02468729, 0.02654913, 
    0.02862076, 0.02900708, 0.02920057, 0.02938818, 0.02893821, 0.02888948, 
    0.0295775, 0.03008535, 0.03082765, 0.03158888, 0.03231109, 0.03706008, 
    0.04323716, 0.04833623, 0.04699172, 0.0412245, 0.03405977, 0.03488784, 
    0.03437638, 0.03260232, 0.03233042, 0.03255163, 0.03301643, 0.03322633, 
    0.03404009, 0.03394748, 0.03358162, 0.03281315, 0.03255188, 0.03596738, 
    0.04021516, 0.04329084, 0.04399862, 0.04302711, 0.04623872, 0.04974987, 
    0.05156622, 0.04763511, 0.04790213, 0.04924455, 0.04857693, 0.04864065, 
    0.04810505, 0.0465131, 0.04451843, 0.04454938, 0.04690765, 0.04310122, 
    0.04411097, 0.04750297, 0.0536674, 0.05221858, 0.0591969, 0.05249681, 
    0.04516535, 0.04131681, 0.04131365, 0.04297125, 0.04156278, 0.03986251, 
    0.03820841, 0.038367, 0.03844306, 0.03924319, 0.04157137, 0.0409135, 
    0.04100684, 0.04278716, 0.04546181, 0.04760295, 0.04753274, 0.04710601, 
    0.04798914, 0.04948514, 0.0511758, 0.0528729, 0.05337649, 0.05040234, 
    0.04738962, 0.04461123, 0.04190491, 0.04094056, 0.04095913, 0.03994371, 
    0.04154563, 0.04307092, 0.04242503, 0.0416563, 0.04128502, 0.04115636, 
    0.04183859, 0.04262061, 0.04253144, 0.04285748, 0.04211228, 0.04051074, 
    0.03923865, 0.0387577, 0.03976529, 0.04082646, 0.04149609, 0.04224632, 
    0.04393258, 0.04473015, 0.04474649, 0.04413119, 0.04489192, 0.04565612, 
    0.04633134, 0.04694059, 0.04886499, 0.05176988, 0.0537718, 0.05675332, 
    0.06085195, 0.06360766, 0.06347732, 0.06389817, 0.06426559, 0.06460677, 
    0.06536183, 0.0670553, 0.06904791, 0.06997377, 0.07276967, 0.073929, 
    0.07414602, 0.07225611, 0.07150038, 0.07172012, 0.07178549, 0.07129362, 
    0.06903721, 0.06713227, 0.06574564, 0.06580285, 0.06354906, 0.06299892, 
    0.06197849, 0.06170841, 0.06131686, 0.05966966, 0.05960434, 0.06034676, 
    0.06174026, 0.06343862, 0.06508336, 0.06602298, 0.06496532, 0.06398751, 
    0.06270327, 0.0609455, 0.06070479, 0.06289799, 0.06646334, 0.0676073, 
    0.06495104, 0.06435637, 0.06350721, 0.06276944, 0.0625688, 0.05784214, 
    0.05480119, 0.05248404, 0.04959929, 0.04624943, 0.0442449, 0.04110882, 
    0.03998068, 0.04084563, 0.04522492, 0.05752108, 0.06045457, 0.1094917, 
    0.039773, 0.03801006, 0.03629366, 0.03042199, 0.02749165, 0.04019714, 
    0.04577166, 0.03870305, 0.04938132, 0.04653253, 0.04125552, 0.04224965, 
    0.03516452, 0.02912178, 0.02284777, 0.02079876, 0.02156829, 0.02138568, 
    0.02036681, 0.02032711, 0.02118359, 0.02287856, 0.0249934, 0.02589203, 
    0.0262411, 0.02702974, 0.02783505, 0.02786598, 0.02832606, 0.02943308, 
    0.02944312, 0.02863683, 0.02944129, 0.03116157, 0.03178553, 0.0317596, 
    0.03287752, 0.03429758, 0.03613228, 0.03786765, 0.03863177, 0.0402466, 
    0.04181644, 0.04253935, 0.04173726, 0.04116941, 0.04085747, 0.04093088, 
    0.04183621, 0.04431884, 0.0484794, 0.05397245, 0.05991538, 0.06616119, 
    0.07653552, 0.0867709, 0.08421389, 0.07033145, 0.05847998, 0.05032317, 
    0.04941724, 0.04958304, 0.04748501, 0.0457765, 0.044891, 0.04756336,
  0.03997828, 0.03870878, 0.03848752, 0.04100916, 0.04582507, 0.04754359, 
    0.04051711, 0.0332262, 0.03262441, 0.0309905, 0.02619477, 0.02411005, 
    0.02620248, 0.02781825, 0.02804486, 0.02684094, 0.02703077, 0.0273814, 
    0.02618516, 0.02476367, 0.024482, 0.02455171, 0.02734926, 0.03071219, 
    0.03365743, 0.03709928, 0.04534244, 0.05431744, 0.08162425, 0.09159822, 
    0.0694828, 0.07243576, 0.05147019, 0.03806145, 0.03563755, 0.03407341, 
    0.03071778, 0.02552128, 0.02281559, 0.02052365, 0.02342955, 0.02160219, 
    0.01946764, 0.01984827, 0.02019606, 0.02153398, 0.02310726, 0.02482209, 
    0.02709345, 0.02845452, 0.02965465, 0.03015797, 0.03075465, 0.03122935, 
    0.03122908, 0.03161474, 0.03243589, 0.03421813, 0.03601543, 0.04453954, 
    0.05373995, 0.05888622, 0.05139828, 0.04740247, 0.03511707, 0.03403303, 
    0.03415851, 0.03442381, 0.03441897, 0.03470892, 0.03480029, 0.03534764, 
    0.03705932, 0.03727532, 0.03561849, 0.03464852, 0.0352032, 0.04017667, 
    0.04377727, 0.04650229, 0.05063318, 0.05323775, 0.05524775, 0.06236084, 
    0.07327502, 0.06391285, 0.04952203, 0.05337176, 0.05462858, 0.0516029, 
    0.05108476, 0.0514176, 0.05034689, 0.04965185, 0.0462477, 0.0457121, 
    0.04656895, 0.04895217, 0.05437922, 0.05315885, 0.05552051, 0.05016448, 
    0.04472202, 0.0433638, 0.04317401, 0.04371766, 0.04307767, 0.04094559, 
    0.03975626, 0.04040264, 0.04040265, 0.04132273, 0.04348723, 0.04272375, 
    0.04153671, 0.04242232, 0.04414303, 0.04534879, 0.04518368, 0.04508527, 
    0.04690743, 0.04920235, 0.0483863, 0.04746491, 0.04641666, 0.04349727, 
    0.04186701, 0.04108496, 0.03923813, 0.0375495, 0.03681505, 0.03567511, 
    0.0365365, 0.03703181, 0.03633812, 0.03612553, 0.03528579, 0.0351278, 
    0.03497874, 0.03545073, 0.03600366, 0.0372095, 0.03588628, 0.03408862, 
    0.03244696, 0.03113566, 0.03131747, 0.03235496, 0.03313051, 0.03391677, 
    0.03540835, 0.03663673, 0.03643131, 0.03578661, 0.03718529, 0.0381637, 
    0.03823485, 0.03881703, 0.04081223, 0.04344816, 0.04404462, 0.04599359, 
    0.04871485, 0.0493684, 0.04893864, 0.05022159, 0.05119708, 0.05249871, 
    0.05236964, 0.05379736, 0.05429583, 0.05529116, 0.05886835, 0.06055584, 
    0.05954501, 0.05877551, 0.05823841, 0.05739383, 0.05772235, 0.05900364, 
    0.0581154, 0.05694794, 0.05558817, 0.05484352, 0.05338345, 0.05227126, 
    0.05213902, 0.0514241, 0.04981751, 0.04918749, 0.04910534, 0.0503267, 
    0.05390897, 0.05547953, 0.05510161, 0.05472238, 0.05310351, 0.05187152, 
    0.04996871, 0.04991869, 0.05149843, 0.05384918, 0.05796472, 0.05870146, 
    0.05493598, 0.05428218, 0.05357856, 0.05278294, 0.05439365, 0.05020693, 
    0.04712667, 0.04558633, 0.04268004, 0.03856858, 0.03711095, 0.03532035, 
    0.03368749, 0.03386727, 0.03748293, 0.04960413, 0.084494, 0.04980523, 
    0.03677262, 0.02761763, 0.02261284, 0.01827079, 0.01613044, 0.02482113, 
    0.03254621, 0.04772742, 0.04250146, 0.02753046, 0.04046216, 0.03085615, 
    0.0221441, 0.01589947, 0.01375737, 0.01753005, 0.01493174, 0.01802761, 
    0.01899662, 0.01940418, 0.0200738, 0.02116543, 0.02248058, 0.02268157, 
    0.02288123, 0.02311584, 0.02342043, 0.02339726, 0.02386734, 0.02514322, 
    0.02506992, 0.02504603, 0.02556923, 0.02671918, 0.02707899, 0.02829147, 
    0.02987824, 0.03103482, 0.03194971, 0.03253546, 0.03245488, 0.0321121, 
    0.0328195, 0.03255368, 0.03206301, 0.03211818, 0.03254857, 0.03354697, 
    0.03486929, 0.03729688, 0.04120562, 0.04538037, 0.04951555, 0.05302873, 
    0.06399308, 0.0694898, 0.06051235, 0.0536248, 0.05099769, 0.04612081, 
    0.04457822, 0.04429559, 0.0424459, 0.04167034, 0.040625, 0.04080464,
  0.03235443, 0.03160951, 0.03173342, 0.03355442, 0.03448526, 0.03144761, 
    0.02741059, 0.02643056, 0.02595047, 0.02293875, 0.02027255, 0.01980363, 
    0.02148061, 0.02296366, 0.02396805, 0.02340095, 0.02387403, 0.02448794, 
    0.02350365, 0.02054721, 0.01966895, 0.01940923, 0.02129643, 0.0233198, 
    0.02423265, 0.02695904, 0.03243052, 0.04113997, 0.06684686, 0.06997207, 
    0.06086294, 0.06914782, 0.04192451, 0.03015241, 0.02962259, 0.02763331, 
    0.02213499, 0.01897665, 0.01971453, 0.02258935, 0.02939256, 0.02092902, 
    0.01815036, 0.01871771, 0.019106, 0.01990863, 0.02143557, 0.02301207, 
    0.0247839, 0.02705208, 0.02918329, 0.02955902, 0.03088156, 0.03257225, 
    0.03311878, 0.03404939, 0.03515854, 0.03616328, 0.0400681, 0.05262887, 
    0.0686128, 0.07111067, 0.05568508, 0.05696884, 0.0424494, 0.03660911, 
    0.03583394, 0.03707758, 0.03778972, 0.03886616, 0.03944859, 0.04024151, 
    0.04241038, 0.04184856, 0.03950355, 0.0383807, 0.0385714, 0.0438203, 
    0.05023097, 0.05195074, 0.05726242, 0.06358664, 0.06750093, 0.07768124, 
    0.09464266, 0.08361024, 0.07163639, 0.0667384, 0.06427932, 0.05305653, 
    0.05103108, 0.05121494, 0.05042944, 0.04922518, 0.04784555, 0.04700495, 
    0.04801448, 0.05117773, 0.05286361, 0.05542836, 0.05507133, 0.04770989, 
    0.04680274, 0.04671932, 0.04610714, 0.04692172, 0.04630291, 0.04455021, 
    0.04361021, 0.04235347, 0.04082491, 0.04142794, 0.04218093, 0.04124021, 
    0.04117119, 0.0418039, 0.0430085, 0.04400562, 0.04459582, 0.04578887, 
    0.04650988, 0.04617547, 0.04304288, 0.0405922, 0.03914492, 0.03758027, 
    0.0360527, 0.03579828, 0.0347192, 0.03346306, 0.03219402, 0.03119597, 
    0.03139577, 0.03154049, 0.03152689, 0.03195115, 0.03129231, 0.03049809, 
    0.02939858, 0.02901844, 0.02979596, 0.03051353, 0.02904061, 0.0278626, 
    0.02724846, 0.02700539, 0.02712077, 0.0282371, 0.02832091, 0.02896069, 
    0.03021099, 0.03133956, 0.03090734, 0.03050237, 0.03199065, 0.03253043, 
    0.03327191, 0.03456939, 0.03591596, 0.03772784, 0.03888216, 0.0397498, 
    0.03975853, 0.03910813, 0.03980574, 0.04060775, 0.04160751, 0.04265528, 
    0.0424456, 0.0442926, 0.04553977, 0.04697709, 0.04924548, 0.04981599, 
    0.04893872, 0.04970983, 0.05082905, 0.04885212, 0.04850848, 0.0495663, 
    0.05005076, 0.05025965, 0.04944378, 0.0477754, 0.04675253, 0.0461644, 
    0.04482148, 0.04360357, 0.04253196, 0.04352214, 0.04497227, 0.04470849, 
    0.04652687, 0.04736081, 0.04592967, 0.04434146, 0.04368911, 0.04444972, 
    0.04437269, 0.04497273, 0.04670236, 0.04822524, 0.05129298, 0.05141786, 
    0.04731738, 0.04569169, 0.04529836, 0.04364087, 0.04423755, 0.04230098, 
    0.04040915, 0.03821307, 0.03452381, 0.03218791, 0.03184417, 0.03182912, 
    0.03283937, 0.03719202, 0.0378615, 0.04305206, 0.05944354, 0.04418153, 
    0.03092393, 0.02348132, 0.01953756, 0.01533191, 0.01266916, 0.0139463, 
    0.01673098, 0.0156757, 0.01359603, 0.01270003, 0.01484409, 0.01137073, 
    0.009053725, 0.009726174, 0.00987025, 0.01196122, 0.01427017, 0.01656247, 
    0.01744114, 0.01758334, 0.01773756, 0.0184305, 0.01947915, 0.0195532, 
    0.01964524, 0.01976613, 0.02045142, 0.02122699, 0.02186241, 0.02245639, 
    0.02233897, 0.02245531, 0.02271058, 0.02391047, 0.02484862, 0.02613353, 
    0.02810287, 0.02925189, 0.0290363, 0.0289737, 0.02929547, 0.02875745, 
    0.02826648, 0.02649315, 0.02519712, 0.02501216, 0.02559157, 0.02632086, 
    0.02723015, 0.02907185, 0.03235396, 0.03584901, 0.03807421, 0.04190736, 
    0.04941771, 0.05107301, 0.0435161, 0.04208193, 0.04372218, 0.03925268, 
    0.03802988, 0.03825099, 0.03732712, 0.03744949, 0.03531939, 0.03335179,
  0.02508, 0.0237471, 0.02350391, 0.02433984, 0.02360442, 0.02110801, 
    0.01984968, 0.01997036, 0.01834631, 0.01657701, 0.01595876, 0.01560086, 
    0.01624833, 0.01765085, 0.01812766, 0.01906255, 0.02118778, 0.02260468, 
    0.02187904, 0.01702643, 0.01454332, 0.01443169, 0.01466806, 0.01513597, 
    0.01630233, 0.01939358, 0.02297171, 0.03059616, 0.04894596, 0.05934116, 
    0.05382782, 0.05810773, 0.03487825, 0.02065819, 0.0256346, 0.0293211, 
    0.02387012, 0.02012681, 0.02009202, 0.02000977, 0.01996903, 0.01956929, 
    0.01637556, 0.01830865, 0.01885176, 0.01983017, 0.02085929, 0.02192293, 
    0.02314929, 0.02513858, 0.02688801, 0.02846748, 0.0299489, 0.0319934, 
    0.03334285, 0.03517732, 0.03649477, 0.03713984, 0.04562338, 0.06421648, 
    0.09533307, 0.07554296, 0.05938982, 0.06379671, 0.05209186, 0.04176853, 
    0.04057616, 0.04236876, 0.04330065, 0.04410454, 0.04527495, 0.04656149, 
    0.04747501, 0.04746003, 0.04410894, 0.04282166, 0.0431476, 0.05108625, 
    0.05953934, 0.05973987, 0.06352647, 0.06831139, 0.07306401, 0.08850303, 
    0.1060327, 0.09862078, 0.0979448, 0.08066456, 0.07022907, 0.05386803, 
    0.05019724, 0.05063876, 0.05028781, 0.04846973, 0.04998714, 0.0509565, 
    0.0515361, 0.05409785, 0.05441127, 0.05331775, 0.05182277, 0.04778581, 
    0.0491035, 0.04924354, 0.0486021, 0.05088037, 0.04893349, 0.0474831, 
    0.04636316, 0.04434868, 0.04242213, 0.04199665, 0.04108701, 0.04069838, 
    0.04070417, 0.04266884, 0.04359921, 0.04383265, 0.04505996, 0.04479852, 
    0.04292936, 0.04058431, 0.03712754, 0.03445945, 0.03363613, 0.0337904, 
    0.03317795, 0.03185156, 0.0313979, 0.0302224, 0.02787724, 0.02646088, 
    0.02645913, 0.02684392, 0.0270083, 0.02783252, 0.02732262, 0.02658915, 
    0.02576494, 0.02528933, 0.0255801, 0.02569103, 0.02490076, 0.02465371, 
    0.024262, 0.02451135, 0.02498387, 0.02527163, 0.02507649, 0.02542402, 
    0.02590176, 0.0261542, 0.02554491, 0.02606412, 0.02792217, 0.02904683, 
    0.02996574, 0.03088211, 0.03223901, 0.03376296, 0.03475104, 0.03483207, 
    0.03464936, 0.03417428, 0.03480877, 0.03505941, 0.03539448, 0.03606908, 
    0.03636238, 0.03759265, 0.03958259, 0.0414315, 0.04323513, 0.04348134, 
    0.04398055, 0.04701229, 0.04657491, 0.04358801, 0.04381506, 0.04547044, 
    0.04688419, 0.04746599, 0.04773137, 0.04579363, 0.04392847, 0.04204032, 
    0.04087346, 0.04043116, 0.03945873, 0.04023384, 0.04155713, 0.04111438, 
    0.04179415, 0.04269164, 0.04064121, 0.03854927, 0.03836688, 0.03976943, 
    0.03999223, 0.04104261, 0.04200591, 0.04275541, 0.04318584, 0.04252132, 
    0.04005878, 0.03793012, 0.03620486, 0.03327337, 0.03340181, 0.03448134, 
    0.0332783, 0.03016024, 0.02712468, 0.02660118, 0.03467583, 0.04541321, 
    0.05027638, 0.05490664, 0.04397576, 0.04217553, 0.05224341, 0.03720846, 
    0.0259142, 0.02008105, 0.01659465, 0.01332657, 0.0109306, 0.009375196, 
    0.009548349, 0.009077369, 0.007893014, 0.007680221, 0.008316291, 
    0.008590562, 0.008568146, 0.009268796, 0.01088908, 0.01331439, 
    0.01486392, 0.01589817, 0.01589695, 0.01594578, 0.01580245, 0.01619194, 
    0.01721928, 0.01731481, 0.01743244, 0.01782529, 0.01847829, 0.01968351, 
    0.02020586, 0.02034675, 0.02086452, 0.0213927, 0.02190096, 0.02280927, 
    0.02434831, 0.02574706, 0.02696109, 0.02756785, 0.02757236, 0.02776943, 
    0.02810557, 0.02761509, 0.02694762, 0.02496507, 0.02246165, 0.02079507, 
    0.01991978, 0.02019412, 0.02066114, 0.02163436, 0.02332892, 0.02595245, 
    0.02798081, 0.03133332, 0.03538832, 0.03694556, 0.03504222, 0.03573772, 
    0.03621411, 0.03224405, 0.03187494, 0.03272185, 0.03305731, 0.03351091, 
    0.03113634, 0.0272391,
  0.02016461, 0.01890352, 0.01836026, 0.01759154, 0.01719389, 0.0156372, 
    0.01445293, 0.01307991, 0.01148957, 0.01122739, 0.01123835, 0.01090671, 
    0.01076702, 0.01182136, 0.01285355, 0.01490209, 0.01783333, 0.01842647, 
    0.01726652, 0.01451435, 0.01197678, 0.01070777, 0.009785932, 0.01001813, 
    0.0116634, 0.01477994, 0.01729565, 0.02285853, 0.03219442, 0.04533694, 
    0.04737991, 0.05026581, 0.02766549, 0.01986459, 0.03088256, 0.03410261, 
    0.02922808, 0.0234494, 0.02004668, 0.01949357, 0.01924444, 0.01851163, 
    0.01835216, 0.01962565, 0.01990469, 0.01975945, 0.02040688, 0.02145388, 
    0.02250167, 0.02335224, 0.02463471, 0.02696016, 0.02965137, 0.03205137, 
    0.03353112, 0.03559409, 0.03760184, 0.03856685, 0.05250308, 0.07442547, 
    0.1081322, 0.0702913, 0.06058434, 0.06553441, 0.05884997, 0.04965983, 
    0.04882069, 0.05072526, 0.05077828, 0.05071115, 0.05087554, 0.05071235, 
    0.05053881, 0.05204379, 0.04885711, 0.04632469, 0.04783949, 0.05717875, 
    0.06495478, 0.06972321, 0.07407786, 0.06819324, 0.07239847, 0.09147375, 
    0.1100793, 0.09913307, 0.0974304, 0.08181103, 0.06637192, 0.05057509, 
    0.04861492, 0.0485304, 0.0479342, 0.04764403, 0.05252648, 0.05328174, 
    0.05336057, 0.05938789, 0.06129044, 0.05562755, 0.05152585, 0.04843422, 
    0.05018037, 0.0506437, 0.05085767, 0.05156999, 0.04984153, 0.05026288, 
    0.04857009, 0.04696216, 0.04526616, 0.04336406, 0.04196451, 0.04060702, 
    0.04070528, 0.04237456, 0.04135104, 0.04165547, 0.04170009, 0.03942548, 
    0.03643261, 0.03443164, 0.03263386, 0.03107194, 0.03062711, 0.03114353, 
    0.03011831, 0.02864169, 0.02864107, 0.02715235, 0.02468558, 0.02311714, 
    0.02297475, 0.02373846, 0.02440787, 0.02472019, 0.02341827, 0.02292974, 
    0.02293397, 0.02304467, 0.02354008, 0.02375446, 0.02300337, 0.02276411, 
    0.02205148, 0.02187134, 0.02251278, 0.02202207, 0.02206808, 0.02307087, 
    0.02364264, 0.02363672, 0.02352009, 0.02456796, 0.02662726, 0.02845205, 
    0.02942184, 0.02958565, 0.03018131, 0.0305812, 0.03031194, 0.03067813, 
    0.02972595, 0.02911891, 0.03003506, 0.03098845, 0.03162929, 0.03193347, 
    0.03217936, 0.03195549, 0.03319522, 0.03459207, 0.03728019, 0.03817628, 
    0.03988243, 0.04254686, 0.04063203, 0.03991577, 0.04204405, 0.04497893, 
    0.04674165, 0.04696953, 0.04618721, 0.04544609, 0.04362508, 0.04166352, 
    0.04030944, 0.0393367, 0.03839951, 0.03827602, 0.03938695, 0.03978297, 
    0.04031254, 0.04022163, 0.03782906, 0.03551507, 0.03451137, 0.03444571, 
    0.03446021, 0.03573702, 0.03730717, 0.0372487, 0.03585201, 0.03492868, 
    0.03377078, 0.03202192, 0.02910334, 0.02691218, 0.02691819, 0.02840791, 
    0.02846156, 0.02629981, 0.02352973, 0.02970744, 0.04404677, 0.05084957, 
    0.05068427, 0.0515268, 0.04605769, 0.05253764, 0.05050614, 0.0350664, 
    0.0252212, 0.01873115, 0.01530928, 0.01268347, 0.01075044, 0.009446532, 
    0.008031462, 0.007466213, 0.007485079, 0.007905619, 0.008582563, 
    0.009154511, 0.009777199, 0.01070218, 0.01223709, 0.01390524, 0.01420817, 
    0.01486544, 0.01497826, 0.01498555, 0.0146468, 0.0148788, 0.01560124, 
    0.01591557, 0.01615644, 0.01668555, 0.01781417, 0.01944618, 0.02006724, 
    0.02031752, 0.02056934, 0.02118727, 0.0223911, 0.02296284, 0.02342036, 
    0.02474072, 0.0255228, 0.02632, 0.02819549, 0.02877143, 0.02875302, 
    0.02784814, 0.02652454, 0.02467916, 0.02277692, 0.0205854, 0.01838764, 
    0.01768175, 0.01687621, 0.01651554, 0.01708195, 0.01895773, 0.02041545, 
    0.02226868, 0.02529737, 0.02822633, 0.02977694, 0.03036153, 0.02937726, 
    0.02698614, 0.02654363, 0.02682755, 0.02658968, 0.02741053, 0.02540664, 
    0.02228396,
  0.01610748, 0.01530338, 0.01458969, 0.01277162, 0.01195156, 0.01069658, 
    0.009553052, 0.008146674, 0.00744105, 0.007483437, 0.007500464, 
    0.007452252, 0.007178525, 0.007601848, 0.008699956, 0.0103371, 
    0.01216961, 0.01181827, 0.01129694, 0.010966, 0.01028316, 0.008702671, 
    0.007549333, 0.007692436, 0.009053268, 0.01083893, 0.01253556, 
    0.01572463, 0.02025844, 0.02811142, 0.03586322, 0.03731788, 0.02254619, 
    0.01844628, 0.03137328, 0.03621767, 0.02752433, 0.02639882, 0.02506506, 
    0.02083658, 0.01909638, 0.01886475, 0.01892813, 0.01938559, 0.0196838, 
    0.01999524, 0.02012827, 0.02113887, 0.02252071, 0.02355783, 0.0250535, 
    0.02720157, 0.02983715, 0.03224938, 0.03438856, 0.03721903, 0.03911769, 
    0.04241756, 0.05854258, 0.0855777, 0.09127122, 0.06400412, 0.06025982, 
    0.06537817, 0.06517261, 0.06009693, 0.05967654, 0.06135421, 0.06012737, 
    0.05819021, 0.05698368, 0.05425395, 0.05285029, 0.05419365, 0.05246112, 
    0.05099699, 0.05358373, 0.06139185, 0.06835663, 0.07800313, 0.08255446, 
    0.06876647, 0.07204833, 0.08742806, 0.1027249, 0.1091911, 0.1285021, 
    0.08667903, 0.06068565, 0.04578502, 0.04609814, 0.04614987, 0.04466036, 
    0.04514412, 0.04823869, 0.05331564, 0.06535714, 0.07146154, 0.06869315, 
    0.0572677, 0.05318153, 0.05123673, 0.05134935, 0.05132017, 0.05204928, 
    0.05131076, 0.04880682, 0.05099926, 0.04930234, 0.04611772, 0.04435293, 
    0.04354419, 0.04208596, 0.0411992, 0.04030648, 0.0396677, 0.03841649, 
    0.03801466, 0.03682688, 0.03424904, 0.03204118, 0.03085395, 0.0297465, 
    0.02918428, 0.02903191, 0.02852723, 0.02683081, 0.02511591, 0.02490269, 
    0.02375532, 0.02206062, 0.02112068, 0.02112664, 0.02199032, 0.02255854, 
    0.02164994, 0.01983338, 0.0197839, 0.02092437, 0.02186719, 0.02222977, 
    0.02162952, 0.02049677, 0.02038684, 0.02031753, 0.02048284, 0.02088097, 
    0.02111072, 0.02118492, 0.02230559, 0.0231877, 0.02290812, 0.02341926, 
    0.02422053, 0.02565358, 0.02682155, 0.02692973, 0.02663684, 0.02730785, 
    0.02772221, 0.02765046, 0.02816879, 0.02738729, 0.0272218, 0.02767554, 
    0.02837571, 0.02908499, 0.02994126, 0.03001635, 0.0296311, 0.02973049, 
    0.03094432, 0.0334142, 0.03514151, 0.03740128, 0.03821503, 0.03764498, 
    0.0399879, 0.04329658, 0.04594672, 0.04661143, 0.046348, 0.04589263, 
    0.04559019, 0.04436357, 0.04322137, 0.04240309, 0.04034182, 0.03929956, 
    0.03972402, 0.04096247, 0.0398926, 0.03871859, 0.03741343, 0.03578497, 
    0.03410967, 0.03302717, 0.03229476, 0.0323512, 0.0329204, 0.03269839, 
    0.03175214, 0.03100688, 0.03141212, 0.03038299, 0.02899104, 0.02530319, 
    0.02290094, 0.02386432, 0.02866611, 0.02975371, 0.0298067, 0.03507595, 
    0.05103573, 0.05427011, 0.07593341, 0.08808193, 0.08407556, 0.06708135, 
    0.06067909, 0.04600238, 0.03211862, 0.02483513, 0.01897454, 0.01538865, 
    0.0130058, 0.01119859, 0.01023908, 0.009414856, 0.008991869, 0.008972801, 
    0.009316781, 0.009793905, 0.01032427, 0.01100173, 0.01187488, 0.01294456, 
    0.01357124, 0.01363117, 0.01451136, 0.01436907, 0.01472216, 0.0144722, 
    0.01435707, 0.01451788, 0.01503122, 0.01570154, 0.01657392, 0.0179755, 
    0.01928156, 0.01954072, 0.01995447, 0.02035363, 0.0205825, 0.02178526, 
    0.02275264, 0.02305509, 0.02442823, 0.02550246, 0.02667584, 0.02912493, 
    0.02964237, 0.0295511, 0.02889361, 0.027102, 0.02467863, 0.022829, 
    0.020093, 0.01663128, 0.01523947, 0.01459019, 0.01398646, 0.01360987, 
    0.01502001, 0.01542962, 0.01638556, 0.01871956, 0.02119825, 0.02310467, 
    0.02293622, 0.02208387, 0.02149703, 0.0215233, 0.02134715, 0.02024815, 
    0.01962199, 0.01802506, 0.01674645,
  0.01168711, 0.01125663, 0.01040068, 0.009871063, 0.009367652, 0.008295923, 
    0.007159337, 0.006268261, 0.005835506, 0.005676517, 0.005568454, 
    0.005490561, 0.005565692, 0.005723927, 0.00598488, 0.006693001, 
    0.007816125, 0.007714409, 0.007261633, 0.006877996, 0.006708515, 
    0.005776621, 0.005417494, 0.005956422, 0.006495594, 0.007309003, 
    0.007951847, 0.009821903, 0.01240129, 0.01512301, 0.02120343, 0.02856301, 
    0.01644387, 0.01580497, 0.02506646, 0.03161482, 0.02344039, 0.01865574, 
    0.01706543, 0.01880082, 0.01950027, 0.02003404, 0.01977356, 0.01937473, 
    0.01818289, 0.01852524, 0.01963137, 0.0208649, 0.02260694, 0.02422219, 
    0.02620189, 0.02868195, 0.03037846, 0.03245668, 0.0354215, 0.03872982, 
    0.04051501, 0.04948655, 0.06665295, 0.1127843, 0.07997327, 0.06634888, 
    0.06443554, 0.06896889, 0.0754276, 0.07304032, 0.07159138, 0.06980636, 
    0.06611226, 0.06225792, 0.05919398, 0.05488981, 0.05110101, 0.0513465, 
    0.05160816, 0.05463478, 0.05676373, 0.06106199, 0.06953989, 0.0788903, 
    0.08076126, 0.06787736, 0.07273587, 0.08806399, 0.09467342, 0.1264091, 
    0.1346252, 0.08780649, 0.05751515, 0.0475416, 0.04654769, 0.04563282, 
    0.04475507, 0.0449142, 0.04632768, 0.05531653, 0.07373435, 0.07419277, 
    0.07163675, 0.05855321, 0.05688618, 0.05685022, 0.05586634, 0.05454532, 
    0.0546784, 0.05183602, 0.04847606, 0.04790471, 0.04684733, 0.04228114, 
    0.04153856, 0.04131879, 0.04088479, 0.04062454, 0.03941935, 0.03802959, 
    0.03635156, 0.03418987, 0.03217062, 0.03079839, 0.02935303, 0.02905495, 
    0.02803302, 0.02756142, 0.02747288, 0.0272177, 0.024925, 0.02281414, 
    0.02218232, 0.021258, 0.01991781, 0.01923054, 0.01955472, 0.02000921, 
    0.01983006, 0.01887439, 0.01797515, 0.01832812, 0.02005161, 0.02121021, 
    0.0210141, 0.02052374, 0.02014542, 0.0198295, 0.01959923, 0.01963758, 
    0.02049076, 0.02085647, 0.02058262, 0.02123697, 0.02195949, 0.0221099, 
    0.0223709, 0.02307172, 0.02409363, 0.02426461, 0.02388683, 0.02399165, 
    0.02476804, 0.02507408, 0.02492851, 0.02534519, 0.0252472, 0.02569964, 
    0.02666848, 0.02751629, 0.0278037, 0.02861944, 0.02820183, 0.02789271, 
    0.02789047, 0.02859508, 0.03068041, 0.03314817, 0.03565761, 0.03594898, 
    0.03681936, 0.03970026, 0.04253916, 0.04446965, 0.04541802, 0.04626308, 
    0.04655289, 0.04701855, 0.04663114, 0.04573386, 0.044753, 0.04295672, 
    0.04109782, 0.04115695, 0.04232922, 0.04054852, 0.03777155, 0.03636487, 
    0.0347858, 0.03215881, 0.03046227, 0.03079485, 0.03106518, 0.03100761, 
    0.03035568, 0.02875252, 0.02883848, 0.03143656, 0.02910277, 0.0282228, 
    0.02539453, 0.02446148, 0.02976687, 0.03496904, 0.02668835, 0.02584716, 
    0.03967413, 0.05393514, 0.06703799, 0.09448882, 0.08914185, 0.07374508, 
    0.08072658, 0.06625652, 0.04109123, 0.02751749, 0.02331533, 0.01866618, 
    0.01574047, 0.01353176, 0.0114681, 0.01037946, 0.009664015, 0.009481376, 
    0.009905308, 0.01081428, 0.01157685, 0.01191023, 0.01221941, 0.01262726, 
    0.01271386, 0.01252627, 0.01314576, 0.01474877, 0.01448852, 0.01468707, 
    0.01440969, 0.0140891, 0.01441581, 0.01506678, 0.01628069, 0.01760649, 
    0.01850324, 0.01961431, 0.02012572, 0.02014493, 0.02079657, 0.02096039, 
    0.02152298, 0.0226778, 0.0238422, 0.02546029, 0.02657239, 0.02741724, 
    0.02916019, 0.03024135, 0.03017853, 0.02955074, 0.02820802, 0.02574763, 
    0.02304897, 0.01928594, 0.01537027, 0.01366877, 0.01316614, 0.01221792, 
    0.01129312, 0.01189723, 0.01226916, 0.01252293, 0.01387507, 0.01580339, 
    0.01667828, 0.01586098, 0.01517809, 0.01549585, 0.01603703, 0.01600219, 
    0.01492347, 0.01337709, 0.01196034, 0.01147327,
  0.00903447, 0.008687605, 0.008115077, 0.0080799, 0.008656112, 0.008676129, 
    0.007554217, 0.005959958, 0.005098039, 0.004513472, 0.004545443, 
    0.004764826, 0.005296148, 0.005576907, 0.005323693, 0.005146592, 
    0.005686069, 0.006047673, 0.00539159, 0.004501959, 0.004033788, 
    0.003736312, 0.003898514, 0.004305294, 0.004891765, 0.005634164, 
    0.005727335, 0.006595725, 0.007651705, 0.00853772, 0.01426199, 
    0.01706542, 0.01102481, 0.01507167, 0.02204272, 0.02102703, 0.01823837, 
    0.01660861, 0.01451515, 0.01389121, 0.01453905, 0.01901018, 0.02165846, 
    0.01886048, 0.01736932, 0.0176933, 0.01875251, 0.02047721, 0.02244449, 
    0.0246772, 0.02721913, 0.03050028, 0.03296695, 0.03541869, 0.03749864, 
    0.04041968, 0.04323931, 0.05596945, 0.07605604, 0.1251301, 0.08207154, 
    0.07769727, 0.0722465, 0.07616086, 0.08760322, 0.08259008, 0.08040725, 
    0.08067239, 0.07070855, 0.06340525, 0.05842065, 0.05427751, 0.05033938, 
    0.04732343, 0.04822573, 0.05759478, 0.06464434, 0.06329452, 0.06688306, 
    0.07298237, 0.07578586, 0.06628214, 0.07794228, 0.08798631, 0.09409662, 
    0.1270689, 0.1074347, 0.07850643, 0.05892977, 0.05241478, 0.04883722, 
    0.04609837, 0.04462536, 0.04536152, 0.04780783, 0.05668653, 0.09171937, 
    0.09242886, 0.07342216, 0.06158974, 0.06355123, 0.06185377, 0.05834008, 
    0.05844238, 0.05907997, 0.05325926, 0.04893709, 0.04630999, 0.04359947, 
    0.04051408, 0.0397518, 0.0400984, 0.04148098, 0.04183143, 0.03997142, 
    0.038159, 0.03512419, 0.03089115, 0.02909359, 0.02839635, 0.0274093, 
    0.02720543, 0.02623811, 0.02588891, 0.02626828, 0.02618465, 0.02468168, 
    0.02285232, 0.02142055, 0.02032265, 0.01899783, 0.01893634, 0.018569, 
    0.01783574, 0.01760287, 0.017641, 0.01797865, 0.01821144, 0.01964547, 
    0.02035365, 0.01982922, 0.01994992, 0.01996625, 0.0193427, 0.01903735, 
    0.0190503, 0.01956642, 0.01979662, 0.0200444, 0.02066992, 0.0218303, 
    0.02227087, 0.02229346, 0.0229654, 0.02366948, 0.02372594, 0.02316443, 
    0.02297304, 0.02316787, 0.02247082, 0.02213397, 0.0228728, 0.02317458, 
    0.02417211, 0.0261612, 0.0268788, 0.02644288, 0.02619787, 0.02601238, 
    0.02619934, 0.02666983, 0.02739176, 0.02970194, 0.03203192, 0.03448027, 
    0.03565126, 0.03695979, 0.03929896, 0.0415764, 0.0436017, 0.04518836, 
    0.04696682, 0.04852352, 0.04843189, 0.04834151, 0.04801503, 0.04594243, 
    0.0439638, 0.0425541, 0.04179562, 0.04112219, 0.03881365, 0.0364126, 
    0.03520785, 0.03324126, 0.03089522, 0.02964217, 0.02978421, 0.02963451, 
    0.02965862, 0.02892733, 0.02779332, 0.02691504, 0.02751839, 0.02720777, 
    0.02847929, 0.02846342, 0.03211563, 0.04541585, 0.04761249, 0.05928206, 
    0.07255484, 0.0781929, 0.08796069, 0.09929927, 0.09425708, 0.07754953, 
    0.06022802, 0.04996587, 0.03588331, 0.02743746, 0.0241184, 0.02150801, 
    0.01770113, 0.01580251, 0.01432933, 0.01335145, 0.01147128, 0.01005833, 
    0.009911046, 0.01084332, 0.01289655, 0.01353359, 0.01336485, 0.01336702, 
    0.01349, 0.01368561, 0.01334596, 0.01448035, 0.01527416, 0.01445956, 
    0.01435115, 0.01407039, 0.01393492, 0.01460835, 0.01577416, 0.01708508, 
    0.01870959, 0.01938493, 0.02012312, 0.02066985, 0.0209128, 0.0210257, 
    0.02092618, 0.02143303, 0.02270133, 0.02450754, 0.02673333, 0.0283173, 
    0.02860226, 0.02970557, 0.03127772, 0.0310281, 0.03012543, 0.02856839, 
    0.02642079, 0.0233781, 0.01886499, 0.01505258, 0.01280864, 0.01173592, 
    0.01007441, 0.008888029, 0.00892054, 0.01015758, 0.01034065, 0.01058313, 
    0.01167832, 0.0119687, 0.01135272, 0.01133673, 0.0111659, 0.01085795, 
    0.01077435, 0.01087875, 0.01000335, 0.008881142, 0.008699339,
  0.007753585, 0.006784381, 0.006525178, 0.007051419, 0.008262324, 
    0.00963832, 0.008135275, 0.005557242, 0.004861161, 0.004164673, 
    0.003822028, 0.004312922, 0.005201898, 0.005969117, 0.005432609, 
    0.004204097, 0.004203511, 0.004637901, 0.004810847, 0.003983392, 
    0.003456997, 0.003135303, 0.0030929, 0.003269239, 0.003931056, 
    0.004601841, 0.004949554, 0.005560398, 0.00569245, 0.007629265, 
    0.01394596, 0.01164523, 0.00985492, 0.01513402, 0.02111028, 0.01672024, 
    0.01588738, 0.01386328, 0.01240266, 0.01223577, 0.01190597, 0.01329463, 
    0.01660659, 0.01543952, 0.01435361, 0.01556101, 0.01692307, 0.01845131, 
    0.02090242, 0.0243173, 0.02794679, 0.0316367, 0.03489561, 0.03832361, 
    0.04103557, 0.04303128, 0.04584913, 0.05829441, 0.09015651, 0.1135034, 
    0.08835796, 0.08815354, 0.08212982, 0.08575658, 0.09718871, 0.08937608, 
    0.08516779, 0.08576433, 0.07351324, 0.06289357, 0.05634611, 0.05140327, 
    0.04698972, 0.04399518, 0.04638458, 0.0568676, 0.06894819, 0.07156204, 
    0.06789406, 0.07109904, 0.07160126, 0.07020257, 0.081749, 0.08671233, 
    0.1110203, 0.1069899, 0.08358923, 0.06319906, 0.06131338, 0.05724051, 
    0.05314726, 0.05028965, 0.04745216, 0.04768857, 0.05079933, 0.05541373, 
    0.08195435, 0.1025977, 0.07948954, 0.0654964, 0.06951401, 0.06838081, 
    0.06299975, 0.06096458, 0.05779035, 0.05375465, 0.05082886, 0.04804054, 
    0.04441456, 0.04098564, 0.03995524, 0.04151735, 0.04227209, 0.04199117, 
    0.04024033, 0.03797745, 0.03452103, 0.0299553, 0.02821023, 0.02756901, 
    0.02640497, 0.02590926, 0.02615049, 0.0256384, 0.02536703, 0.02512555, 
    0.02441938, 0.02264459, 0.02160702, 0.02082807, 0.02060786, 0.02068279, 
    0.01926982, 0.01732746, 0.01707796, 0.01788585, 0.01833704, 0.01882518, 
    0.01953761, 0.01937179, 0.01874192, 0.01910309, 0.01957276, 0.01947834, 
    0.01921107, 0.01939205, 0.01901888, 0.0188888, 0.01968664, 0.02082964, 
    0.02184142, 0.02259798, 0.02343882, 0.02392778, 0.02365396, 0.02302406, 
    0.02273643, 0.02265687, 0.02247604, 0.02143472, 0.02103024, 0.02184869, 
    0.02225151, 0.02408784, 0.02692375, 0.02652416, 0.02534382, 0.02490105, 
    0.02514585, 0.02554682, 0.02605838, 0.02701078, 0.02946508, 0.03239202, 
    0.03492819, 0.03609746, 0.03671659, 0.0386003, 0.04106402, 0.04315009, 
    0.04473774, 0.04639271, 0.04863109, 0.04873926, 0.04888349, 0.04871596, 
    0.04718885, 0.0445472, 0.04264302, 0.04106945, 0.03908262, 0.03643633, 
    0.03474147, 0.03332677, 0.03146177, 0.02924472, 0.0285938, 0.02856735, 
    0.02694348, 0.02627731, 0.02676107, 0.02582738, 0.02335021, 0.02343502, 
    0.02651108, 0.03059348, 0.03535338, 0.04518257, 0.05615528, 0.05404948, 
    0.09427119, 0.097991, 0.08950683, 0.08446787, 0.08044276, 0.06533304, 
    0.0582937, 0.04397235, 0.03864735, 0.02962757, 0.0240549, 0.02123196, 
    0.01980085, 0.01710703, 0.01546524, 0.01345843, 0.01318138, 0.01229056, 
    0.01041116, 0.01116086, 0.01221673, 0.01325252, 0.01368611, 0.01362572, 
    0.01310376, 0.01361919, 0.01411682, 0.01448384, 0.01547239, 0.01543731, 
    0.01462738, 0.01441622, 0.01440334, 0.01461455, 0.01515571, 0.01612421, 
    0.01729459, 0.01852671, 0.01956479, 0.02003212, 0.02083769, 0.02147079, 
    0.02126954, 0.02108756, 0.02166199, 0.02306836, 0.02487036, 0.02680976, 
    0.02910125, 0.02926323, 0.03015749, 0.03090375, 0.03065573, 0.03017648, 
    0.02879002, 0.02632829, 0.02330861, 0.01873624, 0.01465764, 0.01186758, 
    0.01012849, 0.008560187, 0.007468735, 0.006963547, 0.008103327, 
    0.008386553, 0.008350308, 0.008717845, 0.008749854, 0.008661444, 
    0.008847686, 0.008257618, 0.007616691, 0.007633396, 0.00806369, 
    0.007887067, 0.007479053, 0.00760779,
  0.007258384, 0.006235531, 0.005609326, 0.006195896, 0.006787999, 
    0.008346992, 0.007427043, 0.005476501, 0.005013539, 0.004210135, 
    0.003630922, 0.004048037, 0.005113466, 0.006631746, 0.006328603, 
    0.004320565, 0.003520834, 0.003691637, 0.00407452, 0.003775409, 
    0.003578003, 0.003134639, 0.002864667, 0.002856966, 0.00329208, 
    0.003459089, 0.004106801, 0.004930206, 0.005554093, 0.01055085, 
    0.01109976, 0.008218122, 0.009845443, 0.01340653, 0.01718051, 0.01510003, 
    0.01434339, 0.01276099, 0.01142968, 0.01084332, 0.01080952, 0.01088936, 
    0.01033906, 0.01016108, 0.01137423, 0.01355666, 0.01503067, 0.016045, 
    0.01857833, 0.02248329, 0.02682786, 0.03120841, 0.03513503, 0.03869775, 
    0.04127291, 0.04424527, 0.04869985, 0.06008269, 0.1025944, 0.1029485, 
    0.08863429, 0.09067316, 0.08657161, 0.0918187, 0.09885789, 0.0886414, 
    0.07884369, 0.07965294, 0.07150476, 0.06201443, 0.05309238, 0.04711478, 
    0.04314233, 0.04234959, 0.04797936, 0.05933155, 0.0695036, 0.07588621, 
    0.06983854, 0.07390583, 0.07609054, 0.07513173, 0.08656347, 0.09628636, 
    0.1190761, 0.09847705, 0.0681199, 0.06426505, 0.06735731, 0.06201316, 
    0.05782315, 0.05588946, 0.05222413, 0.05240488, 0.05594837, 0.05695086, 
    0.0727002, 0.08842977, 0.07452358, 0.06468296, 0.06848474, 0.06869777, 
    0.06433808, 0.06161974, 0.05897752, 0.05629015, 0.05330674, 0.05023266, 
    0.04646759, 0.04295355, 0.04214499, 0.0452106, 0.04717685, 0.04546073, 
    0.04108043, 0.03848562, 0.0352897, 0.0312847, 0.02897839, 0.02870847, 
    0.02759211, 0.02655273, 0.02663869, 0.02593752, 0.02467429, 0.02378342, 
    0.02259444, 0.02241093, 0.02264327, 0.02208336, 0.0222397, 0.02223055, 
    0.02059823, 0.01868144, 0.0185339, 0.0193912, 0.0196648, 0.02002979, 
    0.02082043, 0.02003868, 0.01899173, 0.01939953, 0.01994325, 0.01996291, 
    0.02066216, 0.0207635, 0.01977862, 0.01910668, 0.01951461, 0.02068508, 
    0.02156102, 0.0222423, 0.02361283, 0.02484868, 0.02429151, 0.02319657, 
    0.02258714, 0.02260891, 0.02229106, 0.02116804, 0.02075163, 0.02090842, 
    0.02164434, 0.02512774, 0.02939842, 0.02729228, 0.0256334, 0.02453121, 
    0.0246805, 0.02499682, 0.02587277, 0.02729139, 0.02985428, 0.03296492, 
    0.03557651, 0.03785349, 0.03853264, 0.04013859, 0.04212809, 0.04426078, 
    0.04611875, 0.04673027, 0.04795553, 0.04839559, 0.04833763, 0.04832437, 
    0.04743496, 0.04491139, 0.04202227, 0.03945553, 0.03710594, 0.03422358, 
    0.0322586, 0.03028214, 0.02856383, 0.02677834, 0.02605002, 0.02516814, 
    0.02304815, 0.02193715, 0.02212961, 0.021927, 0.02124615, 0.02381041, 
    0.02803979, 0.03351258, 0.0423225, 0.05404889, 0.05554513, 0.06725167, 
    0.09084199, 0.08531063, 0.06986044, 0.05585004, 0.04995721, 0.0457255, 
    0.04153714, 0.0330993, 0.03041184, 0.02502768, 0.02136479, 0.01964781, 
    0.01896272, 0.01716661, 0.0151548, 0.01324844, 0.01459256, 0.01360488, 
    0.01252557, 0.01907543, 0.02632431, 0.02602786, 0.01559479, 0.01338338, 
    0.01295793, 0.0142167, 0.01376572, 0.01434357, 0.01499485, 0.01464212, 
    0.0145191, 0.01498643, 0.01511546, 0.0151599, 0.01534853, 0.01629594, 
    0.0172249, 0.01788712, 0.01915288, 0.02013087, 0.02097565, 0.02143888, 
    0.02173948, 0.02207858, 0.02278485, 0.02434298, 0.02520603, 0.02645333, 
    0.02834639, 0.02908856, 0.0300161, 0.03014055, 0.03014223, 0.02982764, 
    0.02844085, 0.02610241, 0.02322197, 0.01961047, 0.01453756, 0.01118798, 
    0.009068477, 0.007411716, 0.006562844, 0.005953458, 0.006577306, 
    0.007176104, 0.007220505, 0.007367639, 0.007271159, 0.007045889, 
    0.00706326, 0.006567909, 0.005992893, 0.006084485, 0.006234759, 
    0.006431158, 0.00655375, 0.0069425,
  0.006786912, 0.005959551, 0.005144694, 0.00543344, 0.005450346, 
    0.006046168, 0.005791393, 0.005259784, 0.004983427, 0.00408761, 
    0.003776548, 0.004161039, 0.005952112, 0.008992709, 0.008491745, 
    0.005099519, 0.003898023, 0.003423208, 0.003390614, 0.003430321, 
    0.003438423, 0.003202312, 0.003042471, 0.002736675, 0.002807983, 
    0.002712051, 0.003320489, 0.004231938, 0.005088241, 0.008270741, 
    0.007640856, 0.007639115, 0.01007217, 0.01251032, 0.01398958, 0.01393702, 
    0.01291193, 0.01166803, 0.01087715, 0.01043979, 0.01009315, 0.009785984, 
    0.009717949, 0.00973177, 0.009744993, 0.01111461, 0.01266648, 0.0140064, 
    0.01580286, 0.01883971, 0.02307505, 0.02806758, 0.03282159, 0.03722422, 
    0.04081502, 0.04568738, 0.05312777, 0.06415325, 0.1030129, 0.09432058, 
    0.08608758, 0.0909962, 0.08980031, 0.09412333, 0.09622307, 0.08469338, 
    0.07513909, 0.07368068, 0.06563134, 0.05762243, 0.0484624, 0.04339559, 
    0.04057851, 0.04310177, 0.05236043, 0.06292811, 0.06701159, 0.07443567, 
    0.07011048, 0.07872681, 0.07906599, 0.08487912, 0.0848465, 0.1080111, 
    0.1123018, 0.09442063, 0.07006019, 0.07789519, 0.07667498, 0.06463084, 
    0.05965644, 0.05969696, 0.05778738, 0.05839674, 0.06084371, 0.06251764, 
    0.06799979, 0.07113765, 0.06631999, 0.06142544, 0.0632911, 0.06488235, 
    0.06293589, 0.06105046, 0.05963137, 0.05710212, 0.05593666, 0.05340295, 
    0.04874035, 0.04543286, 0.04471818, 0.04723703, 0.04924444, 0.04758622, 
    0.04249735, 0.03918325, 0.03597708, 0.03246614, 0.03077402, 0.03065976, 
    0.02991009, 0.02931915, 0.02886926, 0.02715923, 0.02514089, 0.02418847, 
    0.0225292, 0.02298749, 0.0232058, 0.02312192, 0.02220486, 0.02186589, 
    0.02057846, 0.01937942, 0.01968203, 0.02030594, 0.02102918, 0.02228964, 
    0.02303396, 0.02181977, 0.02099428, 0.02130907, 0.02137683, 0.0213566, 
    0.0221076, 0.02172543, 0.02128334, 0.02055104, 0.02042068, 0.02137666, 
    0.02200056, 0.0221584, 0.02312727, 0.02466705, 0.02437697, 0.02395892, 
    0.02344159, 0.02323058, 0.02299155, 0.02148718, 0.0200525, 0.01887509, 
    0.02195331, 0.05703277, 0.0402325, 0.02883429, 0.02602605, 0.02441086, 
    0.02418666, 0.02478022, 0.02577309, 0.02728356, 0.03021421, 0.03270445, 
    0.03625293, 0.03934038, 0.04106831, 0.04258906, 0.0436454, 0.04540715, 
    0.04734493, 0.04796236, 0.04823864, 0.0485394, 0.04835141, 0.04702264, 
    0.04653496, 0.04449639, 0.04175332, 0.03864555, 0.03571478, 0.03269915, 
    0.02984038, 0.02703318, 0.02474549, 0.0235727, 0.02260473, 0.02175616, 
    0.01968192, 0.01853958, 0.01825667, 0.01858922, 0.02152805, 0.02793169, 
    0.03618656, 0.03878286, 0.04819504, 0.05101745, 0.06652027, 0.08150315, 
    0.0961434, 0.07084978, 0.0497671, 0.03731534, 0.03326725, 0.03433823, 
    0.03472437, 0.02946474, 0.0276178, 0.02503158, 0.02219118, 0.01978667, 
    0.01889434, 0.01745579, 0.0162125, 0.01505942, 0.01512322, 0.01469036, 
    0.01459681, 0.02053429, 0.03211814, 0.03504532, 0.01840965, 0.01551427, 
    0.01528328, 0.01505197, 0.01405121, 0.01423585, 0.01509005, 0.01506049, 
    0.01500125, 0.01509749, 0.01519827, 0.01517837, 0.01589777, 0.01692957, 
    0.0178049, 0.01820548, 0.01897114, 0.02025549, 0.0207823, 0.02115879, 
    0.02187787, 0.0228803, 0.02382896, 0.02509996, 0.02558098, 0.02634498, 
    0.0273875, 0.0284514, 0.02875155, 0.02932919, 0.02919143, 0.02915357, 
    0.02781461, 0.02574988, 0.02266401, 0.01927338, 0.01525186, 0.01148103, 
    0.008436374, 0.006553261, 0.006012001, 0.005631275, 0.006080053, 
    0.006764134, 0.007065406, 0.006916829, 0.006645755, 0.006459266, 
    0.006446099, 0.006037058, 0.005453045, 0.005292657, 0.005172027, 
    0.005530572, 0.006101127, 0.006716309,
  0.006482502, 0.005856624, 0.005271276, 0.005342454, 0.005267369, 
    0.005090728, 0.004946326, 0.005148166, 0.005057677, 0.004475717, 
    0.004078032, 0.004385018, 0.006278505, 0.01134105, 0.01122047, 
    0.005783743, 0.004212447, 0.003493889, 0.003346328, 0.003296792, 
    0.003127742, 0.00310378, 0.003001576, 0.002733164, 0.002635605, 
    0.002575582, 0.003014797, 0.003909837, 0.004417506, 0.00678273, 
    0.007049358, 0.007618723, 0.009398847, 0.01312173, 0.01345367, 
    0.01353731, 0.01184887, 0.01132727, 0.01095043, 0.01082108, 0.01057722, 
    0.01010222, 0.009704815, 0.009486226, 0.009361508, 0.009867936, 0.010889, 
    0.01195346, 0.012733, 0.01438062, 0.01776037, 0.02264171, 0.02809866, 
    0.03343439, 0.03870047, 0.04576625, 0.05371612, 0.06327863, 0.09084318, 
    0.08515052, 0.08294441, 0.08799773, 0.08574666, 0.0884596, 0.08858822, 
    0.08043584, 0.07690392, 0.07067405, 0.06405876, 0.0533171, 0.04441018, 
    0.04001372, 0.04056064, 0.04713821, 0.06135855, 0.06565741, 0.06319264, 
    0.06962042, 0.06895236, 0.07891894, 0.08009713, 0.07646167, 0.07894669, 
    0.1070595, 0.1111868, 0.08696473, 0.07591901, 0.07366201, 0.07533359, 
    0.0643488, 0.06243263, 0.06459007, 0.0642117, 0.06360067, 0.0644533, 
    0.06437971, 0.06488286, 0.06607066, 0.06479692, 0.06184218, 0.05980521, 
    0.0606379, 0.06056314, 0.05952831, 0.05856892, 0.05814668, 0.05779451, 
    0.05574928, 0.05106479, 0.04766236, 0.04804677, 0.05037932, 0.05283817, 
    0.05189893, 0.0454793, 0.03977386, 0.03631324, 0.03334597, 0.03237103, 
    0.03203838, 0.03226648, 0.03314139, 0.03237737, 0.02895504, 0.02711754, 
    0.02587244, 0.0243297, 0.02468397, 0.02501604, 0.02437262, 0.02232928, 
    0.02106193, 0.02060015, 0.02037575, 0.02062208, 0.02117652, 0.02214121, 
    0.02335411, 0.02398971, 0.02303747, 0.02323479, 0.02390677, 0.02396804, 
    0.02351183, 0.02389625, 0.02391375, 0.0232365, 0.02298424, 0.02256046, 
    0.02266423, 0.02296414, 0.02285258, 0.02359517, 0.02380285, 0.02368135, 
    0.02480175, 0.02495234, 0.02455355, 0.02399927, 0.02308595, 0.02052762, 
    0.01754444, 0.01889786, 0.04399132, 0.03490548, 0.0286041, 0.02659954, 
    0.02469791, 0.0240936, 0.02471814, 0.02572318, 0.02758139, 0.03087534, 
    0.03353295, 0.03679387, 0.04053675, 0.0429817, 0.04431367, 0.04507616, 
    0.04600725, 0.04731342, 0.0479482, 0.04878477, 0.04886463, 0.04789739, 
    0.04613576, 0.04470126, 0.04256704, 0.04100615, 0.03810282, 0.03387903, 
    0.0304507, 0.02767835, 0.02474538, 0.02202523, 0.02053433, 0.01979425, 
    0.01976464, 0.01791896, 0.01594431, 0.01529086, 0.01601893, 0.02031877, 
    0.02946673, 0.03882503, 0.03941796, 0.04369613, 0.0534738, 0.08932906, 
    0.1029536, 0.0875651, 0.05899986, 0.03779502, 0.02975501, 0.02750646, 
    0.02916544, 0.03018882, 0.02738571, 0.0264942, 0.02517306, 0.02345793, 
    0.02146652, 0.02014598, 0.01796536, 0.01683946, 0.01732296, 0.02047032, 
    0.01995769, 0.01838855, 0.01804377, 0.02010041, 0.01990242, 0.01836594, 
    0.01711259, 0.01749518, 0.01650739, 0.01543539, 0.01584146, 0.01620441, 
    0.01604759, 0.01527713, 0.01513205, 0.01555216, 0.01570036, 0.01677544, 
    0.01794508, 0.01866801, 0.01862623, 0.01858822, 0.02014392, 0.02076034, 
    0.02107724, 0.02185441, 0.02263804, 0.02331249, 0.0249457, 0.02611293, 
    0.02692902, 0.02747577, 0.02741664, 0.02803102, 0.02908113, 0.02931383, 
    0.02855852, 0.02734773, 0.02553531, 0.02264287, 0.01944016, 0.01548604, 
    0.0120232, 0.008966418, 0.006618035, 0.005731559, 0.005497972, 
    0.005619586, 0.006239284, 0.006862614, 0.006677788, 0.00631662, 
    0.006239439, 0.006236044, 0.005797978, 0.005564927, 0.005391151, 
    0.004984442, 0.005154963, 0.005511205, 0.006434164,
  0.005577131, 0.005829426, 0.005688706, 0.005822959, 0.005971479, 
    0.005502129, 0.004912159, 0.005282627, 0.005584556, 0.004998461, 
    0.004733577, 0.004521281, 0.004544316, 0.007565636, 0.008030162, 
    0.004811887, 0.003670011, 0.003254551, 0.003290364, 0.003331782, 
    0.00314265, 0.003093463, 0.002957074, 0.002692109, 0.002636611, 
    0.002564004, 0.002852457, 0.003378658, 0.004365752, 0.006375618, 
    0.006945836, 0.007634068, 0.009526356, 0.01170245, 0.01176113, 
    0.01097625, 0.01069081, 0.01065684, 0.01084204, 0.01094727, 0.01090099, 
    0.01046457, 0.009752125, 0.009891099, 0.01025575, 0.01029529, 0.01048313, 
    0.01056896, 0.01073778, 0.01137485, 0.01320655, 0.01708573, 0.02217932, 
    0.02785538, 0.03435421, 0.04260736, 0.05076848, 0.05771851, 0.07432968, 
    0.07872461, 0.07760906, 0.08266608, 0.0790334, 0.07855423, 0.07574843, 
    0.07378852, 0.07126704, 0.0652772, 0.06071054, 0.05273477, 0.04160447, 
    0.03710376, 0.03909267, 0.04691305, 0.06267873, 0.05704729, 0.05793731, 
    0.06043471, 0.06286747, 0.07564782, 0.07637002, 0.08431598, 0.08666676, 
    0.10868, 0.1076158, 0.08509097, 0.08042751, 0.07878518, 0.07393236, 
    0.06963538, 0.07047258, 0.0699062, 0.06870954, 0.06842973, 0.06684329, 
    0.06353157, 0.06180261, 0.07071985, 0.06724633, 0.06384859, 0.06036063, 
    0.05940781, 0.05948266, 0.05957701, 0.05941902, 0.06016923, 0.06076251, 
    0.05950755, 0.05485146, 0.05118048, 0.05247082, 0.05387544, 0.05603058, 
    0.05488405, 0.04824323, 0.04188568, 0.03842558, 0.0352867, 0.03468961, 
    0.03467597, 0.03500618, 0.03623753, 0.03573525, 0.03185009, 0.02909242, 
    0.02789578, 0.02721845, 0.02760198, 0.0275449, 0.02529776, 0.02308861, 
    0.02245882, 0.02222329, 0.02267079, 0.02330882, 0.0234369, 0.02395166, 
    0.0244896, 0.02462571, 0.0243261, 0.02544345, 0.0259841, 0.02572969, 
    0.02533295, 0.02526516, 0.02604977, 0.02555071, 0.02512627, 0.02448229, 
    0.02364855, 0.02328097, 0.02233439, 0.02237759, 0.02273571, 0.02358338, 
    0.0254407, 0.02631042, 0.02579805, 0.02505793, 0.02463214, 0.02292764, 
    0.02109716, 0.02137196, 0.0274448, 0.02902823, 0.02821661, 0.02727048, 
    0.0249592, 0.02457375, 0.02558223, 0.02690248, 0.02876887, 0.03241229, 
    0.03506074, 0.0383862, 0.04188678, 0.04394599, 0.04466388, 0.04566617, 
    0.04622749, 0.04689841, 0.0476177, 0.0480223, 0.04819742, 0.04678395, 
    0.0446883, 0.04275167, 0.04053487, 0.03886549, 0.03639393, 0.03227878, 
    0.02840574, 0.0251366, 0.02240043, 0.02028603, 0.01847301, 0.0175545, 
    0.01733558, 0.01584753, 0.01405522, 0.01379266, 0.01417583, 0.02002054, 
    0.03326967, 0.0396668, 0.03415149, 0.03803774, 0.05806972, 0.1037917, 
    0.0880763, 0.06758151, 0.04810276, 0.03352451, 0.02776036, 0.02589431, 
    0.02642033, 0.02689392, 0.02654939, 0.02664704, 0.02520811, 0.02377685, 
    0.02226595, 0.02009167, 0.01796005, 0.01811012, 0.02290845, 0.02525747, 
    0.02330487, 0.0214151, 0.01938719, 0.01914225, 0.01887753, 0.01872776, 
    0.01845018, 0.01852399, 0.01788574, 0.01742458, 0.01812595, 0.01825888, 
    0.01741445, 0.01587368, 0.01542005, 0.01585049, 0.01602062, 0.01692407, 
    0.0184187, 0.01965867, 0.01918705, 0.01865076, 0.02025126, 0.02078648, 
    0.0213594, 0.02205504, 0.02259723, 0.02309441, 0.02465369, 0.0264003, 
    0.02722529, 0.02769142, 0.02737784, 0.02775369, 0.02851453, 0.02920859, 
    0.02911742, 0.02786988, 0.02623046, 0.02311265, 0.02002912, 0.01635789, 
    0.01262411, 0.009615386, 0.007204631, 0.005760004, 0.005356533, 
    0.005327039, 0.005483946, 0.006337774, 0.006394655, 0.006256515, 
    0.006260562, 0.006223667, 0.005982285, 0.005886313, 0.005796583, 
    0.005486269, 0.005433848, 0.005314053, 0.005539795,
  0.005110974, 0.005584119, 0.005935582, 0.006738926, 0.00778769, 
    0.006995469, 0.005747412, 0.005512585, 0.005095748, 0.004632665, 
    0.004841229, 0.004497759, 0.003791765, 0.004844537, 0.004916608, 
    0.00392067, 0.003479024, 0.00313364, 0.003136964, 0.003158533, 
    0.003003371, 0.003145556, 0.003133201, 0.002666894, 0.002588174, 
    0.002586426, 0.002669886, 0.003009994, 0.004445644, 0.006161698, 
    0.006880387, 0.008055441, 0.01080621, 0.01145072, 0.0105606, 0.01014002, 
    0.01072176, 0.01064356, 0.01098839, 0.01106919, 0.01085821, 0.01027104, 
    0.009474951, 0.009689223, 0.01003874, 0.009928222, 0.01001152, 
    0.01042624, 0.01010345, 0.01018846, 0.01125518, 0.01337477, 0.01713046, 
    0.02207902, 0.02764299, 0.03365242, 0.03989889, 0.04868915, 0.06296757, 
    0.06992196, 0.06861202, 0.06898309, 0.06813029, 0.06527262, 0.06457211, 
    0.06279363, 0.06203507, 0.05781692, 0.0557932, 0.05026239, 0.04205567, 
    0.03731587, 0.03982704, 0.0454948, 0.05255611, 0.05074007, 0.05499809, 
    0.05335294, 0.06205207, 0.06848888, 0.0740571, 0.08437283, 0.09753788, 
    0.1162404, 0.115696, 0.0974497, 0.09157578, 0.08722328, 0.08736347, 
    0.0905672, 0.08624226, 0.07764793, 0.0725606, 0.07256302, 0.07089254, 
    0.06372716, 0.06706207, 0.08395355, 0.07839529, 0.07067651, 0.06457488, 
    0.06217193, 0.06158967, 0.06145316, 0.06200935, 0.06212397, 0.06228761, 
    0.06182475, 0.05917902, 0.05639062, 0.05635537, 0.05705947, 0.05845433, 
    0.05595805, 0.04950226, 0.04558986, 0.04160998, 0.03835849, 0.03811352, 
    0.03783487, 0.03796947, 0.03822762, 0.03798646, 0.03566658, 0.03234406, 
    0.03122591, 0.03121569, 0.03112335, 0.03006405, 0.02785039, 0.02567652, 
    0.02481176, 0.02469356, 0.02556512, 0.02635291, 0.0261823, 0.02646612, 
    0.02701538, 0.02646262, 0.02656361, 0.02731218, 0.02700479, 0.02614179, 
    0.02614357, 0.02621922, 0.0268909, 0.02653529, 0.02626476, 0.02604689, 
    0.02477181, 0.02393603, 0.02296819, 0.02276674, 0.0229978, 0.02354921, 
    0.02521995, 0.02648476, 0.0269113, 0.02668933, 0.02576651, 0.02727048, 
    0.02618155, 0.0254223, 0.02642614, 0.02726343, 0.02795083, 0.02728129, 
    0.02580543, 0.02551855, 0.02687101, 0.02802647, 0.02989577, 0.03309073, 
    0.03557274, 0.03857412, 0.04118486, 0.04319575, 0.04458717, 0.04518428, 
    0.04550382, 0.04618539, 0.04722391, 0.04663714, 0.04694716, 0.04596035, 
    0.0436523, 0.04165232, 0.03916516, 0.03621383, 0.03320103, 0.02949818, 
    0.02654497, 0.0235622, 0.02059175, 0.01847687, 0.0167836, 0.01581462, 
    0.01550561, 0.01441514, 0.01292059, 0.0126906, 0.01448358, 0.02352865, 
    0.03534466, 0.03532613, 0.03176008, 0.03626277, 0.05490161, 0.08265818, 
    0.05686204, 0.05315127, 0.04408538, 0.03481406, 0.02994826, 0.02767108, 
    0.02752448, 0.02834857, 0.0290083, 0.02806681, 0.02570249, 0.02401173, 
    0.02341583, 0.02281473, 0.02370758, 0.02372846, 0.02447306, 0.02546744, 
    0.02468926, 0.02355162, 0.02235838, 0.02131436, 0.02075942, 0.02057038, 
    0.02072991, 0.02014791, 0.01920745, 0.01937883, 0.02006388, 0.01972394, 
    0.01837608, 0.01722334, 0.01624822, 0.01671367, 0.01649977, 0.01716168, 
    0.01855999, 0.02054522, 0.020441, 0.01989199, 0.02128796, 0.02166375, 
    0.02219076, 0.02282673, 0.02294927, 0.0231625, 0.02460404, 0.02589389, 
    0.02638218, 0.02666597, 0.02672767, 0.02763725, 0.02828555, 0.02879149, 
    0.02884701, 0.02820234, 0.02647009, 0.02387073, 0.02118416, 0.01777688, 
    0.0143098, 0.01090142, 0.007784249, 0.006104231, 0.005539815, 
    0.005229284, 0.005356162, 0.005907376, 0.006043451, 0.00604389, 
    0.00611303, 0.006238542, 0.006188889, 0.006150405, 0.005996175, 
    0.005669183, 0.005274488, 0.005046417, 0.005096803,
  0.004701533, 0.00522145, 0.005978662, 0.007083146, 0.009194633, 
    0.007896988, 0.006493421, 0.005347016, 0.00466193, 0.00455403, 
    0.004874784, 0.004564175, 0.004258334, 0.004637695, 0.004047523, 
    0.003782868, 0.003785474, 0.00349075, 0.003396915, 0.003259251, 
    0.002825754, 0.003137667, 0.003234246, 0.002747295, 0.002773207, 
    0.002511392, 0.002625864, 0.002606966, 0.00373804, 0.005703876, 
    0.00660191, 0.00754075, 0.01035082, 0.01164423, 0.01061252, 0.01060205, 
    0.01105959, 0.01076476, 0.01124313, 0.01140894, 0.01127511, 0.01087878, 
    0.01027767, 0.009885492, 0.008946015, 0.009160734, 0.01007342, 
    0.009798187, 0.009051833, 0.009555568, 0.01089316, 0.0118813, 0.01408213, 
    0.01727306, 0.02101896, 0.02517314, 0.0307137, 0.0391002, 0.05074848, 
    0.05281524, 0.05467172, 0.05528358, 0.0544201, 0.05302807, 0.04960857, 
    0.04802376, 0.0483612, 0.04829097, 0.04821342, 0.04517937, 0.03748034, 
    0.03407465, 0.03799772, 0.04562038, 0.04862718, 0.04833942, 0.0525893, 
    0.05389408, 0.06342432, 0.06878091, 0.07233997, 0.08075731, 0.09398723, 
    0.1100936, 0.1215727, 0.1058848, 0.1027096, 0.09740983, 0.09535264, 
    0.1029174, 0.1006479, 0.09239245, 0.08778685, 0.08121295, 0.07652501, 
    0.07435019, 0.08689091, 0.1325438, 0.09444562, 0.07554264, 0.06941944, 
    0.06682002, 0.06663127, 0.06480979, 0.06377716, 0.06421877, 0.06394491, 
    0.06316791, 0.0618785, 0.06010775, 0.05895537, 0.05830079, 0.05893753, 
    0.05710776, 0.0524856, 0.04930115, 0.04540782, 0.04251254, 0.04238652, 
    0.04138527, 0.0409551, 0.04009757, 0.03918458, 0.03874706, 0.03712513, 
    0.03580621, 0.03475032, 0.03415424, 0.03237911, 0.03017989, 0.02869421, 
    0.02804535, 0.0278181, 0.02790915, 0.02822678, 0.02845215, 0.02856151, 
    0.02923056, 0.02857065, 0.02827086, 0.0282987, 0.0279274, 0.02772589, 
    0.02725346, 0.02738885, 0.02798574, 0.02771517, 0.02762522, 0.02765914, 
    0.02690667, 0.02616758, 0.02527298, 0.02508602, 0.02479309, 0.02455766, 
    0.02568659, 0.02670938, 0.02774147, 0.02896298, 0.02904995, 0.02942551, 
    0.02849455, 0.02772223, 0.02802636, 0.02832712, 0.02839313, 0.02779911, 
    0.02728844, 0.02737303, 0.02805728, 0.02909204, 0.03050262, 0.03307957, 
    0.03534335, 0.03739, 0.0389052, 0.04097648, 0.04289102, 0.04439405, 
    0.0446694, 0.04475732, 0.04521149, 0.04535009, 0.04533327, 0.04476097, 
    0.04303604, 0.04043216, 0.03740494, 0.03398356, 0.03068502, 0.02751154, 
    0.02468619, 0.02222481, 0.01968109, 0.01727744, 0.01508864, 0.01369199, 
    0.01362973, 0.0131061, 0.0115678, 0.01257661, 0.01808636, 0.0285795, 
    0.03468908, 0.03063181, 0.0279131, 0.03012703, 0.04445088, 0.06123623, 
    0.05346398, 0.05164605, 0.04559713, 0.03774104, 0.0340552, 0.03284527, 
    0.0321098, 0.03204455, 0.03256707, 0.03193578, 0.03030377, 0.0286674, 
    0.02757307, 0.02650432, 0.0265091, 0.02584512, 0.02538393, 0.02730186, 
    0.02775932, 0.02742126, 0.02604218, 0.02504039, 0.02421867, 0.02352151, 
    0.02407126, 0.02349823, 0.02241448, 0.02218809, 0.02232125, 0.02135028, 
    0.01991795, 0.01906299, 0.01804393, 0.01803185, 0.01776366, 0.01837281, 
    0.01958863, 0.02108552, 0.02142168, 0.02086573, 0.02170376, 0.02260611, 
    0.02333373, 0.02432005, 0.02413952, 0.02406486, 0.02477726, 0.02540632, 
    0.02510656, 0.0258977, 0.02646005, 0.02720001, 0.02790216, 0.02826789, 
    0.02815324, 0.02848218, 0.02748602, 0.02540386, 0.02284738, 0.01973256, 
    0.01663901, 0.01309914, 0.009265475, 0.00669234, 0.005661954, 
    0.005235418, 0.005267352, 0.005722439, 0.005878287, 0.00587987, 
    0.00586232, 0.006015576, 0.00618666, 0.006219709, 0.005891598, 
    0.005558941, 0.004884411, 0.004439153, 0.004536897,
  0.004374793, 0.005236113, 0.005837959, 0.006478593, 0.007365518, 
    0.006647445, 0.005910256, 0.005222934, 0.005085688, 0.00496728, 
    0.005116644, 0.004835745, 0.004379354, 0.004354406, 0.004046763, 
    0.003791228, 0.00396501, 0.003898834, 0.003779553, 0.003390394, 
    0.002875761, 0.003042647, 0.003114422, 0.002937441, 0.002949693, 
    0.002545106, 0.002928772, 0.00276627, 0.004326764, 0.005560109, 
    0.006733367, 0.007943166, 0.009313837, 0.01093687, 0.01109022, 
    0.01156817, 0.01182138, 0.01174826, 0.01156333, 0.01192601, 0.01216341, 
    0.01199154, 0.01163447, 0.01101758, 0.009519402, 0.01054055, 0.01075385, 
    0.009413969, 0.009038404, 0.01087947, 0.01308032, 0.01348491, 0.01372874, 
    0.01479023, 0.01462808, 0.01714663, 0.02229314, 0.03034891, 0.03772775, 
    0.03897291, 0.03914368, 0.04047237, 0.04055306, 0.04138229, 0.03937301, 
    0.03897712, 0.03905444, 0.04004924, 0.0403542, 0.03839506, 0.03707472, 
    0.03740053, 0.04232617, 0.05074687, 0.04918407, 0.04920008, 0.05523543, 
    0.06491192, 0.07719156, 0.06941175, 0.06678902, 0.07235943, 0.08063527, 
    0.09407004, 0.1021353, 0.1097171, 0.1146249, 0.1090003, 0.1093301, 
    0.1140747, 0.1154011, 0.1037552, 0.09982604, 0.09612308, 0.0906459, 
    0.09487662, 0.1189703, 0.2035925, 0.09994572, 0.08070118, 0.07526029, 
    0.07058164, 0.07064672, 0.06873322, 0.06678773, 0.06740713, 0.06768167, 
    0.06608545, 0.06452153, 0.06203562, 0.0609583, 0.06116968, 0.06093962, 
    0.05828242, 0.05493049, 0.05263942, 0.05012074, 0.04766294, 0.04672358, 
    0.04475557, 0.0433799, 0.04245324, 0.04202794, 0.04259785, 0.04241018, 
    0.04102445, 0.03939132, 0.03791154, 0.03537741, 0.03293893, 0.0314467, 
    0.03121039, 0.03095851, 0.03075589, 0.03061011, 0.03093431, 0.03072059, 
    0.03064917, 0.03016213, 0.02984948, 0.02952404, 0.02941895, 0.02927242, 
    0.0282704, 0.02835369, 0.02926728, 0.02909196, 0.02913919, 0.02897245, 
    0.0288079, 0.02836065, 0.02769922, 0.02764621, 0.0272957, 0.02679115, 
    0.02706487, 0.02751717, 0.02874803, 0.03102697, 0.03192148, 0.03213919, 
    0.03132984, 0.03033735, 0.03017752, 0.03039915, 0.02988604, 0.02922514, 
    0.02876965, 0.02899277, 0.0299094, 0.0302798, 0.03055918, 0.0325537, 
    0.03443649, 0.03630346, 0.03790117, 0.0397189, 0.04148097, 0.04319801, 
    0.04415523, 0.04389976, 0.04361618, 0.04383748, 0.04409703, 0.04346815, 
    0.0413163, 0.03852688, 0.03544191, 0.03189069, 0.0286029, 0.02590288, 
    0.02305872, 0.02076905, 0.01825815, 0.01593909, 0.01366675, 0.01161902, 
    0.01160213, 0.01094674, 0.01058671, 0.01390538, 0.02219702, 0.03139329, 
    0.02663147, 0.0257361, 0.02610564, 0.02534528, 0.03310378, 0.05439693, 
    0.05201445, 0.05239557, 0.04871986, 0.04205787, 0.03868239, 0.03747412, 
    0.03749299, 0.03723905, 0.03751997, 0.03683752, 0.03579234, 0.03314576, 
    0.02955786, 0.02637855, 0.02731581, 0.02875821, 0.02868652, 0.03074371, 
    0.03125504, 0.03167841, 0.03030427, 0.02849999, 0.0277868, 0.0274436, 
    0.02729478, 0.02662825, 0.02596162, 0.02578112, 0.0248718, 0.02354017, 
    0.0222581, 0.02163424, 0.02051674, 0.02004165, 0.02044039, 0.0209052, 
    0.02111141, 0.02220492, 0.02306085, 0.02300834, 0.02327276, 0.02353932, 
    0.02455123, 0.02556102, 0.02539437, 0.02565184, 0.0249476, 0.02447503, 
    0.02467108, 0.02542445, 0.02629921, 0.02697108, 0.02772246, 0.02807799, 
    0.02820721, 0.02852717, 0.02781607, 0.02645377, 0.02448326, 0.0217831, 
    0.0190811, 0.01596572, 0.01184298, 0.008473864, 0.006353809, 0.005609111, 
    0.005351274, 0.005487817, 0.005570605, 0.005608016, 0.005434653, 
    0.005559151, 0.005753845, 0.006075595, 0.006127478, 0.005601659, 
    0.0049066, 0.004206383, 0.004090093,
  0.00412516, 0.0047222, 0.005252996, 0.005736971, 0.006197338, 0.005761692, 
    0.006218825, 0.005848489, 0.005566641, 0.00482873, 0.004967267, 
    0.004907584, 0.004534937, 0.004661199, 0.004532898, 0.004291299, 
    0.004156809, 0.003966182, 0.003810664, 0.003638353, 0.003284023, 
    0.003121496, 0.003164396, 0.003079759, 0.003033631, 0.003014712, 
    0.003018887, 0.0032011, 0.005371904, 0.005587876, 0.006365112, 
    0.008351498, 0.009782528, 0.01092606, 0.01147917, 0.012126, 0.01230601, 
    0.01237919, 0.01249997, 0.01268192, 0.01318179, 0.01322613, 0.01361493, 
    0.013464, 0.01243761, 0.01225617, 0.01152683, 0.01187926, 0.01177842, 
    0.01259064, 0.01310829, 0.01393085, 0.01378484, 0.01277335, 0.01031365, 
    0.01205574, 0.01573105, 0.02001789, 0.02517577, 0.02799357, 0.030673, 
    0.03041508, 0.03055784, 0.03234534, 0.03370387, 0.0340289, 0.03429071, 
    0.03655442, 0.04349421, 0.05237675, 0.05994221, 0.06185523, 0.0624513, 
    0.06506922, 0.0579756, 0.05137278, 0.06033604, 0.07880834, 0.09126364, 
    0.07610301, 0.06308387, 0.06635184, 0.07668863, 0.09444031, 0.1073625, 
    0.1103822, 0.122867, 0.1166747, 0.1210117, 0.1293526, 0.1159652, 
    0.1149126, 0.1051202, 0.1029272, 0.1143728, 0.1249351, 0.1366475, 
    0.1361341, 0.09964421, 0.08808726, 0.08210585, 0.07704697, 0.07609317, 
    0.07417639, 0.07232088, 0.07386303, 0.07302125, 0.07053696, 0.06835588, 
    0.06497912, 0.0618596, 0.06246863, 0.06293088, 0.06092873, 0.05886335, 
    0.05634837, 0.05502212, 0.05355621, 0.05174765, 0.04879487, 0.04753052, 
    0.04748103, 0.04745128, 0.04770574, 0.04785838, 0.04677531, 0.04463176, 
    0.04228141, 0.03985465, 0.03741556, 0.03502103, 0.03418865, 0.03469003, 
    0.03455626, 0.03399155, 0.03426334, 0.03400057, 0.03282827, 0.03224583, 
    0.03170925, 0.03103936, 0.03124552, 0.03119239, 0.03010027, 0.02959113, 
    0.03053199, 0.03090308, 0.03088622, 0.03070157, 0.03058787, 0.03106786, 
    0.03101288, 0.03157119, 0.0310419, 0.03017163, 0.02986076, 0.02956362, 
    0.03062781, 0.03288165, 0.03486571, 0.03473249, 0.03368248, 0.0326224, 
    0.03183243, 0.03170652, 0.03157426, 0.03160075, 0.03163816, 0.03181495, 
    0.0322908, 0.03203779, 0.03190516, 0.03350472, 0.03427884, 0.03592917, 
    0.03793016, 0.03986317, 0.04101191, 0.04275972, 0.04367658, 0.04340111, 
    0.04325703, 0.04300863, 0.04309093, 0.04215518, 0.03953837, 0.03675421, 
    0.0334757, 0.02996342, 0.02639026, 0.02391289, 0.0214919, 0.01917803, 
    0.01644575, 0.01423897, 0.01252815, 0.01039201, 0.009345421, 0.008923097, 
    0.01098622, 0.01727158, 0.02459079, 0.0258252, 0.02485136, 0.02275147, 
    0.02295997, 0.02102102, 0.03501914, 0.05232519, 0.04846537, 0.05113087, 
    0.05025355, 0.04510345, 0.04254676, 0.042181, 0.04257053, 0.0430864, 
    0.04346341, 0.04201435, 0.04000939, 0.03600149, 0.03070047, 0.02807592, 
    0.03101617, 0.03261193, 0.032269, 0.03350957, 0.03454275, 0.03620869, 
    0.03488206, 0.03253283, 0.03142868, 0.03111348, 0.03127817, 0.03093664, 
    0.02984368, 0.02856948, 0.02743594, 0.02659439, 0.02528552, 0.02410159, 
    0.02288165, 0.02257274, 0.02308754, 0.02359127, 0.02348561, 0.02355463, 
    0.02414978, 0.02497326, 0.02616578, 0.02615036, 0.0263327, 0.02727521, 
    0.02694867, 0.02623558, 0.02466394, 0.02404906, 0.02443775, 0.02565111, 
    0.02629106, 0.02657373, 0.02704025, 0.02756131, 0.02837642, 0.02849519, 
    0.02758017, 0.02670584, 0.02559403, 0.02339929, 0.02123833, 0.01928619, 
    0.01559514, 0.01178921, 0.00842404, 0.006549931, 0.006212148, 
    0.005935048, 0.005453953, 0.005435387, 0.004965233, 0.005054217, 
    0.005121383, 0.005666658, 0.006282273, 0.006106319, 0.005152132, 
    0.00427773, 0.003826821,
  0.003769948, 0.003995621, 0.004351347, 0.004721058, 0.005041978, 
    0.005128209, 0.005402307, 0.005421722, 0.004955616, 0.004678086, 
    0.005116433, 0.004860812, 0.004669376, 0.004851955, 0.004979401, 
    0.004841138, 0.004428506, 0.004040421, 0.00380694, 0.003858186, 
    0.003594076, 0.003392414, 0.003324511, 0.003162368, 0.003575483, 
    0.0035152, 0.002804033, 0.004562581, 0.005609964, 0.005432939, 
    0.006452426, 0.008039315, 0.009606568, 0.01100072, 0.01193619, 
    0.01226865, 0.01220976, 0.01226088, 0.01303623, 0.01312216, 0.01370379, 
    0.01533121, 0.01564917, 0.01540794, 0.01512618, 0.01359695, 0.01433578, 
    0.01513304, 0.01505286, 0.0143253, 0.01256586, 0.0125576, 0.0129713, 
    0.01104461, 0.009459231, 0.009300572, 0.0113657, 0.0149327, 0.01922887, 
    0.02309117, 0.02566653, 0.02701795, 0.02723716, 0.02807944, 0.03018155, 
    0.03368044, 0.04087611, 0.05194733, 0.05987344, 0.07323229, 0.09321098, 
    0.1071598, 0.1090612, 0.1014983, 0.08181464, 0.07076734, 0.07578514, 
    0.1098836, 0.09978341, 0.08221541, 0.06036977, 0.06676429, 0.07232782, 
    0.09263557, 0.1122954, 0.1109973, 0.1205287, 0.1199, 0.1280047, 
    0.1293656, 0.1210016, 0.1144593, 0.1111572, 0.1078598, 0.1094467, 
    0.1256666, 0.1314922, 0.1248586, 0.1059547, 0.09683167, 0.08989698, 
    0.08649332, 0.08514061, 0.08284003, 0.08045086, 0.08094423, 0.08060708, 
    0.07764585, 0.07422087, 0.07075761, 0.06716881, 0.06550524, 0.06544553, 
    0.0646929, 0.06411491, 0.06193881, 0.06067535, 0.05994346, 0.05766948, 
    0.05392256, 0.05262041, 0.05266556, 0.0527289, 0.05187374, 0.0524802, 
    0.05211, 0.04949845, 0.04695639, 0.04444886, 0.04201217, 0.03987207, 
    0.038404, 0.03890655, 0.03917075, 0.03862917, 0.03885146, 0.03859312, 
    0.03673898, 0.03492829, 0.0333791, 0.0329727, 0.03349417, 0.0337985, 
    0.03324926, 0.03280565, 0.03355822, 0.03352131, 0.03302119, 0.03308453, 
    0.03303305, 0.03348975, 0.03509204, 0.03618887, 0.03529228, 0.0348072, 
    0.03464409, 0.03427474, 0.03439604, 0.03571423, 0.03783644, 0.03727709, 
    0.03631608, 0.0353574, 0.03402269, 0.03321148, 0.03345423, 0.03425086, 
    0.03460574, 0.0342392, 0.03462021, 0.03443302, 0.03422565, 0.03491802, 
    0.03606633, 0.03660455, 0.03735818, 0.03970106, 0.04116622, 0.04268852, 
    0.04388597, 0.04413727, 0.04340231, 0.04272053, 0.04159998, 0.03995056, 
    0.03774827, 0.03504349, 0.03190528, 0.02826761, 0.02464703, 0.02216104, 
    0.01988167, 0.01757233, 0.01490182, 0.01261075, 0.01148826, 0.009405945, 
    0.007418511, 0.00790707, 0.01220724, 0.01928237, 0.02451148, 0.02673304, 
    0.02065095, 0.02252254, 0.01984123, 0.02468524, 0.042874, 0.04391947, 
    0.04224126, 0.04753492, 0.050244, 0.04765086, 0.04601295, 0.0463451, 
    0.04722922, 0.04799921, 0.04760492, 0.04616738, 0.04327381, 0.03975746, 
    0.03503239, 0.03437326, 0.0377695, 0.03786585, 0.03625091, 0.03588755, 
    0.03712056, 0.03922439, 0.03891563, 0.03692879, 0.03555453, 0.03577012, 
    0.03565289, 0.03573382, 0.03465336, 0.03244006, 0.03121253, 0.03115173, 
    0.02985373, 0.02816144, 0.0264573, 0.02580409, 0.02533159, 0.02595492, 
    0.02562501, 0.02493849, 0.02540203, 0.02665856, 0.02834676, 0.028608, 
    0.02879796, 0.02935681, 0.02868857, 0.02791473, 0.02667058, 0.02558836, 
    0.02562214, 0.02646378, 0.0269652, 0.02658715, 0.0270975, 0.02739754, 
    0.0284024, 0.02882095, 0.02811223, 0.02739409, 0.02620215, 0.02447646, 
    0.02259549, 0.02124678, 0.01868958, 0.01581192, 0.01171541, 0.008218327, 
    0.007544251, 0.007723886, 0.007044368, 0.006814868, 0.006044919, 
    0.005126776, 0.004906324, 0.005189889, 0.005815879, 0.00609007, 
    0.005497498, 0.004653995, 0.003950988,
  0.003651618, 0.003727021, 0.004154443, 0.004482444, 0.004897554, 
    0.004980606, 0.004834104, 0.004908749, 0.004737942, 0.004991498, 
    0.005397819, 0.005170973, 0.005100745, 0.00574503, 0.005789613, 
    0.005271467, 0.004859832, 0.004500946, 0.004184469, 0.004019404, 
    0.003958563, 0.003962947, 0.00380964, 0.003641072, 0.004424067, 
    0.004117721, 0.00373383, 0.005424477, 0.004831088, 0.005792529, 
    0.00636083, 0.007663541, 0.00922164, 0.01045784, 0.01159378, 0.01241208, 
    0.01230632, 0.01174877, 0.01220464, 0.01278366, 0.01473835, 0.01670171, 
    0.01706061, 0.01652379, 0.01718551, 0.01657417, 0.01442986, 0.0140549, 
    0.01536323, 0.01338535, 0.01141169, 0.01149731, 0.01318989, 0.01319269, 
    0.01237451, 0.009785061, 0.01011907, 0.01231645, 0.01572572, 0.01971033, 
    0.02313931, 0.02690764, 0.02861484, 0.03017326, 0.03786948, 0.04331453, 
    0.05415044, 0.06515238, 0.071738, 0.09310758, 0.1200619, 0.1335538, 
    0.1300134, 0.1343707, 0.1600647, 0.1567213, 0.1128582, 0.1247252, 
    0.1304356, 0.09248017, 0.06725904, 0.07540544, 0.09316947, 0.1232897, 
    0.1286953, 0.113342, 0.1205159, 0.1225235, 0.1282275, 0.1377092, 
    0.1232194, 0.1123455, 0.1119568, 0.1122853, 0.1073319, 0.1316329, 
    0.1308393, 0.1214072, 0.1098122, 0.1022209, 0.09606105, 0.09559623, 
    0.09671097, 0.09488017, 0.09123932, 0.08845142, 0.08608142, 0.08440244, 
    0.08105737, 0.07776784, 0.07475739, 0.07305181, 0.07226212, 0.07088423, 
    0.06855693, 0.06699181, 0.06594766, 0.06536313, 0.0633906, 0.06035182, 
    0.05909224, 0.05913207, 0.05872625, 0.05801146, 0.05748376, 0.05703418, 
    0.05465395, 0.05169531, 0.04881158, 0.04679512, 0.0457847, 0.04506212, 
    0.04500403, 0.04496541, 0.04452052, 0.04429059, 0.04335849, 0.04175039, 
    0.03982151, 0.0378224, 0.03738341, 0.03799255, 0.03771679, 0.03711646, 
    0.03674928, 0.03724704, 0.03737195, 0.03682052, 0.03671409, 0.03651102, 
    0.03728426, 0.03916997, 0.03991624, 0.03907449, 0.03911308, 0.03959481, 
    0.03975502, 0.03979128, 0.04072126, 0.0422387, 0.04097633, 0.03944801, 
    0.03907058, 0.03768712, 0.03611444, 0.03578194, 0.03705066, 0.03709189, 
    0.036368, 0.0360113, 0.036479, 0.03640053, 0.03609205, 0.03717089, 
    0.03823107, 0.03844742, 0.03961929, 0.04127324, 0.0428677, 0.04375963, 
    0.04435538, 0.04433431, 0.04271625, 0.04062483, 0.03865733, 0.03654943, 
    0.03365992, 0.03078256, 0.02795996, 0.02436732, 0.0213713, 0.01894516, 
    0.01636686, 0.01360032, 0.01161526, 0.0105082, 0.008036006, 0.006819515, 
    0.008995933, 0.01354132, 0.01923263, 0.02269311, 0.02107067, 0.02057876, 
    0.01909794, 0.01855347, 0.03070363, 0.03968889, 0.03902657, 0.0402956, 
    0.04640249, 0.04937446, 0.04934725, 0.04947841, 0.04985484, 0.04981102, 
    0.05024798, 0.04917083, 0.04691059, 0.04398202, 0.04241655, 0.04013795, 
    0.04297632, 0.04552556, 0.04515838, 0.04238943, 0.04089464, 0.04153362, 
    0.04287938, 0.04326718, 0.04236625, 0.04082103, 0.04065667, 0.04101949, 
    0.04062932, 0.03931952, 0.03750842, 0.03673391, 0.03698979, 0.03562637, 
    0.03362042, 0.03104264, 0.02950604, 0.0282492, 0.02779818, 0.02790789, 
    0.02707037, 0.02740222, 0.02873369, 0.02959408, 0.02926478, 0.02997555, 
    0.03108247, 0.02996938, 0.02921302, 0.02837919, 0.02785977, 0.02774375, 
    0.027937, 0.02772527, 0.02713897, 0.02685922, 0.02717695, 0.02841788, 
    0.02916202, 0.02875702, 0.02822326, 0.02739377, 0.02597998, 0.02429508, 
    0.02283093, 0.02101379, 0.0188563, 0.01313139, 0.008057855, 0.008196671, 
    0.009432735, 0.01051962, 0.0119355, 0.01046625, 0.006505662, 0.00515838, 
    0.005023406, 0.005242244, 0.0053321, 0.005136999, 0.004525273, 0.003913922,
  0.003999753, 0.004046967, 0.004285935, 0.004667906, 0.004978556, 
    0.004954003, 0.004974904, 0.005353593, 0.005565025, 0.005797094, 
    0.006299602, 0.006741091, 0.007055648, 0.00727181, 0.006657801, 
    0.005892084, 0.005541586, 0.005339833, 0.00495251, 0.004689439, 
    0.004572522, 0.004624715, 0.004563767, 0.004425234, 0.005147939, 
    0.005226662, 0.006025321, 0.005925218, 0.005457669, 0.006552892, 
    0.007465504, 0.008172153, 0.00947174, 0.01050791, 0.01111939, 0.01210862, 
    0.01232889, 0.01194553, 0.01267103, 0.01455616, 0.01750144, 0.01940428, 
    0.01858128, 0.01756032, 0.01829314, 0.0218639, 0.01692929, 0.01470057, 
    0.0143104, 0.01221584, 0.0121113, 0.01145416, 0.01256741, 0.0151966, 
    0.01543826, 0.01119012, 0.0106454, 0.0119958, 0.01458928, 0.0184509, 
    0.02219061, 0.02867866, 0.03501729, 0.04411468, 0.0583897, 0.06561161, 
    0.0815855, 0.1031809, 0.09404176, 0.06551349, 0.05575763, 0.06168977, 
    0.06830671, 0.08501939, 0.1364366, 0.222153, 0.1762915, 0.1568734, 
    0.1166439, 0.08302768, 0.06318223, 0.09141596, 0.1413706, 0.1735282, 
    0.13787, 0.113127, 0.1237874, 0.1263209, 0.1223857, 0.1280892, 0.1151584, 
    0.1075244, 0.1126852, 0.1138872, 0.1082832, 0.118077, 0.1288985, 
    0.1160975, 0.1087205, 0.1037697, 0.09828868, 0.09920492, 0.1022861, 
    0.1033057, 0.10042, 0.09609911, 0.09330947, 0.09043952, 0.08637583, 
    0.08262651, 0.08035972, 0.07966376, 0.08058865, 0.08042175, 0.07719225, 
    0.07365161, 0.07218159, 0.07084275, 0.06908344, 0.06723817, 0.06595116, 
    0.06535121, 0.06498586, 0.06399518, 0.062773, 0.06252892, 0.06126783, 
    0.05797765, 0.05439056, 0.05277168, 0.05235641, 0.0518908, 0.05158226, 
    0.05112211, 0.05094688, 0.05055727, 0.04931863, 0.04836604, 0.04691427, 
    0.04494785, 0.04396297, 0.0433111, 0.04274733, 0.0421116, 0.04192881, 
    0.04227152, 0.04214872, 0.04154299, 0.04166448, 0.04126729, 0.04199892, 
    0.04335511, 0.04360773, 0.04198224, 0.04281297, 0.04418123, 0.04501742, 
    0.04610132, 0.0471962, 0.04802677, 0.04605827, 0.04399975, 0.04369185, 
    0.04293696, 0.04059051, 0.03880912, 0.03965032, 0.03989167, 0.03871246, 
    0.03843656, 0.03786851, 0.03715349, 0.03788646, 0.03861061, 0.03970812, 
    0.04026145, 0.04052947, 0.0416711, 0.04316225, 0.04348052, 0.0437629, 
    0.04442982, 0.04329201, 0.04125163, 0.03873434, 0.03687301, 0.03376127, 
    0.03064461, 0.02818878, 0.02497323, 0.0214204, 0.01872884, 0.01616542, 
    0.01341244, 0.01180321, 0.009255136, 0.006804896, 0.007508174, 
    0.01035556, 0.0138281, 0.01842065, 0.0212074, 0.01911051, 0.02004156, 
    0.01791105, 0.01910352, 0.03231913, 0.03843586, 0.03780235, 0.04101038, 
    0.04597111, 0.0486099, 0.05036793, 0.05225606, 0.05236929, 0.05171407, 
    0.05134647, 0.04999967, 0.04797725, 0.04573825, 0.04508527, 0.04508395, 
    0.04994645, 0.05250742, 0.0521529, 0.04867113, 0.04674463, 0.04700726, 
    0.04777006, 0.04827731, 0.04840811, 0.04753013, 0.04612449, 0.04607064, 
    0.04577935, 0.04532856, 0.0438753, 0.04363128, 0.0435369, 0.04114017, 
    0.03836474, 0.03542342, 0.03351196, 0.032066, 0.03100318, 0.03209012, 
    0.03161993, 0.03126993, 0.03241142, 0.03186553, 0.03075612, 0.0309947, 
    0.03199952, 0.03177294, 0.03108247, 0.03042004, 0.0301897, 0.02997126, 
    0.02976197, 0.02969551, 0.02927194, 0.02861824, 0.02827104, 0.02872289, 
    0.02901248, 0.02873688, 0.02824814, 0.02751924, 0.02704594, 0.02628656, 
    0.02504916, 0.02375276, 0.0216721, 0.01601096, 0.0128317, 0.01304721, 
    0.01164067, 0.01230299, 0.01287381, 0.01249943, 0.008749961, 0.00607443, 
    0.005148184, 0.004818873, 0.004796295, 0.004710414, 0.004419427, 
    0.004105396,
  0.00456723, 0.004470623, 0.004704718, 0.004808228, 0.0049192, 0.005190399, 
    0.005769289, 0.006341211, 0.006742009, 0.006936071, 0.007695673, 
    0.008559275, 0.00920009, 0.009028884, 0.008443143, 0.008242271, 
    0.007451307, 0.006451292, 0.005983905, 0.005757787, 0.005376271, 
    0.005344043, 0.005221069, 0.005444761, 0.006538914, 0.008005723, 
    0.009546283, 0.01050705, 0.009782151, 0.007954516, 0.009016618, 
    0.008550731, 0.009365267, 0.01031684, 0.01082954, 0.01152457, 0.01246511, 
    0.01328847, 0.01502138, 0.0187507, 0.0210739, 0.02347635, 0.02018444, 
    0.01525281, 0.01684171, 0.01603023, 0.01460629, 0.01364864, 0.01097793, 
    0.01223465, 0.01209733, 0.01255629, 0.01382227, 0.01579391, 0.01569449, 
    0.01303598, 0.01280724, 0.01288218, 0.01478816, 0.01921702, 0.02523014, 
    0.03576012, 0.04628357, 0.06158032, 0.0854648, 0.08186582, 0.06315645, 
    0.04507371, 0.035053, 0.02833806, 0.0273349, 0.03010853, 0.03234613, 
    0.03845667, 0.06505229, 0.1308658, 0.1416631, 0.08743163, 0.05572136, 
    0.05194442, 0.05130345, 0.08048445, 0.1828022, 0.1495156, 0.1031618, 
    0.1087637, 0.1109796, 0.1156024, 0.1225082, 0.1212497, 0.1076191, 
    0.1059387, 0.1069317, 0.1049418, 0.109813, 0.1187788, 0.1216242, 
    0.113866, 0.1053122, 0.1009451, 0.09598147, 0.09905657, 0.1028916, 
    0.1035024, 0.10127, 0.09870154, 0.0977359, 0.09569173, 0.09045974, 
    0.08705372, 0.08532589, 0.08451596, 0.08558063, 0.08643753, 0.08469531, 
    0.08167456, 0.07960629, 0.07827614, 0.07617553, 0.07348856, 0.07210211, 
    0.07171968, 0.07135394, 0.07012799, 0.06831799, 0.06772804, 0.06859841, 
    0.06567325, 0.06176001, 0.05984366, 0.05955232, 0.06041202, 0.06062594, 
    0.0589046, 0.05739286, 0.05693683, 0.05636368, 0.05497339, 0.05417675, 
    0.05248075, 0.05119725, 0.04947541, 0.04834718, 0.04768557, 0.04777955, 
    0.04809373, 0.04827296, 0.04738834, 0.04757139, 0.04770103, 0.04800613, 
    0.04822023, 0.04835872, 0.04716532, 0.04717254, 0.04829999, 0.04987386, 
    0.05131606, 0.05272183, 0.05280253, 0.05108734, 0.04856716, 0.04702711, 
    0.04742487, 0.04623984, 0.04397396, 0.0432495, 0.04334462, 0.0419441, 
    0.04144816, 0.04027111, 0.03902546, 0.03903674, 0.04053419, 0.04148072, 
    0.04241797, 0.04236534, 0.04278236, 0.04339611, 0.04391731, 0.04410691, 
    0.04396394, 0.0434681, 0.04220676, 0.03961596, 0.03700234, 0.03395956, 
    0.03113852, 0.0278813, 0.02499093, 0.0219159, 0.01927233, 0.0167996, 
    0.01538054, 0.01242369, 0.007485864, 0.006745988, 0.008948452, 
    0.01106455, 0.01421732, 0.01799095, 0.01747761, 0.01565376, 0.0173093, 
    0.01630105, 0.01899812, 0.02821712, 0.0345432, 0.03805256, 0.0440464, 
    0.04828206, 0.05159786, 0.05384694, 0.0554499, 0.05627696, 0.05649981, 
    0.05466823, 0.05281933, 0.05180693, 0.05022702, 0.04912437, 0.05105353, 
    0.0557515, 0.05786971, 0.05697883, 0.05539346, 0.05333447, 0.05292209, 
    0.05203972, 0.05195732, 0.05218908, 0.05104903, 0.05010973, 0.04979273, 
    0.05076659, 0.05083923, 0.04944406, 0.04988431, 0.05020396, 0.04805745, 
    0.04452615, 0.04010198, 0.03798476, 0.03635469, 0.03528952, 0.03661613, 
    0.03697492, 0.03793886, 0.03760282, 0.03505485, 0.03360918, 0.03235547, 
    0.03280457, 0.0336665, 0.03309725, 0.03224537, 0.03195652, 0.03214814, 
    0.03182449, 0.03141607, 0.03136152, 0.03074783, 0.02992181, 0.02982472, 
    0.02965774, 0.02933498, 0.02880468, 0.02875878, 0.02898416, 0.02790781, 
    0.02682157, 0.02557944, 0.02412375, 0.02119567, 0.01821455, 0.01694724, 
    0.0139698, 0.01226917, 0.01236389, 0.01184909, 0.01062657, 0.008685664, 
    0.006650997, 0.005697876, 0.005092919, 0.004865486, 0.004906424, 
    0.004857294,
  0.005785842, 0.005549765, 0.005825224, 0.005679201, 0.005470953, 
    0.00589817, 0.006638296, 0.007325258, 0.007717925, 0.008588697, 
    0.009770332, 0.01023899, 0.01046347, 0.01113347, 0.01139841, 0.01184921, 
    0.01000969, 0.008110809, 0.007364359, 0.006938488, 0.007212041, 
    0.007928261, 0.008235509, 0.008756152, 0.009403445, 0.01058058, 
    0.01331358, 0.01661365, 0.01613976, 0.01154835, 0.01013084, 0.009107797, 
    0.009106358, 0.01007056, 0.01042743, 0.01176458, 0.01325002, 0.01496128, 
    0.01909784, 0.02296244, 0.02963564, 0.02755267, 0.01497992, 0.01252295, 
    0.01182728, 0.01215023, 0.0159928, 0.01277937, 0.01135336, 0.01311973, 
    0.01284994, 0.01369714, 0.01507195, 0.01889828, 0.01589349, 0.01684562, 
    0.01714903, 0.01459298, 0.01571487, 0.02245049, 0.03425323, 0.04918133, 
    0.06264174, 0.07433187, 0.06346318, 0.04466917, 0.02605646, 0.01947808, 
    0.01737224, 0.0162076, 0.01764837, 0.01944655, 0.0222606, 0.02717816, 
    0.03536845, 0.05650507, 0.06321947, 0.04120337, 0.03206087, 0.03554215, 
    0.03804819, 0.07916573, 0.156093, 0.1160528, 0.09258255, 0.1023445, 
    0.09987763, 0.1019111, 0.1124373, 0.1086621, 0.1017343, 0.09681256, 
    0.09373278, 0.1017623, 0.1071018, 0.1143094, 0.1101851, 0.1033055, 
    0.09849041, 0.09678009, 0.09340531, 0.09704743, 0.1008223, 0.1010491, 
    0.09730842, 0.09796206, 0.09943736, 0.09926825, 0.09550188, 0.09170355, 
    0.09014843, 0.08864548, 0.08925509, 0.09028072, 0.08975887, 0.08855143, 
    0.08655528, 0.08483701, 0.08303815, 0.08039567, 0.07954492, 0.07924804, 
    0.0784074, 0.07697187, 0.0754536, 0.07501186, 0.07579702, 0.07425829, 
    0.07095867, 0.0691491, 0.06822985, 0.06829111, 0.06820032, 0.06681692, 
    0.06541313, 0.0646193, 0.0631753, 0.06159781, 0.0608938, 0.05944663, 
    0.05799183, 0.05646692, 0.05471076, 0.05412109, 0.05433499, 0.05475651, 
    0.05540223, 0.05410841, 0.053584, 0.05398789, 0.05437659, 0.05431935, 
    0.05457671, 0.05446195, 0.05421485, 0.0543045, 0.05445789, 0.05501227, 
    0.05693343, 0.05821076, 0.05601759, 0.05310571, 0.05100412, 0.05140315, 
    0.05162438, 0.05100681, 0.04957069, 0.04888743, 0.04689576, 0.04574344, 
    0.04400501, 0.04249143, 0.04206889, 0.04351845, 0.04459305, 0.04525734, 
    0.04513573, 0.04537329, 0.04521352, 0.04484322, 0.04425162, 0.04392715, 
    0.04322641, 0.04244391, 0.03992599, 0.03682606, 0.03405325, 0.03150869, 
    0.02787144, 0.02460959, 0.0218059, 0.01947377, 0.01709642, 0.01798262, 
    0.01237205, 0.008934046, 0.008028573, 0.01081841, 0.0123152, 0.01541103, 
    0.0171841, 0.0158437, 0.01485456, 0.01467359, 0.01622154, 0.02032279, 
    0.02582178, 0.0295556, 0.03594408, 0.04371949, 0.04867326, 0.05328501, 
    0.05705246, 0.05954409, 0.06080029, 0.06247237, 0.06154153, 0.05917801, 
    0.05728995, 0.05657687, 0.05680973, 0.05737357, 0.05935, 0.0603366, 
    0.06161631, 0.06220876, 0.06092765, 0.06022766, 0.05877761, 0.05784182, 
    0.05668852, 0.05558584, 0.05474332, 0.05457274, 0.05514583, 0.05527539, 
    0.05433467, 0.05499487, 0.05546792, 0.05426003, 0.05082246, 0.04689219, 
    0.04461863, 0.04300637, 0.04065809, 0.04169397, 0.04240528, 0.04337975, 
    0.04240301, 0.03933728, 0.03743591, 0.03556706, 0.03468807, 0.03502769, 
    0.03443017, 0.03346115, 0.03339814, 0.0341818, 0.03437179, 0.03426626, 
    0.03347699, 0.03323458, 0.03251954, 0.03213334, 0.03190809, 0.03133494, 
    0.0308997, 0.03081602, 0.03080318, 0.02972643, 0.02841917, 0.02727256, 
    0.02578109, 0.02326784, 0.02122737, 0.01979793, 0.01619091, 0.01329449, 
    0.01241085, 0.01204667, 0.01306948, 0.0149572, 0.011859, 0.009728142, 
    0.007869643, 0.006443527, 0.006064469, 0.006216401,
  0.007702785, 0.007202177, 0.007241657, 0.007240824, 0.006855425, 
    0.006871633, 0.007266527, 0.007905065, 0.009355527, 0.01214083, 
    0.01364843, 0.01299774, 0.01289559, 0.01372928, 0.01440604, 0.01416517, 
    0.01244876, 0.01080748, 0.0100405, 0.01027019, 0.01109705, 0.01224135, 
    0.01270843, 0.01187592, 0.01161346, 0.01241835, 0.01352596, 0.01967999, 
    0.02380824, 0.01760996, 0.01278313, 0.01096481, 0.009203539, 0.009436044, 
    0.01021398, 0.01258801, 0.01606756, 0.01913337, 0.0242442, 0.02914364, 
    0.03355455, 0.01848138, 0.01214631, 0.01214587, 0.01299873, 0.01383652, 
    0.01413138, 0.0117729, 0.01347039, 0.01498307, 0.01480434, 0.01715752, 
    0.01816238, 0.01735566, 0.01607412, 0.01789683, 0.02119102, 0.01663239, 
    0.01904109, 0.03136082, 0.04561248, 0.05954093, 0.06183754, 0.04349394, 
    0.02616005, 0.01579968, 0.01250528, 0.01219133, 0.01283104, 0.01395856, 
    0.01520811, 0.01640825, 0.01777063, 0.02092593, 0.02362951, 0.03041007, 
    0.03217885, 0.02755413, 0.02745416, 0.02948223, 0.03391225, 0.06055184, 
    0.1114153, 0.1242085, 0.09681721, 0.09241401, 0.09007484, 0.09681591, 
    0.1190677, 0.1100515, 0.09253266, 0.08657434, 0.09204021, 0.09822105, 
    0.0956039, 0.09830134, 0.09829932, 0.09707402, 0.09336299, 0.09303288, 
    0.09130894, 0.09419025, 0.09730496, 0.09746855, 0.09871069, 0.09911104, 
    0.09882084, 0.100272, 0.09910451, 0.09512925, 0.09388231, 0.09271462, 
    0.09360343, 0.09506825, 0.0952318, 0.09451299, 0.09199613, 0.0896496, 
    0.08776873, 0.08665646, 0.08717053, 0.08694018, 0.08515701, 0.08331536, 
    0.08166904, 0.08116927, 0.08270828, 0.08348184, 0.0818115, 0.07997812, 
    0.07829089, 0.07646949, 0.07556945, 0.07471247, 0.07363842, 0.07315337, 
    0.07174486, 0.06992877, 0.06860125, 0.06694146, 0.06532927, 0.0642202, 
    0.06279985, 0.06170065, 0.06096869, 0.06128743, 0.06184585, 0.06096357, 
    0.059576, 0.05889075, 0.05937621, 0.0596026, 0.06039957, 0.06153199, 
    0.0621085, 0.06199883, 0.05997753, 0.05908462, 0.06001336, 0.06162939, 
    0.06125964, 0.05806154, 0.05536518, 0.05513403, 0.0561679, 0.05648759, 
    0.05492525, 0.05378427, 0.051285, 0.04976443, 0.04827218, 0.0471526, 
    0.04645033, 0.04751719, 0.04831155, 0.04872405, 0.04804708, 0.04742165, 
    0.04676427, 0.04604665, 0.04535789, 0.04466965, 0.0433539, 0.04257442, 
    0.04060633, 0.03805286, 0.03489672, 0.03194331, 0.02837553, 0.02487509, 
    0.02156414, 0.0193832, 0.01773181, 0.01901403, 0.01305764, 0.01246868, 
    0.008458099, 0.01077873, 0.01397014, 0.01722193, 0.01719726, 0.0157354, 
    0.01384213, 0.01340648, 0.01559222, 0.01939878, 0.02258429, 0.02691547, 
    0.03180879, 0.03927828, 0.04556859, 0.0516292, 0.05759864, 0.06152161, 
    0.06269756, 0.06417903, 0.0653841, 0.06428628, 0.06205937, 0.06088642, 
    0.06113383, 0.06181365, 0.06219049, 0.0621651, 0.06452105, 0.06791762, 
    0.06971915, 0.06972919, 0.06792641, 0.06541996, 0.06424841, 0.06325252, 
    0.06137078, 0.05962456, 0.05905711, 0.05921366, 0.05852098, 0.05784984, 
    0.0578548, 0.05727201, 0.05539107, 0.0537995, 0.0520474, 0.05064392, 
    0.04880779, 0.04857126, 0.04755056, 0.04737921, 0.04679589, 0.04381391, 
    0.04117589, 0.0398793, 0.03883892, 0.03818434, 0.03691622, 0.03553404, 
    0.03490043, 0.03582041, 0.03623437, 0.03616021, 0.0361199, 0.0362346, 
    0.03554299, 0.03417617, 0.03388758, 0.03364896, 0.03355668, 0.03347963, 
    0.0329606, 0.03186177, 0.03057545, 0.02895045, 0.02770053, 0.02588935, 
    0.02284811, 0.02146141, 0.01859891, 0.01628218, 0.01476946, 0.01484872, 
    0.0185331, 0.02229206, 0.02061357, 0.01779174, 0.01220696, 0.009481939, 
    0.008117607, 0.00811334,
  0.01111596, 0.009986917, 0.009116527, 0.009051984, 0.008708533, 
    0.008417395, 0.008923099, 0.009716745, 0.01243591, 0.01506473, 
    0.01656579, 0.01617047, 0.01560694, 0.01565029, 0.01565772, 0.01589199, 
    0.01621505, 0.01688696, 0.01636635, 0.01663998, 0.0165628, 0.01591851, 
    0.01465099, 0.01347483, 0.01236972, 0.01275933, 0.01407964, 0.01911747, 
    0.03169802, 0.02416412, 0.01504253, 0.01246471, 0.01063403, 0.01036631, 
    0.0111493, 0.01467762, 0.01985026, 0.02487534, 0.03330473, 0.0380624, 
    0.03034054, 0.01407087, 0.01353705, 0.01363728, 0.01354002, 0.01396587, 
    0.0124218, 0.01446531, 0.01566331, 0.016807, 0.01743367, 0.02030065, 
    0.02023391, 0.01998223, 0.01528221, 0.01932623, 0.02259622, 0.02129974, 
    0.0275757, 0.0423193, 0.05286578, 0.05233381, 0.03280684, 0.01675237, 
    0.01250789, 0.01230216, 0.01234705, 0.01305125, 0.01483361, 0.01416091, 
    0.01552746, 0.01608333, 0.01950982, 0.02144975, 0.02260116, 0.0251757, 
    0.02650953, 0.02673158, 0.0283056, 0.02829988, 0.03287845, 0.04092025, 
    0.07546392, 0.1126065, 0.09865422, 0.08961054, 0.0908939, 0.09216218, 
    0.09903374, 0.09241159, 0.0806573, 0.08122134, 0.08101371, 0.0814764, 
    0.08316753, 0.08767092, 0.09065105, 0.09169296, 0.08961662, 0.09006844, 
    0.0880419, 0.09127013, 0.09368603, 0.09468377, 0.1067408, 0.1009549, 
    0.0980103, 0.09975378, 0.09882048, 0.09770036, 0.09699258, 0.09791368, 
    0.09868345, 0.100628, 0.1013915, 0.1006537, 0.09865303, 0.09637851, 
    0.09431265, 0.09346336, 0.09445629, 0.0942307, 0.09277916, 0.09102129, 
    0.08887067, 0.08723839, 0.08779725, 0.08947233, 0.08937856, 0.08930377, 
    0.08840916, 0.08623625, 0.08509147, 0.08388659, 0.08275138, 0.0814668, 
    0.07972521, 0.07824124, 0.07721604, 0.07516614, 0.07281904, 0.07143617, 
    0.07059535, 0.06989351, 0.06877694, 0.06796867, 0.06793984, 0.06774347, 
    0.06636217, 0.06472427, 0.06457573, 0.06442475, 0.06424456, 0.06543444, 
    0.06658924, 0.06682502, 0.06482281, 0.06413951, 0.06318856, 0.0636308, 
    0.06491556, 0.06277741, 0.06040328, 0.05960365, 0.060506, 0.06093474, 
    0.05933668, 0.05804759, 0.05511319, 0.05345815, 0.05245303, 0.051663, 
    0.05097593, 0.05205816, 0.05234743, 0.05271281, 0.05158115, 0.05029447, 
    0.04942387, 0.04875187, 0.04777267, 0.046308, 0.04463447, 0.04312471, 
    0.04145503, 0.03877668, 0.03603686, 0.03276804, 0.02941649, 0.02594423, 
    0.02240826, 0.02024314, 0.01876068, 0.01851326, 0.01776348, 0.01142095, 
    0.01055364, 0.01246902, 0.01646909, 0.01925272, 0.01804842, 0.01572601, 
    0.01328557, 0.01446534, 0.01611969, 0.01878511, 0.02197379, 0.02611405, 
    0.03077502, 0.0373926, 0.04343975, 0.04970783, 0.05649955, 0.06173996, 
    0.06337028, 0.0638376, 0.0661332, 0.06734022, 0.06670226, 0.06646419, 
    0.0663607, 0.06607094, 0.06613592, 0.06349724, 0.06455725, 0.07104186, 
    0.07669693, 0.07811049, 0.07676157, 0.07475986, 0.07370916, 0.07213446, 
    0.06957897, 0.06680939, 0.06470434, 0.06367537, 0.06246288, 0.06093329, 
    0.06073003, 0.06017403, 0.05907326, 0.05845834, 0.05687613, 0.05517319, 
    0.05375144, 0.05566449, 0.05395289, 0.05230462, 0.05097532, 0.04722549, 
    0.04453163, 0.04339833, 0.04235368, 0.04110925, 0.04024861, 0.03884504, 
    0.03711714, 0.03697244, 0.03751992, 0.03783867, 0.03835328, 0.03877336, 
    0.03868683, 0.03688674, 0.03615808, 0.03609205, 0.03605814, 0.03558928, 
    0.0347676, 0.03416104, 0.03270534, 0.030948, 0.02976325, 0.02737022, 
    0.02487746, 0.02351483, 0.02137131, 0.01940271, 0.01762813, 0.0181999, 
    0.02092737, 0.0261527, 0.02946194, 0.02900968, 0.01912925, 0.01395531, 
    0.01290811, 0.01181668,
  0.01746594, 0.01538051, 0.01211247, 0.01205783, 0.01321285, 0.01315823, 
    0.01199865, 0.01247683, 0.01474915, 0.016809, 0.01743297, 0.0178513, 
    0.01770493, 0.01711205, 0.0173209, 0.01865074, 0.01951562, 0.02114483, 
    0.02201308, 0.02048652, 0.01778022, 0.01615675, 0.01522499, 0.01434528, 
    0.01302634, 0.01325675, 0.01364628, 0.01758118, 0.03518008, 0.02844577, 
    0.01513071, 0.01368276, 0.01323343, 0.01302908, 0.01411349, 0.01860064, 
    0.02461747, 0.03306279, 0.03822659, 0.03371357, 0.02015364, 0.0169686, 
    0.01754847, 0.01445789, 0.01354593, 0.01403955, 0.01519293, 0.01548033, 
    0.01736778, 0.01725372, 0.01718942, 0.02059472, 0.01828102, 0.01885096, 
    0.0167604, 0.0195177, 0.02881199, 0.03076928, 0.0415757, 0.05107898, 
    0.05691709, 0.03383255, 0.01632625, 0.01202293, 0.01563491, 0.01801452, 
    0.01786623, 0.01677781, 0.01589382, 0.01271996, 0.01239296, 0.01357613, 
    0.01775507, 0.0219226, 0.02123135, 0.02378104, 0.02685745, 0.02689346, 
    0.02764001, 0.02826482, 0.03372522, 0.03808283, 0.05482568, 0.08593382, 
    0.08918605, 0.08228, 0.08940327, 0.09266552, 0.08910593, 0.08354303, 
    0.07770605, 0.07098353, 0.06642859, 0.0672583, 0.07185608, 0.07869349, 
    0.08219524, 0.08225308, 0.08330455, 0.08476745, 0.08515283, 0.09008037, 
    0.09240736, 0.09648879, 0.1010108, 0.09212814, 0.1030885, 0.09961738, 
    0.1002232, 0.1022497, 0.1011291, 0.1002656, 0.1011596, 0.1027733, 
    0.1038984, 0.1045722, 0.1036065, 0.1015884, 0.1003106, 0.1000719, 
    0.1004769, 0.1001561, 0.0982759, 0.09706972, 0.09563832, 0.09411392, 
    0.09345754, 0.09451842, 0.09495272, 0.09502756, 0.09527335, 0.09499998, 
    0.09438775, 0.09296374, 0.09149025, 0.08986254, 0.08758634, 0.08566698, 
    0.08576308, 0.08454651, 0.08170635, 0.07954271, 0.07832479, 0.07739746, 
    0.07647037, 0.07537008, 0.07462896, 0.0747222, 0.07396091, 0.07241262, 
    0.07130452, 0.07008538, 0.06913119, 0.06921601, 0.06949332, 0.06907261, 
    0.06904007, 0.06989937, 0.06842909, 0.06809635, 0.06856763, 0.06780322, 
    0.06498362, 0.06394248, 0.06418331, 0.06457032, 0.06352288, 0.0628282, 
    0.06004624, 0.05839392, 0.05745579, 0.05584345, 0.05496617, 0.05643062, 
    0.05622154, 0.05622053, 0.05554437, 0.05352155, 0.05194654, 0.05131572, 
    0.05022933, 0.04826024, 0.04603292, 0.04389391, 0.04175187, 0.03918521, 
    0.03688796, 0.0336183, 0.03001066, 0.02770049, 0.0251797, 0.02172663, 
    0.01905944, 0.01792645, 0.02051962, 0.01148717, 0.01350394, 0.01573176, 
    0.01986062, 0.02196619, 0.01922195, 0.01653947, 0.01390613, 0.01584462, 
    0.01635148, 0.01881581, 0.02221041, 0.02651523, 0.03041961, 0.03565004, 
    0.04167236, 0.04781783, 0.05462564, 0.06040992, 0.06383572, 0.06556483, 
    0.06719989, 0.07002868, 0.07180583, 0.07210096, 0.07455251, 0.07255716, 
    0.07120787, 0.06767525, 0.06608675, 0.06955972, 0.07818141, 0.08326257, 
    0.08448081, 0.08324505, 0.08228307, 0.08162006, 0.07890512, 0.07552085, 
    0.0722106, 0.06992558, 0.06756778, 0.06624347, 0.06554347, 0.06525733, 
    0.06420222, 0.06327455, 0.06124215, 0.05835992, 0.05618419, 0.0585724, 
    0.0590586, 0.05742267, 0.05543291, 0.05263465, 0.0493577, 0.04695642, 
    0.0462642, 0.04489508, 0.04410337, 0.04299046, 0.04128137, 0.03983794, 
    0.03960465, 0.03983018, 0.04060962, 0.04026766, 0.04039424, 0.03975814, 
    0.03899817, 0.0386235, 0.03873048, 0.0382665, 0.0368122, 0.0361022, 
    0.03534195, 0.03398187, 0.03332516, 0.03183383, 0.02901712, 0.02668456, 
    0.02452204, 0.0225431, 0.02041864, 0.0196026, 0.02141988, 0.0270209, 
    0.03275333, 0.03915533, 0.03045883, 0.02210893, 0.02195533, 0.02015205,
  0.03190061, 0.02861509, 0.02040225, 0.01717739, 0.01729947, 0.01714558, 
    0.01795104, 0.01896921, 0.01884736, 0.01848995, 0.01957365, 0.02054489, 
    0.02037113, 0.01960263, 0.01951013, 0.02072939, 0.02272785, 0.02417885, 
    0.02262759, 0.01883844, 0.01686952, 0.01667002, 0.01642375, 0.01542344, 
    0.01430379, 0.01447945, 0.01436229, 0.01569628, 0.02600362, 0.03012158, 
    0.01744035, 0.01522478, 0.01531739, 0.01595777, 0.01887704, 0.02486075, 
    0.03130488, 0.03511679, 0.02723609, 0.02252588, 0.01933275, 0.01978305, 
    0.01634748, 0.01434919, 0.01356437, 0.0151145, 0.01594515, 0.01716007, 
    0.01938133, 0.02120448, 0.01993105, 0.01868982, 0.01878911, 0.01788838, 
    0.01634578, 0.02095607, 0.03225104, 0.03961439, 0.04805453, 0.055603, 
    0.03761397, 0.01883567, 0.01120892, 0.01345779, 0.01681249, 0.02053034, 
    0.01967555, 0.01821843, 0.01822277, 0.01239731, 0.01278404, 0.01536245, 
    0.01899402, 0.02215226, 0.02251262, 0.02515891, 0.02640126, 0.02713736, 
    0.02535859, 0.02772281, 0.0317228, 0.03956061, 0.05041928, 0.0697338, 
    0.07233902, 0.07744594, 0.07940111, 0.07034053, 0.06957179, 0.07188441, 
    0.06622445, 0.0590132, 0.05639899, 0.05706885, 0.06143714, 0.06771497, 
    0.07048136, 0.07123715, 0.07277457, 0.07638816, 0.08011579, 0.08372024, 
    0.08635587, 0.090965, 0.0973651, 0.09951139, 0.09474859, 0.09880047, 
    0.09939201, 0.1039746, 0.1068945, 0.1006364, 0.1004031, 0.1029777, 
    0.1048542, 0.10552, 0.1047917, 0.1030421, 0.1025841, 0.1023587, 
    0.1027311, 0.1033788, 0.1031714, 0.102528, 0.1015266, 0.1002162, 
    0.0995919, 0.09973503, 0.09961156, 0.1001376, 0.1006148, 0.1010199, 
    0.1013594, 0.1007662, 0.09931656, 0.09828383, 0.09637339, 0.09426758, 
    0.09443168, 0.09401425, 0.09098703, 0.08836053, 0.08696324, 0.08576622, 
    0.0845679, 0.08300712, 0.08174333, 0.08131916, 0.08081357, 0.08059967, 
    0.07936386, 0.07792122, 0.07709207, 0.07563405, 0.07483378, 0.0737128, 
    0.07397866, 0.07600378, 0.07539073, 0.07500592, 0.07470814, 0.07376413, 
    0.07081442, 0.06921431, 0.06870851, 0.06821184, 0.0677986, 0.06797623, 
    0.06659594, 0.06512559, 0.06279764, 0.05825403, 0.05751454, 0.06068995, 
    0.06085333, 0.06001671, 0.05919243, 0.05788381, 0.05601826, 0.05413562, 
    0.05252583, 0.04998043, 0.04751821, 0.0450665, 0.04237961, 0.03988803, 
    0.03735538, 0.03469108, 0.03120513, 0.03028043, 0.02684843, 0.02405054, 
    0.02330963, 0.01984179, 0.01589381, 0.01318038, 0.01598375, 0.02023447, 
    0.02246168, 0.02051709, 0.01751969, 0.01525372, 0.01418551, 0.01655047, 
    0.01654014, 0.01853738, 0.02208541, 0.02635347, 0.02975144, 0.03435825, 
    0.04041836, 0.04748812, 0.05555832, 0.06084787, 0.06521536, 0.06714357, 
    0.06875461, 0.07207622, 0.07687203, 0.07862182, 0.07911944, 0.08429705, 
    0.07981386, 0.07561602, 0.07338119, 0.0724215, 0.07786427, 0.0857144, 
    0.09028246, 0.09016886, 0.09017589, 0.08963481, 0.08787088, 0.08506184, 
    0.08105826, 0.07822187, 0.0752258, 0.07333867, 0.0718476, 0.07145646, 
    0.07005199, 0.06836751, 0.06508251, 0.06071417, 0.05923263, 0.06128274, 
    0.06274089, 0.06209114, 0.05945735, 0.05700788, 0.05435481, 0.05186808, 
    0.05114539, 0.05112612, 0.05031082, 0.04916129, 0.04784143, 0.04550716, 
    0.04422083, 0.04407448, 0.04381982, 0.04274179, 0.04300522, 0.04336794, 
    0.04268906, 0.04207643, 0.04202314, 0.04178028, 0.04016201, 0.03888994, 
    0.03830495, 0.03736042, 0.0364745, 0.03499484, 0.03293252, 0.03036648, 
    0.02805363, 0.02588197, 0.02338213, 0.02134623, 0.02058057, 0.02288681, 
    0.02864956, 0.03609339, 0.03360033, 0.03193428, 0.03595137, 0.0339033,
  0.03528801, 0.04084082, 0.03203811, 0.02674182, 0.02974573, 0.03455781, 
    0.03353352, 0.02857655, 0.02383387, 0.02176163, 0.0224294, 0.02295853, 
    0.02248874, 0.02243132, 0.02334931, 0.02464806, 0.02660646, 0.02631318, 
    0.02383978, 0.02322789, 0.02043633, 0.01939515, 0.01881931, 0.01743416, 
    0.01688098, 0.01750728, 0.01747507, 0.01806017, 0.02543532, 0.02816975, 
    0.02216134, 0.01924454, 0.01923412, 0.02194142, 0.02557302, 0.03139441, 
    0.03876485, 0.03238606, 0.02112527, 0.02162511, 0.02475047, 0.02827056, 
    0.02762039, 0.01956709, 0.01637077, 0.01675448, 0.0182095, 0.01977542, 
    0.02413873, 0.02563146, 0.026098, 0.02484458, 0.02214598, 0.01956011, 
    0.02301839, 0.02467229, 0.03336103, 0.03960921, 0.04754495, 0.034323, 
    0.02701691, 0.01907323, 0.01841358, 0.0142225, 0.0177462, 0.01936362, 
    0.02035329, 0.01710286, 0.01672192, 0.01495298, 0.01638083, 0.01961188, 
    0.02346651, 0.02708328, 0.0285851, 0.02710475, 0.0263004, 0.0254832, 
    0.02488622, 0.02773106, 0.03088713, 0.03823053, 0.0465743, 0.0467936, 
    0.05454955, 0.06562273, 0.07305701, 0.07067204, 0.06829161, 0.06402514, 
    0.05747692, 0.05577671, 0.05185765, 0.04896141, 0.05317352, 0.06003851, 
    0.06007282, 0.06029914, 0.06291817, 0.07041337, 0.07888734, 0.07919123, 
    0.08728545, 0.08392996, 0.09043255, 0.09966941, 0.1052723, 0.1059026, 
    0.1034222, 0.1091632, 0.1399949, 0.1189405, 0.1039307, 0.09996921, 
    0.1036281, 0.1051553, 0.1054647, 0.1052722, 0.1054425, 0.105109, 
    0.1047876, 0.1058753, 0.1072287, 0.1075988, 0.107572, 0.1063929, 
    0.1052366, 0.1051836, 0.105248, 0.1048975, 0.1043968, 0.1044682, 
    0.1046762, 0.1043373, 0.1035286, 0.103546, 0.1021033, 0.1005108, 
    0.1003998, 0.1006252, 0.09882135, 0.09577073, 0.09381008, 0.09272122, 
    0.0909436, 0.08938599, 0.08808373, 0.0868566, 0.08617878, 0.08645174, 
    0.08626927, 0.08583946, 0.08590508, 0.0847249, 0.08339286, 0.08132224, 
    0.08058802, 0.0820637, 0.08289639, 0.08210922, 0.08147711, 0.08087914, 
    0.07828607, 0.07571352, 0.0743585, 0.07368144, 0.07319881, 0.0732208, 
    0.07184593, 0.06965494, 0.06520473, 0.06182472, 0.06342975, 0.06500436, 
    0.06498595, 0.06425335, 0.0632422, 0.06231133, 0.06053412, 0.05760019, 
    0.05511631, 0.05276264, 0.04996751, 0.0466284, 0.04307041, 0.0407166, 
    0.03787699, 0.03510327, 0.03260573, 0.0323272, 0.03018622, 0.03125244, 
    0.02559697, 0.01877759, 0.01286712, 0.01450397, 0.01750398, 0.01983034, 
    0.01797057, 0.01649716, 0.01717466, 0.01635363, 0.01567105, 0.01582987, 
    0.01625075, 0.01807074, 0.02150563, 0.02605774, 0.03096531, 0.03595543, 
    0.04170066, 0.04694962, 0.05402264, 0.06086541, 0.06586319, 0.06791881, 
    0.07012461, 0.0744274, 0.08043888, 0.08309651, 0.08825433, 0.08656718, 
    0.08621321, 0.08396605, 0.08052991, 0.07776875, 0.07811267, 0.0837266, 
    0.08954158, 0.09246077, 0.09410181, 0.09563102, 0.09576352, 0.09337255, 
    0.08980234, 0.08715574, 0.08425066, 0.08142035, 0.07857464, 0.07739921, 
    0.07593726, 0.07184324, 0.06561626, 0.06415686, 0.06602275, 0.06561596, 
    0.06536181, 0.06656635, 0.06604441, 0.06332437, 0.06103538, 0.05810628, 
    0.05645872, 0.05686807, 0.05639332, 0.05504815, 0.05396966, 0.05174006, 
    0.04949917, 0.04884738, 0.04849221, 0.04673491, 0.04679098, 0.04782287, 
    0.04760197, 0.0462175, 0.04477285, 0.04507923, 0.04455355, 0.04346017, 
    0.04248635, 0.04185801, 0.0407882, 0.03895551, 0.03669228, 0.0342778, 
    0.03192878, 0.02951072, 0.02638089, 0.02332512, 0.02165655, 0.02119774, 
    0.02464468, 0.0310335, 0.02871304, 0.03108479, 0.02810752, 0.03089389,
  0.02657738, 0.03090815, 0.0362053, 0.04612613, 0.04806787, 0.04148809, 
    0.03970605, 0.03567774, 0.0269144, 0.025593, 0.02426643, 0.02296703, 
    0.02405585, 0.02669443, 0.02854173, 0.03003098, 0.03091663, 0.03013233, 
    0.02785692, 0.02660879, 0.02310771, 0.02201774, 0.02694539, 0.04010286, 
    0.03514135, 0.04428552, 0.04971707, 0.03679192, 0.03224021, 0.0415859, 
    0.03326391, 0.02451313, 0.02599656, 0.02991056, 0.0343339, 0.04086294, 
    0.03677997, 0.03139848, 0.02726421, 0.04720385, 0.05902017, 0.05705322, 
    0.04089927, 0.03530259, 0.02641551, 0.02062428, 0.02281589, 0.02316922, 
    0.02617401, 0.02481807, 0.02490285, 0.02851625, 0.03128221, 0.0299415, 
    0.03490641, 0.03352585, 0.03062758, 0.02258383, 0.0219853, 0.021051, 
    0.02251294, 0.01934702, 0.0156457, 0.01971498, 0.01701875, 0.01726917, 
    0.01953766, 0.01986992, 0.02089755, 0.01789398, 0.01763549, 0.01853344, 
    0.02284813, 0.02514915, 0.02361653, 0.02007161, 0.0183431, 0.01875429, 
    0.02033256, 0.02538056, 0.02933321, 0.03662539, 0.03651395, 0.03302515, 
    0.03784966, 0.04614569, 0.0496957, 0.05560592, 0.05353939, 0.05074103, 
    0.05055138, 0.05321518, 0.04775044, 0.04402233, 0.04962955, 0.05122773, 
    0.05117424, 0.0538689, 0.05935841, 0.0664425, 0.07378972, 0.07779068, 
    0.07673334, 0.08056045, 0.08245205, 0.08953117, 0.09606395, 0.09968918, 
    0.1054512, 0.1153287, 0.119799, 0.1102449, 0.1080522, 0.09705032, 
    0.09826684, 0.1033007, 0.1060163, 0.1081182, 0.109324, 0.1092331, 
    0.1087651, 0.1091732, 0.1105756, 0.1119588, 0.1129006, 0.1121988, 
    0.1106586, 0.1094983, 0.1090927, 0.1086696, 0.1081259, 0.1074889, 
    0.1066361, 0.1064344, 0.1063704, 0.1055384, 0.1045155, 0.1030226, 
    0.1030303, 0.1036806, 0.1031423, 0.1005915, 0.09847894, 0.0974789, 
    0.09621055, 0.09541325, 0.09443447, 0.09301557, 0.09167912, 0.0916828, 
    0.09150668, 0.09198647, 0.09306788, 0.09281877, 0.09159441, 0.08905793, 
    0.08730913, 0.08794845, 0.08885989, 0.08855269, 0.08818256, 0.08761884, 
    0.08603176, 0.08405764, 0.08197993, 0.08069365, 0.07846809, 0.07590491, 
    0.07212438, 0.07118396, 0.07320445, 0.07334724, 0.07166632, 0.07045334, 
    0.06992024, 0.06841966, 0.06701238, 0.06599136, 0.06423615, 0.06179352, 
    0.05847532, 0.05565923, 0.05233953, 0.04891682, 0.04514544, 0.0419339, 
    0.03857651, 0.03551905, 0.0342752, 0.03443597, 0.03998564, 0.03488401, 
    0.03148773, 0.02043119, 0.01374237, 0.01601001, 0.01739408, 0.01895351, 
    0.01486228, 0.01507694, 0.0188652, 0.01966688, 0.01814363, 0.01653621, 
    0.01667767, 0.01977881, 0.02287751, 0.02726925, 0.0326114, 0.0380611, 
    0.04285042, 0.04825753, 0.0560795, 0.06478675, 0.06901842, 0.07093713, 
    0.07226765, 0.07655127, 0.08106604, 0.08454854, 0.08330059, 0.0867613, 
    0.08840986, 0.0853766, 0.08332749, 0.08141104, 0.07966659, 0.0825066, 
    0.08720079, 0.09139403, 0.09485837, 0.09829929, 0.1006189, 0.1005772, 
    0.0973845, 0.09345997, 0.09018108, 0.08795546, 0.08378163, 0.07970339, 
    0.07599057, 0.07404473, 0.07473668, 0.07490262, 0.07322403, 0.07108711, 
    0.07000932, 0.0699352, 0.0705454, 0.07024855, 0.06868964, 0.06623441, 
    0.06379641, 0.06288283, 0.06206673, 0.06015568, 0.05871642, 0.05725506, 
    0.05577279, 0.05494652, 0.05439211, 0.05251594, 0.05127336, 0.05265076, 
    0.05346876, 0.05268105, 0.05044344, 0.04995129, 0.05060989, 0.04946997, 
    0.04728674, 0.04584975, 0.04499405, 0.04313792, 0.04125714, 0.03901226, 
    0.03639219, 0.03330058, 0.02985153, 0.02702835, 0.02432158, 0.02259763, 
    0.0253789, 0.03142175, 0.0322036, 0.02843173, 0.02227671, 0.02336618,
  0.0217677, 0.02281153, 0.02600558, 0.02949497, 0.03235905, 0.03389651, 
    0.03247138, 0.02898149, 0.0269528, 0.0275199, 0.02638372, 0.03134943, 
    0.03067197, 0.03064165, 0.03192446, 0.03242294, 0.03415293, 0.05198728, 
    0.03930805, 0.03091771, 0.02632649, 0.02762528, 0.04130503, 0.04802873, 
    0.04651294, 0.05269199, 0.03298747, 0.04367891, 0.05289525, 0.05206367, 
    0.04384334, 0.03757684, 0.03664189, 0.03911293, 0.04474816, 0.04243525, 
    0.02685192, 0.02679838, 0.04046333, 0.06751722, 0.05311635, 0.0394306, 
    0.03248311, 0.03015099, 0.03250324, 0.03072042, 0.02535082, 0.02623317, 
    0.02538497, 0.01986568, 0.01885906, 0.022305, 0.02535244, 0.02405533, 
    0.02743978, 0.03387768, 0.03131848, 0.02093022, 0.01133825, 0.01182568, 
    0.01860026, 0.02063757, 0.02041134, 0.01714322, 0.01217306, 0.009611398, 
    0.009696502, 0.01252325, 0.01621763, 0.02015996, 0.02054155, 0.01791563, 
    0.01809904, 0.01794293, 0.01490932, 0.01102711, 0.01348782, 0.01830809, 
    0.02490792, 0.03012181, 0.03297153, 0.03529236, 0.0302604, 0.0261338, 
    0.02639097, 0.03025765, 0.03464751, 0.03977492, 0.0413917, 0.04227654, 
    0.04314953, 0.05021503, 0.04295394, 0.03910645, 0.04265007, 0.04377675, 
    0.04718107, 0.05046318, 0.05367614, 0.06003761, 0.06766, 0.07165402, 
    0.08442254, 0.08411714, 0.0788463, 0.07897808, 0.08246048, 0.08784815, 
    0.0953125, 0.1056883, 0.1068597, 0.1142088, 0.1072008, 0.09653702, 
    0.09345049, 0.09869108, 0.1041358, 0.1077409, 0.1112894, 0.1122409, 
    0.1119529, 0.1122025, 0.11234, 0.1128325, 0.1137019, 0.1138325, 0.11285, 
    0.1121515, 0.1116771, 0.1112567, 0.1111154, 0.1104523, 0.1093683, 
    0.1089031, 0.1089093, 0.1081249, 0.1068007, 0.1053061, 0.104707, 
    0.1047483, 0.1052575, 0.1047146, 0.1028025, 0.1020387, 0.1016351, 
    0.1015656, 0.1014912, 0.100049, 0.09829204, 0.09745868, 0.09672171, 
    0.09705582, 0.09846905, 0.09843653, 0.09776678, 0.09576004, 0.09415313, 
    0.0933122, 0.09359922, 0.09417224, 0.09431983, 0.09374472, 0.0934583, 
    0.09240799, 0.08939816, 0.08500148, 0.07954565, 0.07678316, 0.07925273, 
    0.0825463, 0.08267865, 0.08003312, 0.07774004, 0.07572974, 0.07355057, 
    0.07230906, 0.07189542, 0.07038681, 0.06700826, 0.06471034, 0.06224311, 
    0.0586508, 0.05478476, 0.05119878, 0.04707834, 0.04321396, 0.03991112, 
    0.03732433, 0.03744612, 0.03843624, 0.04250112, 0.03975403, 0.03778687, 
    0.0185605, 0.01391589, 0.0163123, 0.01781816, 0.01844816, 0.01729162, 
    0.01466013, 0.02118368, 0.02410177, 0.02438294, 0.01469257, 0.01797185, 
    0.02103244, 0.02382378, 0.02859209, 0.03463355, 0.03937027, 0.04388626, 
    0.04974231, 0.05708685, 0.06440689, 0.06946143, 0.07237957, 0.0737029, 
    0.0768654, 0.08099788, 0.08449844, 0.08723166, 0.08737041, 0.08784232, 
    0.08883356, 0.08520276, 0.08436541, 0.08245218, 0.08115657, 0.08343475, 
    0.08826824, 0.09421687, 0.09966578, 0.1020104, 0.1024554, 0.1016288, 
    0.0990991, 0.09621935, 0.09231292, 0.08603954, 0.08269184, 0.08503722, 
    0.08748802, 0.08607799, 0.08195944, 0.07973085, 0.07839298, 0.07713819, 
    0.07600043, 0.07556175, 0.07518145, 0.07479636, 0.07368284, 0.07220609, 
    0.07041268, 0.06872135, 0.06662628, 0.06421141, 0.06218112, 0.06080905, 
    0.06184522, 0.06152833, 0.05999162, 0.05796338, 0.05758531, 0.05854512, 
    0.05843553, 0.05662278, 0.05514772, 0.05475205, 0.0544349, 0.05183014, 
    0.05037106, 0.04957863, 0.04777248, 0.04575442, 0.04392082, 0.04128746, 
    0.03809334, 0.03457781, 0.03227899, 0.03043664, 0.03175489, 0.03357984, 
    0.03696828, 0.03891862, 0.03598714, 0.02351075, 0.02244309,
  0.02296671, 0.01956274, 0.02084469, 0.02427148, 0.02637105, 0.02756848, 
    0.0277799, 0.02620885, 0.02632625, 0.0287625, 0.02878714, 0.03310172, 
    0.03590739, 0.03667276, 0.03485438, 0.03590055, 0.03940766, 0.0564314, 
    0.05096595, 0.04200652, 0.0307769, 0.03687795, 0.04882458, 0.04799355, 
    0.04336839, 0.03867025, 0.03459547, 0.03501843, 0.04044332, 0.04315966, 
    0.03999236, 0.04180036, 0.04785277, 0.04599041, 0.03362447, 0.03179336, 
    0.02556898, 0.0336372, 0.05468859, 0.06086767, 0.03454703, 0.02309696, 
    0.01947111, 0.02117213, 0.02721082, 0.02873607, 0.02742006, 0.02455911, 
    0.01911496, 0.0167211, 0.01749767, 0.02063829, 0.02380193, 0.02867288, 
    0.03322182, 0.0427628, 0.03966686, 0.02730205, 0.01332883, 0.011915, 
    0.02121608, 0.02366861, 0.01255746, 0.006696028, 0.005961561, 
    0.006032153, 0.006455214, 0.006930431, 0.008456758, 0.01149745, 
    0.01736573, 0.01919211, 0.01591683, 0.01299045, 0.01005999, 0.01079328, 
    0.01852604, 0.02053137, 0.02568923, 0.02904687, 0.02846318, 0.02300612, 
    0.01921467, 0.01773576, 0.0200005, 0.0222814, 0.02505408, 0.03037374, 
    0.03203749, 0.03474978, 0.03694912, 0.04596516, 0.04122649, 0.03877633, 
    0.03979504, 0.04149336, 0.04290563, 0.04546275, 0.04935263, 0.05648309, 
    0.06373618, 0.07096955, 0.07660516, 0.06867811, 0.06968514, 0.07130475, 
    0.07430509, 0.07666371, 0.07960449, 0.08637345, 0.1002515, 0.104656, 
    0.09456084, 0.08933623, 0.09036735, 0.09266078, 0.09846322, 0.1030715, 
    0.1074585, 0.1110846, 0.1128119, 0.1140091, 0.1140351, 0.1134841, 
    0.1134303, 0.1132805, 0.1125347, 0.1123183, 0.1125, 0.1120718, 0.1120236, 
    0.1122391, 0.1118265, 0.1113226, 0.1109038, 0.1104689, 0.1097034, 
    0.1084148, 0.107213, 0.106474, 0.1071582, 0.1079943, 0.1070367, 
    0.1064322, 0.1058267, 0.1056498, 0.1055129, 0.1046248, 0.1032788, 
    0.1021265, 0.1014189, 0.1017797, 0.1025051, 0.1023634, 0.1021652, 
    0.1015258, 0.1003765, 0.09918484, 0.09910995, 0.09937214, 0.09968002, 
    0.09897543, 0.09806346, 0.09508792, 0.08979344, 0.08749875, 0.08923312, 
    0.09037165, 0.08972759, 0.08826765, 0.08659859, 0.08473796, 0.08289883, 
    0.08055523, 0.07831218, 0.07610168, 0.07463734, 0.07362304, 0.07198932, 
    0.06815536, 0.06503621, 0.06134621, 0.05777181, 0.0539711, 0.04929965, 
    0.04484799, 0.04156431, 0.04180237, 0.04371461, 0.04518721, 0.04320109, 
    0.04686266, 0.03575751, 0.01567353, 0.01460813, 0.01486736, 0.0146058, 
    0.01685501, 0.01684129, 0.01414944, 0.0194489, 0.02578055, 0.02210362, 
    0.01674452, 0.02134035, 0.02344741, 0.02644008, 0.03172937, 0.03686608, 
    0.04086905, 0.04568132, 0.05206994, 0.058298, 0.06358862, 0.06767643, 
    0.06943902, 0.07138054, 0.07504468, 0.07878207, 0.08196237, 0.08509706, 
    0.08915468, 0.09089872, 0.09331498, 0.09088067, 0.08623645, 0.08460069, 
    0.08119702, 0.08333939, 0.08764371, 0.09343947, 0.09827956, 0.09979011, 
    0.1006237, 0.1019671, 0.1010906, 0.09775373, 0.0955321, 0.09694228, 
    0.09855299, 0.09776523, 0.09559894, 0.09365989, 0.09135629, 0.08938093, 
    0.08833193, 0.08708932, 0.08481231, 0.08330178, 0.08192596, 0.08102062, 
    0.08013907, 0.07798894, 0.07630832, 0.07538424, 0.07319099, 0.07085965, 
    0.06945444, 0.06786631, 0.06805201, 0.06789136, 0.06643905, 0.06471027, 
    0.06363641, 0.06415846, 0.06423356, 0.06149882, 0.05936678, 0.05816605, 
    0.05768834, 0.05635783, 0.05580905, 0.05431111, 0.05227226, 0.05110205, 
    0.04911942, 0.04594756, 0.04300874, 0.04053634, 0.03958107, 0.04058256, 
    0.04330438, 0.04347946, 0.04430283, 0.04172881, 0.03766224, 0.03191133, 
    0.02557473,
  0.02749713, 0.02178955, 0.02058662, 0.02281234, 0.0248695, 0.02671688, 
    0.02756687, 0.02850359, 0.02724988, 0.03002688, 0.03253771, 0.03675822, 
    0.04010719, 0.04019118, 0.03850866, 0.04242481, 0.06507979, 0.07097032, 
    0.06294995, 0.05128786, 0.04146392, 0.05268553, 0.06343538, 0.06841326, 
    0.05561257, 0.04468272, 0.0429352, 0.04208143, 0.04143338, 0.04038415, 
    0.04185422, 0.04381797, 0.04405566, 0.03636824, 0.02936303, 0.02985077, 
    0.03827522, 0.05871955, 0.05752824, 0.04661476, 0.02883621, 0.023438, 
    0.02045135, 0.02138097, 0.02362169, 0.02493371, 0.0232124, 0.01966652, 
    0.01741908, 0.01775122, 0.01928959, 0.02173383, 0.02492139, 0.03156098, 
    0.03697169, 0.0483635, 0.03732872, 0.02394859, 0.0167472, 0.01335818, 
    0.01841104, 0.01588448, 0.009278811, 0.008112933, 0.00665712, 
    0.005666666, 0.00525643, 0.005599291, 0.00639461, 0.007234303, 
    0.008334531, 0.009990718, 0.01212123, 0.01244138, 0.01134941, 0.01373991, 
    0.01901979, 0.02128027, 0.01976541, 0.02025691, 0.01583453, 0.0122864, 
    0.01106042, 0.0122956, 0.01508285, 0.01648929, 0.01970649, 0.02406557, 
    0.02537257, 0.02877727, 0.03061797, 0.0430294, 0.04466505, 0.04153652, 
    0.04039136, 0.04141286, 0.04361679, 0.04737808, 0.05219486, 0.05889215, 
    0.06536592, 0.07184027, 0.06936385, 0.06477687, 0.06063507, 0.06278803, 
    0.06718475, 0.06963681, 0.07181439, 0.07520672, 0.08169809, 0.08768384, 
    0.09734681, 0.09500744, 0.08916912, 0.08888935, 0.09195255, 0.0957489, 
    0.1017166, 0.1064467, 0.1089224, 0.1107275, 0.1116325, 0.1123574, 
    0.1126144, 0.1123922, 0.1118895, 0.1110952, 0.1107233, 0.109724, 
    0.1088296, 0.1097311, 0.1104902, 0.1105963, 0.110337, 0.1106471, 
    0.1103447, 0.1094978, 0.1090454, 0.108507, 0.108297, 0.1089361, 
    0.1085866, 0.1082182, 0.1077674, 0.106771, 0.1065738, 0.1064784, 
    0.1060475, 0.1041099, 0.1033636, 0.103666, 0.1038356, 0.1037323, 
    0.1038514, 0.1045978, 0.104654, 0.1046243, 0.103962, 0.1030526, 
    0.1019919, 0.0991545, 0.09706634, 0.09804067, 0.1006714, 0.1016152, 
    0.1001954, 0.09626956, 0.09335323, 0.0919237, 0.09115642, 0.08980945, 
    0.08756875, 0.08551686, 0.08401457, 0.08215726, 0.07992302, 0.07764718, 
    0.0758532, 0.07289734, 0.06946747, 0.06501668, 0.06033824, 0.05587157, 
    0.05135902, 0.0472197, 0.04424644, 0.04790555, 0.05142221, 0.05129855, 
    0.04952889, 0.049732, 0.02850285, 0.01948284, 0.0211359, 0.01507326, 
    0.01460153, 0.01576137, 0.01843936, 0.0157855, 0.01984718, 0.02312983, 
    0.02857143, 0.01882109, 0.02380945, 0.02632719, 0.02994337, 0.03496162, 
    0.0387787, 0.04244135, 0.0475417, 0.05320527, 0.0579684, 0.06213665, 
    0.06593391, 0.0683694, 0.07084293, 0.07313375, 0.07698715, 0.08089609, 
    0.08299191, 0.08530562, 0.08816475, 0.08874742, 0.08920014, 0.08636145, 
    0.08589567, 0.08319785, 0.08329298, 0.08740954, 0.09158085, 0.09377605, 
    0.09412324, 0.09455191, 0.09682965, 0.1009, 0.1044486, 0.1065528, 
    0.1065131, 0.1059197, 0.1049142, 0.1039323, 0.1034996, 0.1024676, 
    0.1006607, 0.098461, 0.09744567, 0.09621016, 0.094674, 0.09264452, 
    0.09088057, 0.0891452, 0.08679855, 0.08331664, 0.080423, 0.07870039, 
    0.077186, 0.07662769, 0.07551687, 0.07465259, 0.07374006, 0.07257737, 
    0.07106401, 0.07038273, 0.07003134, 0.06869818, 0.06658871, 0.06483117, 
    0.06279468, 0.06248945, 0.06181329, 0.06060519, 0.05897596, 0.05758232, 
    0.05672169, 0.05486951, 0.05153075, 0.0488475, 0.04693336, 0.04795728, 
    0.0530996, 0.060973, 0.05464267, 0.05128893, 0.04880899, 0.03897588, 
    0.03435656, 0.02991412,
  0.03676881, 0.02989335, 0.02653757, 0.025911, 0.02561498, 0.02705185, 
    0.02971318, 0.03300631, 0.02911216, 0.03217326, 0.03624387, 0.03700568, 
    0.05385138, 0.04062817, 0.04475374, 0.04784571, 0.08156218, 0.06994871, 
    0.06487147, 0.05515066, 0.05039846, 0.05733498, 0.06511418, 0.07429702, 
    0.0814553, 0.07598065, 0.05940824, 0.05167248, 0.06105803, 0.07827087, 
    0.09091559, 0.1084317, 0.08967068, 0.07175527, 0.04307422, 0.04095761, 
    0.04988444, 0.05264683, 0.0609715, 0.04973309, 0.03171586, 0.0257701, 
    0.02325596, 0.02257261, 0.02355758, 0.02303529, 0.02116834, 0.01955477, 
    0.01938029, 0.02032254, 0.02175582, 0.02269897, 0.02555664, 0.02898133, 
    0.03615971, 0.03551846, 0.03251539, 0.03262365, 0.04357388, 0.03886511, 
    0.0202713, 0.01764661, 0.01735195, 0.01745824, 0.01245958, 0.00805888, 
    0.006489329, 0.00603241, 0.006437859, 0.006862533, 0.007290101, 
    0.007086771, 0.006574982, 0.006416553, 0.007363969, 0.008688821, 
    0.009927988, 0.0105626, 0.01082384, 0.008994242, 0.007238162, 
    0.007589396, 0.009210009, 0.01024091, 0.01118641, 0.01243752, 0.01445899, 
    0.01899363, 0.02329672, 0.02606203, 0.02761289, 0.03160004, 0.03922746, 
    0.04518835, 0.04489448, 0.04522447, 0.04542049, 0.04670229, 0.05532632, 
    0.06567261, 0.06975805, 0.07910325, 0.06929859, 0.06047815, 0.0581899, 
    0.05584553, 0.05965872, 0.06396894, 0.06701565, 0.07085023, 0.07658965, 
    0.08428985, 0.08966635, 0.08193357, 0.08796675, 0.08674007, 0.08764568, 
    0.09084215, 0.09465848, 0.09886713, 0.1030183, 0.1050546, 0.1060065, 
    0.1068866, 0.1075659, 0.1084434, 0.1083621, 0.1074285, 0.1070907, 
    0.1071347, 0.1065404, 0.1061018, 0.1069337, 0.1078203, 0.1085812, 
    0.1089417, 0.10906, 0.1088514, 0.1082154, 0.107225, 0.1069023, 0.1068917, 
    0.1069195, 0.1067166, 0.1066464, 0.1060743, 0.106117, 0.1066268, 
    0.1069343, 0.1058592, 0.1050394, 0.1047955, 0.1051896, 0.1055364, 
    0.1056127, 0.1060909, 0.1061866, 0.105384, 0.1025674, 0.1003092, 
    0.1008697, 0.1047713, 0.1085968, 0.1092802, 0.1081678, 0.1061117, 
    0.1033529, 0.1000028, 0.09775407, 0.0967878, 0.09585041, 0.09453404, 
    0.09340946, 0.0913605, 0.0891905, 0.08658844, 0.08437332, 0.08216918, 
    0.07970591, 0.07604957, 0.07264392, 0.06855479, 0.06392093, 0.05897142, 
    0.05391987, 0.04978645, 0.04759344, 0.05378363, 0.05989235, 0.05705593, 
    0.04683335, 0.04092682, 0.02220173, 0.0222827, 0.02065813, 0.01719823, 
    0.01449668, 0.01797529, 0.02381818, 0.02172594, 0.01600742, 0.02156149, 
    0.02549407, 0.02204619, 0.02474875, 0.02712716, 0.03138766, 0.03721078, 
    0.04110075, 0.04509855, 0.04829605, 0.05177836, 0.05663308, 0.05994722, 
    0.0636429, 0.06591575, 0.06812894, 0.07066821, 0.07459552, 0.07823657, 
    0.07894683, 0.07968945, 0.0839648, 0.0868482, 0.09034866, 0.08630339, 
    0.08615687, 0.08640331, 0.08535213, 0.0857168, 0.08730651, 0.08829312, 
    0.09048482, 0.0957337, 0.1022644, 0.1070962, 0.1090158, 0.1087333, 
    0.1080927, 0.1085062, 0.1095169, 0.1103429, 0.1105942, 0.110473, 
    0.1100939, 0.1086413, 0.1072838, 0.1059651, 0.105267, 0.1047593, 
    0.1031719, 0.1002335, 0.09686188, 0.09251671, 0.08892401, 0.08656643, 
    0.08504752, 0.08388264, 0.082691, 0.08107101, 0.08005713, 0.07911357, 
    0.07802863, 0.07660721, 0.07598121, 0.07433082, 0.07222643, 0.0705833, 
    0.06843976, 0.06794471, 0.06745852, 0.06643075, 0.06555288, 0.06420784, 
    0.0622654, 0.06007234, 0.05688527, 0.05397981, 0.05244721, 0.05506855, 
    0.06361842, 0.07910796, 0.07431775, 0.0651367, 0.0551317, 0.04687332, 
    0.04586085, 0.04186793,
  0.03980635, 0.04192683, 0.03676122, 0.0331765, 0.02790927, 0.02837492, 
    0.02914482, 0.03257228, 0.03224352, 0.03531555, 0.04736388, 0.05497104, 
    0.04706616, 0.04773879, 0.05184959, 0.06193518, 0.07635914, 0.06659808, 
    0.07177365, 0.08150133, 0.06697979, 0.06202786, 0.06612743, 0.07031468, 
    0.0732023, 0.0767046, 0.07767351, 0.08064853, 0.07000139, 0.07105269, 
    0.06839159, 0.08168641, 0.08533558, 0.09955238, 0.08195205, 0.06563796, 
    0.05404667, 0.06367705, 0.07520482, 0.05170875, 0.03750598, 0.02914776, 
    0.02568186, 0.02584347, 0.02600649, 0.02467997, 0.02343823, 0.02204233, 
    0.02209202, 0.02229744, 0.02321179, 0.0243915, 0.02371203, 0.02476435, 
    0.02921635, 0.03044016, 0.03308219, 0.02250081, 0.0251653, 0.02501429, 
    0.01746733, 0.01822, 0.01748156, 0.01813481, 0.01770578, 0.01407811, 
    0.01112356, 0.01062151, 0.0118865, 0.01189385, 0.01053354, 0.008554431, 
    0.006511536, 0.006071694, 0.006448301, 0.007070504, 0.008270686, 
    0.007850236, 0.00644878, 0.006394661, 0.006437217, 0.006598915, 
    0.007217047, 0.008489455, 0.00949561, 0.01183537, 0.01440925, 0.01861951, 
    0.02104703, 0.02223834, 0.02304521, 0.02543556, 0.03189456, 0.03812814, 
    0.03913787, 0.03941058, 0.04251502, 0.04629328, 0.05013971, 0.06041276, 
    0.06498, 0.06082484, 0.05829427, 0.05864189, 0.05802429, 0.05304607, 
    0.05380594, 0.05895615, 0.06250497, 0.06646786, 0.07296803, 0.07923455, 
    0.08329943, 0.08243283, 0.08759481, 0.083182, 0.0822009, 0.08476844, 
    0.08787002, 0.0912949, 0.09556583, 0.09977391, 0.1013853, 0.1020606, 
    0.102144, 0.1029382, 0.1035858, 0.1035888, 0.1033836, 0.1034271, 
    0.1036955, 0.104138, 0.104583, 0.1053731, 0.1068016, 0.1074042, 
    0.1074852, 0.1073796, 0.1069091, 0.1056531, 0.1047248, 0.104733, 
    0.1045769, 0.1047802, 0.105164, 0.1054366, 0.1051235, 0.1054358, 
    0.1058062, 0.1064017, 0.1064767, 0.1063351, 0.1065933, 0.1070534, 
    0.1066473, 0.1050844, 0.1042393, 0.1043356, 0.1053319, 0.1074905, 
    0.1099265, 0.1120893, 0.1121891, 0.1098671, 0.1077931, 0.1067884, 
    0.1062863, 0.1050297, 0.1032477, 0.1013272, 0.09975393, 0.09880994, 
    0.09855486, 0.09669168, 0.09433462, 0.09134743, 0.08879401, 0.0860398, 
    0.08270779, 0.07957058, 0.07648063, 0.07253789, 0.0676111, 0.06213355, 
    0.05651491, 0.05284422, 0.05114412, 0.05880193, 0.06652944, 0.06375775, 
    0.04435749, 0.03194279, 0.02281886, 0.02147972, 0.0227381, 0.02057553, 
    0.01690633, 0.01912517, 0.02360901, 0.02292642, 0.01410481, 0.01783853, 
    0.02010923, 0.02506446, 0.02458705, 0.02846833, 0.03267856, 0.03726629, 
    0.04215924, 0.04620448, 0.04830205, 0.05049121, 0.05462527, 0.05820927, 
    0.06169847, 0.06477798, 0.0666576, 0.06962762, 0.0730509, 0.07642881, 
    0.07755146, 0.07703353, 0.08117572, 0.08523336, 0.0889332, 0.09017964, 
    0.084472, 0.08726984, 0.08780495, 0.08882044, 0.08734442, 0.08759975, 
    0.09139077, 0.09665307, 0.1008517, 0.1035774, 0.1060968, 0.1080852, 
    0.1093422, 0.1109987, 0.1126941, 0.1142152, 0.1152344, 0.1161245, 
    0.1165715, 0.1158094, 0.1148623, 0.1141586, 0.1134312, 0.1134282, 
    0.1127152, 0.1107104, 0.1075862, 0.1032582, 0.09890371, 0.09602717, 
    0.09388005, 0.09244923, 0.09121903, 0.08809631, 0.08608861, 0.08514094, 
    0.08416351, 0.08381944, 0.0821996, 0.07905564, 0.076668, 0.07540873, 
    0.07364596, 0.07290992, 0.07269226, 0.0725266, 0.07186846, 0.07053016, 
    0.06792007, 0.06505378, 0.06154968, 0.0591243, 0.05839814, 0.0626445, 
    0.07406975, 0.09322003, 0.08061729, 0.06293496, 0.0568357, 0.05907122, 
    0.04983938, 0.04144244,
  0.1113938, 0.07888833, 0.05153847, 0.04144896, 0.03374708, 0.03190461, 
    0.03906627, 0.04559081, 0.03485248, 0.04699481, 0.0740794, 0.0560114, 
    0.05040957, 0.05276781, 0.06252328, 0.09250935, 0.08361027, 0.06901169, 
    0.07277527, 0.0688237, 0.06894746, 0.0696459, 0.06450003, 0.06442238, 
    0.06352463, 0.06329618, 0.0630411, 0.06076022, 0.05624234, 0.04637861, 
    0.04415152, 0.04696034, 0.06287347, 0.09908244, 0.09622751, 0.0691539, 
    0.07122816, 0.069669, 0.06128941, 0.05255588, 0.03369566, 0.03155575, 
    0.02897599, 0.02960175, 0.02976377, 0.02848378, 0.02680907, 0.02480649, 
    0.02408673, 0.02434615, 0.02424245, 0.02422626, 0.02367736, 0.023727, 
    0.02602695, 0.02630371, 0.02700568, 0.02372438, 0.03056097, 0.02630498, 
    0.02326215, 0.02225678, 0.02447265, 0.0280453, 0.02836361, 0.01958001, 
    0.01604676, 0.01884779, 0.02391281, 0.01999095, 0.01665582, 0.01396416, 
    0.008956182, 0.007316416, 0.006956147, 0.007279823, 0.006497055, 
    0.006081574, 0.00526497, 0.005311864, 0.005800744, 0.006864217, 
    0.008348125, 0.009839904, 0.01109311, 0.01260482, 0.01347158, 0.01453877, 
    0.01621768, 0.01800142, 0.01979741, 0.02118801, 0.0232443, 0.02783888, 
    0.03095893, 0.03257349, 0.03542052, 0.03975244, 0.04565558, 0.05416246, 
    0.05932275, 0.05939659, 0.0579774, 0.05575637, 0.0588121, 0.05349102, 
    0.05225073, 0.05336807, 0.0578232, 0.06192019, 0.06727097, 0.07438206, 
    0.08031175, 0.08176324, 0.08348095, 0.0745641, 0.07778005, 0.07978243, 
    0.0829718, 0.08569112, 0.08898257, 0.09295448, 0.09620748, 0.09752431, 
    0.0976438, 0.09829683, 0.09893787, 0.09898812, 0.09915394, 0.09899701, 
    0.0996722, 0.1010124, 0.1020689, 0.102947, 0.1038369, 0.1048022, 
    0.1050507, 0.1049664, 0.1047199, 0.1034699, 0.1030494, 0.1037602, 
    0.1041571, 0.1044806, 0.1049273, 0.1052551, 0.1053152, 0.1044694, 
    0.1040067, 0.1045137, 0.1040041, 0.1030957, 0.1033336, 0.1043969, 
    0.1069031, 0.1095121, 0.1120885, 0.1134037, 0.1132279, 0.1120762, 
    0.111202, 0.1109149, 0.1110457, 0.1105917, 0.1100148, 0.1099757, 
    0.1096183, 0.1075976, 0.1056713, 0.1043878, 0.1032495, 0.1021453, 
    0.1013801, 0.1003493, 0.09834313, 0.09576757, 0.09313682, 0.08948186, 
    0.08569184, 0.08299747, 0.08020661, 0.07699752, 0.07248184, 0.06707645, 
    0.06104102, 0.05679461, 0.05625574, 0.06365355, 0.07751187, 0.06966083, 
    0.0505326, 0.02977713, 0.02530443, 0.02396941, 0.02525328, 0.0227161, 
    0.01981826, 0.02164511, 0.02867536, 0.02398432, 0.01683885, 0.01695909, 
    0.01846796, 0.02177922, 0.02523921, 0.0292568, 0.03526812, 0.03905614, 
    0.0421701, 0.04518921, 0.04666009, 0.04905066, 0.05252082, 0.05664868, 
    0.06127214, 0.06471611, 0.0667382, 0.06860118, 0.07550102, 0.07596262, 
    0.07534042, 0.07637553, 0.07881268, 0.0807643, 0.07925414, 0.08306254, 
    0.08290333, 0.09022694, 0.09113404, 0.09040459, 0.08921122, 0.08510704, 
    0.08683837, 0.09060955, 0.0953414, 0.09881087, 0.1017909, 0.1038001, 
    0.1061109, 0.1077409, 0.110012, 0.1130492, 0.1155746, 0.1178129, 
    0.1188465, 0.1191798, 0.1187974, 0.1178535, 0.1172337, 0.1173829, 
    0.1176483, 0.1179288, 0.1160627, 0.1126896, 0.1087147, 0.1044504, 
    0.1017856, 0.1001805, 0.09889393, 0.09592687, 0.093057, 0.09123865, 
    0.0901456, 0.08952039, 0.08737672, 0.08432958, 0.0815082, 0.07994034, 
    0.07862177, 0.07857744, 0.07863008, 0.07852133, 0.07752635, 0.07617863, 
    0.07402974, 0.070539, 0.0665336, 0.06430135, 0.06451603, 0.07008344, 
    0.08309419, 0.1104141, 0.1086644, 0.09376837, 0.08255991, 0.08423597, 
    0.0814134, 0.09889945,
  0.08203508, 0.07981997, 0.06933554, 0.05437207, 0.05224568, 0.05143939, 
    0.04725135, 0.04027321, 0.04472325, 0.05576004, 0.05762516, 0.05182862, 
    0.05343891, 0.0750327, 0.09956983, 0.09712866, 0.07964758, 0.07502092, 
    0.07810076, 0.07674213, 0.07390448, 0.07156234, 0.06976917, 0.06714903, 
    0.06576762, 0.06154414, 0.05715623, 0.05410633, 0.05025563, 0.0476946, 
    0.04743666, 0.06340504, 0.1087907, 0.08989388, 0.07601663, 0.07904874, 
    0.07872798, 0.06271104, 0.05328027, 0.03953799, 0.03625235, 0.03261562, 
    0.03359762, 0.03236548, 0.03188309, 0.0307665, 0.02900045, 0.02747638, 
    0.02650626, 0.02532995, 0.02479669, 0.02408833, 0.02336484, 0.02320287, 
    0.02416156, 0.02663718, 0.02943439, 0.03140495, 0.03181626, 0.02807376, 
    0.02739169, 0.02933983, 0.03053007, 0.02454919, 0.02089719, 0.02036336, 
    0.02869088, 0.03004454, 0.02463693, 0.02113496, 0.017835, 0.01314695, 
    0.008903529, 0.007639794, 0.00852416, 0.0076349, 0.007495303, 0.00678598, 
    0.005782855, 0.006351816, 0.007638157, 0.008945436, 0.009887098, 
    0.01188723, 0.0124467, 0.01309102, 0.01332718, 0.01384896, 0.01483076, 
    0.01601942, 0.01783161, 0.01969601, 0.02157399, 0.02357039, 0.02583369, 
    0.03004084, 0.03112243, 0.03278821, 0.03778578, 0.04692416, 0.05450888, 
    0.05921442, 0.05647421, 0.05295222, 0.05679339, 0.05503825, 0.05625081, 
    0.05885329, 0.0542501, 0.05779077, 0.06254514, 0.06886408, 0.07380701, 
    0.07815281, 0.0779324, 0.07102741, 0.07246443, 0.07691061, 0.08109162, 
    0.08442447, 0.08622684, 0.08792976, 0.09012102, 0.09184523, 0.09220427, 
    0.09200601, 0.09254671, 0.09302992, 0.09350518, 0.09369873, 0.09477195, 
    0.09636179, 0.09752837, 0.09848706, 0.09953237, 0.1003493, 0.1008459, 
    0.1014694, 0.1013712, 0.09991118, 0.09891456, 0.09988584, 0.1005614, 
    0.1007413, 0.1009983, 0.1009685, 0.1017765, 0.1020087, 0.1016559, 
    0.1028004, 0.1038706, 0.1050235, 0.1066774, 0.1082385, 0.1102207, 
    0.1119326, 0.1129212, 0.1125721, 0.1120662, 0.1116389, 0.1111114, 
    0.111454, 0.1120267, 0.111964, 0.1115991, 0.111216, 0.1109102, 0.1099021, 
    0.1079614, 0.1059707, 0.1047059, 0.1034408, 0.1023387, 0.1014668, 
    0.100165, 0.09783071, 0.09517606, 0.09265335, 0.0890551, 0.0860618, 
    0.08290505, 0.07923868, 0.07521202, 0.0703311, 0.06492409, 0.06042488, 
    0.06025349, 0.06685072, 0.07375215, 0.07692689, 0.06575657, 0.04087495, 
    0.0307061, 0.02824939, 0.0310671, 0.03510556, 0.03007027, 0.02248254, 
    0.02724695, 0.03475626, 0.02051955, 0.01752838, 0.02063639, 0.0230564, 
    0.02814518, 0.03240946, 0.03702641, 0.03872503, 0.03999711, 0.04153336, 
    0.04444735, 0.04839744, 0.05153206, 0.05594957, 0.06002944, 0.06361876, 
    0.06539466, 0.06786171, 0.07569428, 0.07387663, 0.07155096, 0.07398594, 
    0.08099714, 0.08202482, 0.07975685, 0.08584388, 0.08895419, 0.09444065, 
    0.09209027, 0.08757037, 0.08780383, 0.08276167, 0.08427017, 0.08806215, 
    0.09206637, 0.09497495, 0.0952379, 0.09743448, 0.09839708, 0.1011583, 
    0.1047503, 0.1080322, 0.1113643, 0.1149943, 0.1180094, 0.1198182, 
    0.1211179, 0.1203714, 0.1195316, 0.1199162, 0.1206238, 0.1213765, 
    0.1211424, 0.1195994, 0.1174067, 0.1131635, 0.1090444, 0.106311, 
    0.1044974, 0.1019021, 0.09900184, 0.09689078, 0.09575268, 0.09491934, 
    0.09253563, 0.08934876, 0.08681878, 0.08475932, 0.08288302, 0.08264996, 
    0.08272306, 0.08218303, 0.08118661, 0.08012918, 0.07852182, 0.07492517, 
    0.07134333, 0.06957733, 0.0701581, 0.0747659, 0.0834653, 0.09213686, 
    0.09356271, 0.08861422, 0.08192863, 0.08079179, 0.08072044, 0.08684546,
  0.08795065, 0.09208293, 0.09806655, 0.07026345, 0.07862904, 0.08253876, 
    0.06601311, 0.07251579, 0.07430736, 0.06591796, 0.05721573, 0.0558426, 
    0.06805255, 0.08508848, 0.08511999, 0.08084236, 0.08110025, 0.08464397, 
    0.08178212, 0.07953969, 0.07859192, 0.07102809, 0.07065172, 0.07029733, 
    0.07113142, 0.06754961, 0.06099632, 0.06055247, 0.05647087, 0.05453732, 
    0.05949755, 0.0673674, 0.06209644, 0.06734067, 0.07567224, 0.07280688, 
    0.05651918, 0.04688289, 0.04322335, 0.0416129, 0.03801093, 0.03711852, 
    0.03635903, 0.03626277, 0.03350636, 0.03184542, 0.02905678, 0.02749526, 
    0.0268073, 0.02605917, 0.0254808, 0.02491174, 0.02529237, 0.02485369, 
    0.02465523, 0.0233507, 0.02327622, 0.02167704, 0.01737957, 0.01641778, 
    0.01879061, 0.02142841, 0.02846151, 0.02703468, 0.02160902, 0.01714604, 
    0.02236717, 0.02308455, 0.02433656, 0.01955136, 0.01204186, 0.01111861, 
    0.01172507, 0.01081744, 0.008402817, 0.007119476, 0.007093906, 
    0.007254045, 0.007982713, 0.008628157, 0.008877598, 0.009819274, 
    0.01100324, 0.0118465, 0.01263201, 0.01293616, 0.01318862, 0.01326298, 
    0.01442946, 0.01575224, 0.01723911, 0.01934472, 0.02055047, 0.02258935, 
    0.02600332, 0.02814743, 0.03011874, 0.03067602, 0.03355931, 0.04052335, 
    0.04714962, 0.05421457, 0.05755349, 0.0548539, 0.0513856, 0.05236789, 
    0.05153873, 0.05712175, 0.05921094, 0.05651834, 0.05941395, 0.06559233, 
    0.0690774, 0.07266577, 0.06643695, 0.06784035, 0.07224528, 0.07502034, 
    0.07864607, 0.08018406, 0.08232899, 0.08377582, 0.08583379, 0.08745486, 
    0.08856113, 0.08870677, 0.08909652, 0.08978675, 0.09082673, 0.09110993, 
    0.09124599, 0.0920784, 0.09309009, 0.09389072, 0.09492306, 0.09508324, 
    0.0954753, 0.09703916, 0.09783181, 0.09655471, 0.09540676, 0.09575228, 
    0.09617808, 0.09680805, 0.0976397, 0.09829593, 0.1002718, 0.1031818, 
    0.1047304, 0.1059695, 0.1069692, 0.107721, 0.1076658, 0.1066791, 
    0.1057373, 0.1062718, 0.1078819, 0.1092137, 0.1097168, 0.1104025, 
    0.1107084, 0.1106478, 0.1106253, 0.110305, 0.1104672, 0.1106539, 
    0.1105815, 0.1097593, 0.1086475, 0.1066922, 0.10436, 0.103367, 0.1028088, 
    0.102157, 0.1006106, 0.09866779, 0.09636673, 0.09422744, 0.09147443, 
    0.08828914, 0.08500541, 0.08115542, 0.07716495, 0.07248463, 0.06726633, 
    0.06312116, 0.0619919, 0.06754469, 0.0756195, 0.08148125, 0.07379005, 
    0.05103153, 0.04596731, 0.04130925, 0.0392205, 0.04642979, 0.03339173, 
    0.02347795, 0.02802544, 0.03623817, 0.02918851, 0.02594258, 0.02982091, 
    0.0303148, 0.03207401, 0.03623542, 0.03714628, 0.0381965, 0.0383779, 
    0.04161479, 0.04655584, 0.04987204, 0.05252838, 0.05566986, 0.05963699, 
    0.06293421, 0.06563152, 0.06787788, 0.07553394, 0.07685371, 0.07477721, 
    0.07894316, 0.08433054, 0.08344151, 0.07910965, 0.08037419, 0.08205006, 
    0.08511437, 0.0903606, 0.08812979, 0.09123938, 0.08532794, 0.08317214, 
    0.08724993, 0.0898622, 0.09417725, 0.09414849, 0.09162101, 0.0918263, 
    0.09336942, 0.09781205, 0.1017009, 0.1054991, 0.1094057, 0.1126261, 
    0.1151692, 0.117552, 0.1193516, 0.1198739, 0.1200058, 0.1205183, 
    0.1211522, 0.1217478, 0.1222766, 0.1208014, 0.1176157, 0.1130994, 
    0.1097517, 0.1078616, 0.1061567, 0.1045507, 0.1025655, 0.1009705, 
    0.09953876, 0.09729187, 0.09477326, 0.09288243, 0.09132263, 0.08964099, 
    0.08748405, 0.08572169, 0.08478656, 0.08464576, 0.08376208, 0.08206869, 
    0.07836872, 0.07588062, 0.07471767, 0.07443093, 0.07559707, 0.07982557, 
    0.08171052, 0.08155385, 0.08115225, 0.07537494, 0.06820328, 0.07096332, 
    0.08240636,
  0.0836534, 0.09530294, 0.0934526, 0.08574619, 0.09113117, 0.1034089, 
    0.08814745, 0.09366011, 0.08937619, 0.09480598, 0.08484399, 0.08389562, 
    0.08137435, 0.07644969, 0.07409547, 0.07373476, 0.0747431, 0.08243819, 
    0.09104055, 0.08784739, 0.08599463, 0.07906435, 0.07301984, 0.06993554, 
    0.07095256, 0.07074603, 0.06890348, 0.07000764, 0.06791507, 0.06570805, 
    0.06435357, 0.06398471, 0.06473574, 0.06423265, 0.06024011, 0.0549722, 
    0.05053634, 0.04570321, 0.04174756, 0.03937872, 0.03932565, 0.03840359, 
    0.03690113, 0.03544934, 0.03403697, 0.03203283, 0.02893537, 0.02625604, 
    0.02581657, 0.02591548, 0.02536604, 0.0249246, 0.02549703, 0.02625402, 
    0.02599252, 0.02498792, 0.02332855, 0.02024321, 0.01754707, 0.01599954, 
    0.01587388, 0.01822518, 0.01990282, 0.03107691, 0.02446504, 0.01746011, 
    0.01599745, 0.01347161, 0.01266537, 0.0105421, 0.009835352, 0.0112329, 
    0.01096103, 0.008974032, 0.009177767, 0.008283495, 0.009642176, 
    0.008566478, 0.009845862, 0.008910028, 0.01013325, 0.01163176, 
    0.01268305, 0.01237119, 0.01265501, 0.01243906, 0.01281247, 0.01368448, 
    0.01502582, 0.01614145, 0.01799677, 0.02103543, 0.02168888, 0.02195384, 
    0.0240737, 0.02756265, 0.03037871, 0.03240871, 0.03344223, 0.03667064, 
    0.04231218, 0.04840798, 0.05148653, 0.05248114, 0.05091854, 0.05231242, 
    0.05280747, 0.05562053, 0.0622035, 0.06134635, 0.05653123, 0.06096757, 
    0.06460927, 0.0648929, 0.06462041, 0.06508361, 0.06726091, 0.07046372, 
    0.07500812, 0.07694405, 0.07909981, 0.08094893, 0.08252729, 0.08331753, 
    0.08424, 0.08506157, 0.08559874, 0.0869565, 0.08869276, 0.08983883, 
    0.09007572, 0.0906284, 0.09087303, 0.0909987, 0.09176509, 0.0924865, 
    0.09354309, 0.09571724, 0.09734133, 0.09761669, 0.09656511, 0.09632891, 
    0.09622724, 0.09606241, 0.09583233, 0.09590926, 0.09695908, 0.09898005, 
    0.1008424, 0.1019976, 0.1028579, 0.1039904, 0.1041102, 0.1031639, 
    0.1021378, 0.1021657, 0.1030812, 0.1042112, 0.1054703, 0.1065833, 
    0.1073314, 0.1080005, 0.1077235, 0.1077152, 0.1084221, 0.1095871, 
    0.1098947, 0.1084984, 0.10732, 0.1062692, 0.1041241, 0.1026979, 
    0.1022683, 0.1018077, 0.1001726, 0.0984263, 0.09676734, 0.09546114, 
    0.09382346, 0.09063433, 0.08683199, 0.08299775, 0.0785089, 0.07369282, 
    0.06923235, 0.06541322, 0.06441262, 0.06775326, 0.07626739, 0.08423916, 
    0.07567319, 0.05646095, 0.05175578, 0.05454523, 0.05470567, 0.04849311, 
    0.03676293, 0.0275214, 0.02593771, 0.03142186, 0.02967362, 0.03142142, 
    0.03331763, 0.03009979, 0.03325854, 0.03508033, 0.03707042, 0.0366667, 
    0.03865153, 0.04092667, 0.04557849, 0.04783443, 0.05161687, 0.05491988, 
    0.05824963, 0.06194049, 0.06473703, 0.06535821, 0.0701751, 0.07465575, 
    0.07389634, 0.07724178, 0.0820177, 0.08132084, 0.08028448, 0.07958621, 
    0.07740492, 0.07916953, 0.08295283, 0.08556765, 0.09134579, 0.09155411, 
    0.08534195, 0.08847443, 0.09111417, 0.09232404, 0.09257879, 0.09234126, 
    0.09120692, 0.08883829, 0.09120295, 0.09528822, 0.09903351, 0.1035637, 
    0.1061831, 0.1080476, 0.1103535, 0.1129224, 0.1153843, 0.1170491, 
    0.1179399, 0.1188983, 0.1202328, 0.1211142, 0.1199419, 0.1183309, 
    0.1158595, 0.113108, 0.1111616, 0.1093515, 0.1080095, 0.1069921, 
    0.1057556, 0.1043836, 0.102426, 0.1005044, 0.09810955, 0.09614659, 
    0.09446901, 0.09182288, 0.08908592, 0.08826549, 0.0888048, 0.08832753, 
    0.08619823, 0.08293314, 0.08071315, 0.07868747, 0.07806434, 0.07803043, 
    0.07676192, 0.07447819, 0.07105763, 0.06611165, 0.06067383, 0.05843334, 
    0.06186777, 0.07140863,
  0.07956576, 0.08416602, 0.0882827, 0.09430947, 0.1039367, 0.1120481, 
    0.1059431, 0.1095602, 0.1043373, 0.1079389, 0.1118615, 0.09992161, 
    0.0895742, 0.07956823, 0.07120088, 0.06552562, 0.06905123, 0.08109983, 
    0.08831586, 0.08675568, 0.08756387, 0.08681095, 0.07981342, 0.07392094, 
    0.06991788, 0.07003245, 0.07073946, 0.07091509, 0.07314925, 0.07141332, 
    0.06799076, 0.06801461, 0.06767426, 0.06323384, 0.06062774, 0.05711771, 
    0.05009837, 0.04499736, 0.04042508, 0.03755337, 0.03718097, 0.03639949, 
    0.03546751, 0.03534164, 0.0345397, 0.03281597, 0.03115089, 0.02911656, 
    0.02731578, 0.02682578, 0.02649575, 0.02673811, 0.02696898, 0.02795179, 
    0.02734555, 0.02692722, 0.02572533, 0.02299423, 0.01995394, 0.01719848, 
    0.01613525, 0.0167288, 0.01964126, 0.02129047, 0.0209737, 0.01973352, 
    0.01823112, 0.0152745, 0.01110283, 0.01369917, 0.01397468, 0.01232192, 
    0.01597398, 0.01329608, 0.01188746, 0.01105342, 0.01099002, 0.01224808, 
    0.01145986, 0.01278017, 0.01691935, 0.01964542, 0.01914808, 0.01754821, 
    0.01604816, 0.01476819, 0.01485513, 0.01623264, 0.01703916, 0.01888276, 
    0.01927505, 0.0207895, 0.02238098, 0.02351598, 0.02545453, 0.02896361, 
    0.03056481, 0.0328295, 0.03403686, 0.03538151, 0.0391328, 0.04389248, 
    0.04879963, 0.0493459, 0.04781689, 0.04913647, 0.05267814, 0.05502459, 
    0.05918983, 0.06490222, 0.06140669, 0.0595035, 0.06228098, 0.06183514, 
    0.05973227, 0.05954874, 0.06304144, 0.06788462, 0.07212118, 0.07533807, 
    0.07768026, 0.07891912, 0.07985467, 0.0807291, 0.08142675, 0.08169914, 
    0.08218694, 0.08359607, 0.0853347, 0.08670183, 0.0868957, 0.08720338, 
    0.0872879, 0.08683348, 0.086904, 0.08783825, 0.08932609, 0.0913026, 
    0.09317356, 0.09485528, 0.09523735, 0.09450933, 0.09387973, 0.09367166, 
    0.09303964, 0.09323278, 0.0938666, 0.09483214, 0.09627496, 0.09732207, 
    0.0984726, 0.09994151, 0.1005373, 0.1005233, 0.1004204, 0.1002534, 
    0.1000699, 0.1005144, 0.101553, 0.102562, 0.103403, 0.1039071, 0.1044796, 
    0.1050289, 0.1057302, 0.1066737, 0.107276, 0.1059775, 0.104942, 
    0.1044113, 0.1036943, 0.1027009, 0.1022215, 0.10152, 0.09986471, 
    0.09788346, 0.09611629, 0.09480361, 0.09348477, 0.09137226, 0.08823581, 
    0.0842211, 0.07949167, 0.0741429, 0.06991828, 0.06738359, 0.06697613, 
    0.07214412, 0.07862259, 0.08779927, 0.08774934, 0.05967775, 0.04725728, 
    0.05392772, 0.05939113, 0.0607378, 0.04816378, 0.03705602, 0.02817934, 
    0.0319215, 0.02934742, 0.02867447, 0.02757704, 0.02863569, 0.03164398, 
    0.0353149, 0.03709419, 0.03777565, 0.03990352, 0.0412863, 0.04368605, 
    0.04661031, 0.05061439, 0.05337076, 0.05741694, 0.05974965, 0.06364542, 
    0.06631637, 0.06800058, 0.07168106, 0.07356742, 0.07315435, 0.07502442, 
    0.07696154, 0.07871649, 0.07934242, 0.07786869, 0.07979745, 0.08337273, 
    0.08226074, 0.08389702, 0.08515415, 0.08611625, 0.08547276, 0.08877301, 
    0.08855983, 0.08701237, 0.08777889, 0.08895386, 0.09781843, 0.09403546, 
    0.09699877, 0.1003049, 0.1020584, 0.1030318, 0.1032197, 0.1036393, 
    0.1062106, 0.1089696, 0.111559, 0.1128869, 0.1138972, 0.11528, 0.1174928, 
    0.1187022, 0.1182979, 0.1163821, 0.1144258, 0.1130718, 0.1115177, 
    0.1099999, 0.1090504, 0.1083105, 0.1075147, 0.1055392, 0.1032608, 
    0.1009389, 0.09920616, 0.0982871, 0.09613355, 0.09381114, 0.09228531, 
    0.09160692, 0.09045088, 0.0878524, 0.08509625, 0.08316203, 0.08143352, 
    0.08046541, 0.07997811, 0.07864826, 0.07660237, 0.07396121, 0.07082865, 
    0.06775986, 0.06566423, 0.06786529, 0.07450761,
  0.07773039, 0.08250708, 0.08846572, 0.09381397, 0.0990283, 0.1039395, 
    0.1018861, 0.09896985, 0.1008654, 0.09839638, 0.1059513, 0.0935018, 
    0.08871276, 0.08165985, 0.07702721, 0.07498597, 0.07846891, 0.08589322, 
    0.09133589, 0.1067113, 0.09610169, 0.08846229, 0.0822915, 0.07727818, 
    0.07505445, 0.07524998, 0.07493724, 0.07409957, 0.07431447, 0.07551374, 
    0.07282234, 0.07187934, 0.06982805, 0.06564271, 0.06158535, 0.05654718, 
    0.05068082, 0.04654969, 0.04366539, 0.04136703, 0.03929803, 0.03764416, 
    0.03702551, 0.03688979, 0.03668079, 0.03560932, 0.03378259, 0.03259836, 
    0.03126186, 0.03058766, 0.02967456, 0.02886626, 0.02963221, 0.0300164, 
    0.02920854, 0.02973564, 0.02906121, 0.02765042, 0.02493257, 0.02150635, 
    0.01940644, 0.01842638, 0.01876793, 0.01971938, 0.02151549, 0.02155285, 
    0.02144581, 0.02224883, 0.0188347, 0.01627218, 0.01585229, 0.02156045, 
    0.02136685, 0.01431998, 0.01493608, 0.01392695, 0.01370869, 0.01711266, 
    0.01866297, 0.01540023, 0.01710432, 0.02119548, 0.02337581, 0.0235769, 
    0.02125283, 0.02057472, 0.01936716, 0.02000055, 0.02177296, 0.02288855, 
    0.02268706, 0.02241054, 0.022093, 0.02286001, 0.02469999, 0.02936804, 
    0.032168, 0.03255225, 0.03412312, 0.03540128, 0.03825853, 0.04313336, 
    0.04816316, 0.05007456, 0.04787459, 0.04770735, 0.05035776, 0.05421518, 
    0.05790623, 0.06436933, 0.06216514, 0.05894053, 0.06008754, 0.05882261, 
    0.05771858, 0.05821593, 0.06082264, 0.06390613, 0.06909426, 0.07272841, 
    0.07474151, 0.07689735, 0.07704273, 0.07765642, 0.07811013, 0.07788581, 
    0.07814968, 0.0794346, 0.08110917, 0.08248366, 0.08274847, 0.08329977, 
    0.08379386, 0.08390906, 0.08405425, 0.08470631, 0.08604401, 0.08767178, 
    0.08925588, 0.09118927, 0.09220286, 0.09216201, 0.09142429, 0.09106515, 
    0.0911162, 0.09183746, 0.09294164, 0.09309351, 0.09357663, 0.09381538, 
    0.09451437, 0.09609004, 0.0967718, 0.09697961, 0.09785015, 0.09840902, 
    0.09789833, 0.09768775, 0.09817939, 0.09908181, 0.09979522, 0.1003116, 
    0.1007225, 0.101849, 0.102792, 0.1033964, 0.1040477, 0.103814, 0.1026493, 
    0.102138, 0.1020466, 0.1018912, 0.1018677, 0.1015358, 0.1002462, 
    0.09811249, 0.09567152, 0.09334793, 0.09178296, 0.09025251, 0.08791397, 
    0.08446258, 0.07964559, 0.07532261, 0.07206099, 0.07060581, 0.07195304, 
    0.07654235, 0.08432275, 0.09039155, 0.07902924, 0.06873474, 0.04786246, 
    0.0518447, 0.05681357, 0.05841524, 0.04526979, 0.04030317, 0.02594484, 
    0.02852773, 0.02819238, 0.0265943, 0.02645935, 0.02771357, 0.03096403, 
    0.03514556, 0.03798101, 0.03859752, 0.04037683, 0.0420718, 0.04360061, 
    0.04687559, 0.05031793, 0.05471509, 0.05712192, 0.05989852, 0.06259795, 
    0.06672839, 0.06841933, 0.0700286, 0.06855842, 0.07220707, 0.07198091, 
    0.07229776, 0.07328048, 0.07563929, 0.0773733, 0.07673525, 0.07728294, 
    0.07721576, 0.08311382, 0.08228885, 0.07732833, 0.08214426, 0.07978525, 
    0.08123248, 0.08005168, 0.08414761, 0.08775009, 0.09472755, 0.1005572, 
    0.1092631, 0.1038394, 0.1026604, 0.09945495, 0.09777825, 0.09750132, 
    0.1014149, 0.104465, 0.1072044, 0.1089746, 0.1101106, 0.1113778, 
    0.1130618, 0.1148472, 0.1162169, 0.1162438, 0.1146254, 0.1129794, 
    0.1114443, 0.1102283, 0.1094715, 0.1087804, 0.1078341, 0.1051398, 
    0.1026585, 0.1008208, 0.1002301, 0.1004115, 0.09858324, 0.09583354, 
    0.09386187, 0.09271508, 0.09141333, 0.08917981, 0.08661851, 0.084383, 
    0.08302479, 0.08159315, 0.08048516, 0.07912823, 0.078082, 0.07645064, 
    0.07512125, 0.07456992, 0.07455049, 0.07551815, 0.07718746,
  0.08279104, 0.0827708, 0.08541322, 0.0898177, 0.09103057, 0.09703558, 
    0.0998041, 0.09953862, 0.09473066, 0.09044228, 0.08847453, 0.08339782, 
    0.08404388, 0.0859189, 0.09085036, 0.1013835, 0.09940422, 0.09741567, 
    0.109743, 0.109042, 0.09201077, 0.08878416, 0.08670046, 0.08297957, 
    0.08192629, 0.08122938, 0.08076217, 0.07925566, 0.0785304, 0.07720555, 
    0.07673887, 0.07504096, 0.07129884, 0.06681405, 0.06226704, 0.05760811, 
    0.05331828, 0.04951533, 0.04736886, 0.04546051, 0.04419125, 0.04336453, 
    0.04291315, 0.04214014, 0.04125732, 0.04013761, 0.03807566, 0.0361847, 
    0.03487764, 0.03348831, 0.03233196, 0.03192225, 0.0321704, 0.03182669, 
    0.03159179, 0.03188534, 0.03183995, 0.03130579, 0.03006002, 0.02818513, 
    0.02497746, 0.02359149, 0.02358039, 0.02422811, 0.0249327, 0.02664839, 
    0.02904348, 0.02954751, 0.02652088, 0.02474844, 0.02421691, 0.02057762, 
    0.0143723, 0.01547143, 0.01654263, 0.0144728, 0.01649381, 0.02002125, 
    0.01955784, 0.01863267, 0.02055993, 0.02330121, 0.02469031, 0.02590717, 
    0.02579638, 0.0293294, 0.03201633, 0.02716902, 0.02479831, 0.02501856, 
    0.02496215, 0.02341697, 0.02213846, 0.02212259, 0.02376675, 0.02724721, 
    0.03216464, 0.03372673, 0.03558541, 0.03673033, 0.03843792, 0.04318349, 
    0.04758338, 0.04938129, 0.04984643, 0.05003056, 0.05105985, 0.05379857, 
    0.05560798, 0.05882848, 0.061741, 0.05990146, 0.05680833, 0.05645812, 
    0.05486664, 0.0553172, 0.05967863, 0.0619775, 0.06562141, 0.06866065, 
    0.07171974, 0.07386877, 0.07481068, 0.0751917, 0.07507838, 0.07423552, 
    0.07384622, 0.07501689, 0.07677566, 0.07800777, 0.07821792, 0.07893779, 
    0.0801002, 0.08099776, 0.0816133, 0.08213249, 0.08307681, 0.08432361, 
    0.08511645, 0.08674444, 0.08860075, 0.08989648, 0.09015702, 0.09009381, 
    0.09010904, 0.09007515, 0.09059882, 0.09087789, 0.09067128, 0.09046076, 
    0.09105229, 0.09219986, 0.09295957, 0.09335902, 0.09394235, 0.09488922, 
    0.0947246, 0.09464674, 0.0945639, 0.09576382, 0.09682447, 0.09716712, 
    0.09737337, 0.09816187, 0.09896514, 0.09968754, 0.1006215, 0.1014742, 
    0.1012713, 0.1006188, 0.1001899, 0.1001817, 0.1000474, 0.09967123, 
    0.09871735, 0.09722359, 0.09524845, 0.09289736, 0.09114534, 0.0895137, 
    0.08722353, 0.08394095, 0.08043893, 0.07722271, 0.07615551, 0.07737809, 
    0.08126063, 0.08093094, 0.08962888, 0.08588777, 0.09785559, 0.07518127, 
    0.04992361, 0.05148366, 0.05520536, 0.04885897, 0.04502919, 0.03770464, 
    0.02615627, 0.02716949, 0.0263667, 0.02611998, 0.02637101, 0.02847158, 
    0.03139084, 0.03439067, 0.03707843, 0.03774152, 0.03912809, 0.04129327, 
    0.04275445, 0.04684407, 0.05006068, 0.05210913, 0.05414318, 0.05625366, 
    0.05844954, 0.06138267, 0.06303, 0.0632324, 0.06585236, 0.06759853, 
    0.06815721, 0.06799487, 0.06823681, 0.07117786, 0.07297023, 0.07300407, 
    0.07357186, 0.07199869, 0.07004656, 0.07640338, 0.0734838, 0.07244906, 
    0.07591734, 0.07591338, 0.07433434, 0.07582252, 0.08204586, 0.09196153, 
    0.09651882, 0.1062033, 0.101007, 0.09725288, 0.0938376, 0.09037922, 
    0.09394915, 0.09801278, 0.1010373, 0.1038155, 0.1062279, 0.1081395, 
    0.1095959, 0.1107128, 0.1126588, 0.1149192, 0.1161677, 0.1143395, 
    0.1122962, 0.1110301, 0.1101933, 0.1098434, 0.1085312, 0.106741, 
    0.1046964, 0.1024752, 0.1006541, 0.1000818, 0.100285, 0.09968206, 
    0.09798677, 0.09604944, 0.09454495, 0.09313699, 0.09114047, 0.08856925, 
    0.08582152, 0.08491726, 0.08402296, 0.08322917, 0.08209364, 0.08068908, 
    0.08031187, 0.08113018, 0.08488786, 0.08842906, 0.08410623, 0.08442354,
  0.0825615, 0.08647542, 0.08661712, 0.09292375, 0.09609766, 0.09201676, 
    0.0897673, 0.09046526, 0.0887439, 0.08787113, 0.08452336, 0.08406488, 
    0.08711067, 0.09313229, 0.09975896, 0.1107354, 0.1092261, 0.1016882, 
    0.09768563, 0.09542567, 0.09280265, 0.09100835, 0.08728459, 0.08577964, 
    0.08498496, 0.08341807, 0.08287838, 0.08282559, 0.08233652, 0.08066811, 
    0.07827923, 0.07566307, 0.07293585, 0.0691542, 0.0644481, 0.05939083, 
    0.05508978, 0.05231126, 0.05099057, 0.04916839, 0.04763458, 0.04665228, 
    0.04690959, 0.0466418, 0.04604937, 0.0442643, 0.04216685, 0.03986724, 
    0.03781935, 0.03546172, 0.03419005, 0.03459968, 0.03478011, 0.03533145, 
    0.03389498, 0.03422685, 0.03490575, 0.03405686, 0.03363874, 0.03234848, 
    0.03045252, 0.02836607, 0.02887781, 0.02969307, 0.03072839, 0.03364788, 
    0.03379336, 0.03355848, 0.03439165, 0.0298358, 0.0204789, 0.01283624, 
    0.01525011, 0.02018784, 0.02177698, 0.01840293, 0.02255202, 0.02198382, 
    0.02125258, 0.01762383, 0.02074361, 0.02249892, 0.02407272, 0.02631101, 
    0.02896678, 0.03243527, 0.03665916, 0.03665178, 0.03193266, 0.02805346, 
    0.0256875, 0.02560595, 0.02428468, 0.02327723, 0.02445145, 0.02646742, 
    0.02938303, 0.03231729, 0.0360738, 0.0368316, 0.0385427, 0.04189776, 
    0.04443424, 0.04625592, 0.05002405, 0.05210344, 0.0540616, 0.05405713, 
    0.05497995, 0.05329214, 0.05559493, 0.05350998, 0.05219407, 0.05625799, 
    0.05543301, 0.05191116, 0.05809152, 0.06162642, 0.06443327, 0.06710296, 
    0.06950442, 0.07149809, 0.07298552, 0.07392337, 0.07317954, 0.07175663, 
    0.07134265, 0.07152468, 0.07271288, 0.0740752, 0.07435737, 0.07429765, 
    0.0750974, 0.07640396, 0.07761776, 0.07900502, 0.07987318, 0.08066025, 
    0.08101958, 0.08291526, 0.08501932, 0.08663786, 0.08747577, 0.08782744, 
    0.08786571, 0.08749545, 0.08732904, 0.08831794, 0.08870824, 0.08814413, 
    0.08851388, 0.08943699, 0.09004473, 0.09036825, 0.09081995, 0.09144148, 
    0.0915219, 0.09161544, 0.09206149, 0.0924651, 0.09305472, 0.09353211, 
    0.09399003, 0.09481209, 0.09569297, 0.0965967, 0.09766289, 0.09860826, 
    0.09954362, 0.0995309, 0.09951448, 0.09873047, 0.09775268, 0.09706987, 
    0.09632714, 0.09521933, 0.09365479, 0.09209839, 0.09029883, 0.08866776, 
    0.08637146, 0.08393372, 0.08185398, 0.08021308, 0.08194272, 0.08505184, 
    0.0969816, 0.09722412, 0.09840426, 0.09480525, 0.09262381, 0.05596667, 
    0.04821047, 0.05078996, 0.05003156, 0.03804777, 0.03252531, 0.02685174, 
    0.02707161, 0.02649026, 0.02744654, 0.0275878, 0.03000888, 0.0322241, 
    0.03304904, 0.03431233, 0.03323276, 0.03440172, 0.03690018, 0.03847948, 
    0.04002029, 0.0442463, 0.04727901, 0.05046192, 0.05217596, 0.05324153, 
    0.05432452, 0.05490819, 0.0570704, 0.05883259, 0.06167458, 0.06284351, 
    0.06402159, 0.06491906, 0.06532989, 0.06787398, 0.06955591, 0.07022852, 
    0.07087255, 0.07083615, 0.0703038, 0.06932766, 0.06913816, 0.06655961, 
    0.06733505, 0.06981979, 0.07251057, 0.07392848, 0.07885714, 0.08659385, 
    0.09101755, 0.09675016, 0.09586521, 0.08936568, 0.09013391, 0.0905432, 
    0.09170796, 0.09474926, 0.09845456, 0.1019718, 0.1050385, 0.1075229, 
    0.1087406, 0.1097497, 0.1113882, 0.113266, 0.114636, 0.1131041, 
    0.1110022, 0.1097174, 0.1090783, 0.109055, 0.1081118, 0.1062842, 
    0.1043066, 0.1028734, 0.1013773, 0.1005494, 0.1004631, 0.1002271, 
    0.09947237, 0.09775557, 0.09615997, 0.09434042, 0.09267703, 0.09113538, 
    0.08943126, 0.0882098, 0.08813772, 0.08713528, 0.08491917, 0.08319531, 
    0.08354782, 0.08603445, 0.08701681, 0.08524786, 0.0847353, 0.08480402,
  0.08371221, 0.08765515, 0.08766367, 0.09269185, 0.09678902, 0.0956047, 
    0.0939877, 0.09259091, 0.09160864, 0.08949471, 0.0889547, 0.08888227, 
    0.09445633, 0.09826382, 0.09840356, 0.09923952, 0.09899521, 0.09615152, 
    0.09647682, 0.09505282, 0.09093148, 0.08896228, 0.08751131, 0.08709747, 
    0.08698458, 0.08667892, 0.08688139, 0.08606668, 0.08511139, 0.08328182, 
    0.07921707, 0.07568995, 0.07287775, 0.06996787, 0.06582896, 0.06106165, 
    0.05648215, 0.05375091, 0.05237762, 0.05077768, 0.04923915, 0.04866253, 
    0.04899842, 0.04921096, 0.04907738, 0.04735169, 0.0456343, 0.04247573, 
    0.03971544, 0.03721115, 0.03595552, 0.03657685, 0.03715095, 0.03734719, 
    0.03649922, 0.03701448, 0.03645588, 0.03548119, 0.03473331, 0.03326451, 
    0.03216297, 0.03068136, 0.03016597, 0.03002136, 0.03179502, 0.03476833, 
    0.04179179, 0.04185332, 0.04029842, 0.03384523, 0.02940972, 0.02464129, 
    0.01893891, 0.02424719, 0.02220408, 0.02128715, 0.02560567, 0.0279502, 
    0.0244574, 0.01988834, 0.02040185, 0.02385001, 0.02732943, 0.03130346, 
    0.03116989, 0.03122068, 0.03496142, 0.03823594, 0.03804348, 0.03349881, 
    0.02865771, 0.02568891, 0.02556696, 0.02546041, 0.02596839, 0.02609785, 
    0.02930922, 0.03154041, 0.03339048, 0.03507857, 0.03706039, 0.03850154, 
    0.04152488, 0.04542317, 0.04876127, 0.04875882, 0.05333345, 0.05547771, 
    0.05707611, 0.04838258, 0.04920714, 0.05507503, 0.0502746, 0.05223343, 
    0.05693176, 0.05248876, 0.05706982, 0.05960551, 0.06286014, 0.06524371, 
    0.06654849, 0.06856455, 0.07110085, 0.07296287, 0.0737403, 0.07142176, 
    0.0693204, 0.06925429, 0.06897873, 0.06927699, 0.06999851, 0.0699072, 
    0.07041988, 0.07155466, 0.07326197, 0.07508221, 0.0764485, 0.07738224, 
    0.07769756, 0.07941426, 0.08137031, 0.08300009, 0.08429206, 0.08514743, 
    0.0853492, 0.08544254, 0.08546238, 0.08609622, 0.08668617, 0.08654514, 
    0.08637431, 0.08687975, 0.08746195, 0.08756953, 0.08817953, 0.08883464, 
    0.08929221, 0.08967832, 0.08984363, 0.09000394, 0.0904319, 0.09093938, 
    0.09183695, 0.09280757, 0.09360544, 0.09396177, 0.09447719, 0.09541012, 
    0.09608819, 0.09644261, 0.09667461, 0.09629122, 0.09498995, 0.09349366, 
    0.09318307, 0.09257083, 0.09186024, 0.09106684, 0.08976904, 0.08801883, 
    0.08542484, 0.08403085, 0.08284189, 0.08263192, 0.08942081, 0.09891972, 
    0.108688, 0.1001177, 0.0931968, 0.08211855, 0.05158988, 0.04743491, 
    0.05042857, 0.05174709, 0.04334046, 0.03163747, 0.02909792, 0.02879947, 
    0.02733606, 0.02506753, 0.02690505, 0.02908636, 0.03134696, 0.03269255, 
    0.03324141, 0.03294627, 0.03264625, 0.03409983, 0.03532813, 0.03751139, 
    0.03905915, 0.04250368, 0.0452918, 0.04849194, 0.05031521, 0.05192375, 
    0.0521, 0.05202628, 0.05353397, 0.05457732, 0.05623339, 0.05713446, 
    0.05793629, 0.0600587, 0.06375109, 0.06603649, 0.06822418, 0.06918143, 
    0.06952715, 0.0708444, 0.06893747, 0.0677058, 0.06414966, 0.06509022, 
    0.06602614, 0.06812756, 0.072108, 0.07297475, 0.07557698, 0.08138416, 
    0.08656927, 0.08954749, 0.09543096, 0.08618597, 0.08588056, 0.08619898, 
    0.08785684, 0.09173444, 0.09570087, 0.09989282, 0.1037606, 0.1063903, 
    0.1077785, 0.1086077, 0.1094788, 0.1105331, 0.1110853, 0.1101138, 
    0.1084585, 0.1071889, 0.1063212, 0.1058719, 0.1055155, 0.1042811, 
    0.1027944, 0.1017549, 0.100997, 0.09998761, 0.09920827, 0.09885447, 
    0.0986516, 0.09786046, 0.09652874, 0.09483761, 0.09287547, 0.09238208, 
    0.09176423, 0.09106898, 0.09204943, 0.09113197, 0.08755592, 0.0844412, 
    0.0852695, 0.08818348, 0.09566173, 0.09005162, 0.08693987, 0.08403363,
  0.08574859, 0.08482164, 0.08638621, 0.09017257, 0.09311842, 0.09551628, 
    0.0943242, 0.09301448, 0.08911811, 0.08567094, 0.08722814, 0.08892899, 
    0.08966501, 0.0907836, 0.09342041, 0.09528777, 0.09361967, 0.09153229, 
    0.09077474, 0.08981614, 0.08932032, 0.08856487, 0.08811302, 0.08868165, 
    0.08918448, 0.08990002, 0.08914412, 0.08701933, 0.0848555, 0.08340723, 
    0.07962517, 0.07653724, 0.07364222, 0.07049206, 0.0668163, 0.06326031, 
    0.05916246, 0.05620232, 0.05352537, 0.0520157, 0.05144667, 0.05125301, 
    0.05138303, 0.05104852, 0.05154894, 0.05041355, 0.04778197, 0.04368981, 
    0.04165451, 0.03931359, 0.03843472, 0.03876848, 0.04013171, 0.03993829, 
    0.03923372, 0.03854844, 0.03754022, 0.03625621, 0.03509345, 0.03351689, 
    0.03260899, 0.03081757, 0.02955417, 0.02916129, 0.03122026, 0.03544559, 
    0.04121903, 0.04541872, 0.04613568, 0.04960314, 0.04616094, 0.03689239, 
    0.03154972, 0.02963307, 0.02807239, 0.02528298, 0.02831359, 0.03387219, 
    0.03136987, 0.02820509, 0.0254843, 0.032648, 0.03850187, 0.0388272, 
    0.03326992, 0.03101244, 0.03111477, 0.03228156, 0.03199897, 0.03028864, 
    0.02812829, 0.02513984, 0.02501844, 0.02636627, 0.02760999, 0.02813557, 
    0.0290967, 0.03172307, 0.03386761, 0.03513787, 0.03593405, 0.03724905, 
    0.03973722, 0.04203745, 0.04749487, 0.04937752, 0.05236911, 0.05060516, 
    0.053167, 0.04934867, 0.04997921, 0.04810456, 0.04643663, 0.04781494, 
    0.04939002, 0.05126603, 0.05505419, 0.05742025, 0.0597071, 0.06219774, 
    0.06382959, 0.06632724, 0.06856788, 0.07259259, 0.07210412, 0.07422783, 
    0.0695732, 0.06507336, 0.06610834, 0.06556954, 0.06630965, 0.06684429, 
    0.06743963, 0.06865901, 0.06978212, 0.07104681, 0.07278711, 0.07410732, 
    0.07430661, 0.07568805, 0.07741555, 0.07923619, 0.0809944, 0.08170491, 
    0.08228137, 0.08284554, 0.08337416, 0.08396251, 0.08372831, 0.08435337, 
    0.08472841, 0.0851911, 0.08579512, 0.08602547, 0.08644567, 0.08661252, 
    0.0869827, 0.08792157, 0.08865527, 0.08898579, 0.08903756, 0.0892107, 
    0.08988267, 0.09045271, 0.09069611, 0.09072268, 0.0909689, 0.09145845, 
    0.09187967, 0.09219348, 0.0924357, 0.09200827, 0.09128509, 0.09089706, 
    0.09076186, 0.09069788, 0.0904491, 0.08926196, 0.08796315, 0.08648956, 
    0.08585246, 0.08462922, 0.08348929, 0.08792669, 0.09487607, 0.105464, 
    0.1155846, 0.09081049, 0.05731233, 0.04130711, 0.04186738, 0.05086747, 
    0.05333212, 0.04915331, 0.04665057, 0.02862379, 0.02936206, 0.02940006, 
    0.02684147, 0.02580055, 0.02701294, 0.02902285, 0.03093762, 0.03202439, 
    0.03222129, 0.03276709, 0.03380711, 0.03526674, 0.03676694, 0.03852249, 
    0.0402512, 0.04297546, 0.04601233, 0.04827234, 0.05012013, 0.05123797, 
    0.0512388, 0.05116378, 0.05156881, 0.05243335, 0.05335642, 0.05398007, 
    0.05418961, 0.05681115, 0.0605892, 0.06408688, 0.06630125, 0.0674411, 
    0.06749709, 0.0674331, 0.06621892, 0.06400026, 0.06120453, 0.06006876, 
    0.06231416, 0.06277756, 0.06532156, 0.06632192, 0.06842475, 0.07250951, 
    0.07811408, 0.07868353, 0.0800239, 0.07941609, 0.0796359, 0.08240834, 
    0.0851803, 0.08853132, 0.09243807, 0.09663661, 0.1008535, 0.1039388, 
    0.1055817, 0.1062119, 0.1064223, 0.1063182, 0.1063285, 0.106066, 0.1053, 
    0.1046128, 0.1035665, 0.1026396, 0.1023759, 0.1022217, 0.1015225, 
    0.100567, 0.09897294, 0.09755172, 0.09693841, 0.09649425, 0.09612861, 
    0.09581725, 0.09528933, 0.09400834, 0.09236579, 0.0921405, 0.09240095, 
    0.0924983, 0.09500292, 0.09571651, 0.09874006, 0.08944634, 0.08760949, 
    0.0905669, 0.1010586, 0.09578606, 0.09208249, 0.08953271,
  0.08658437, 0.0845841, 0.0851331, 0.08778448, 0.09135638, 0.09100523, 
    0.09152486, 0.09017173, 0.08793707, 0.08690297, 0.08465729, 0.08514574, 
    0.08670107, 0.08727293, 0.08609547, 0.08688774, 0.08709402, 0.08816636, 
    0.0889649, 0.08937928, 0.09006149, 0.08961896, 0.08996411, 0.09116072, 
    0.0915722, 0.09111604, 0.0896443, 0.08636374, 0.08281654, 0.07978303, 
    0.07754751, 0.07608151, 0.07353812, 0.07129269, 0.06857555, 0.06546474, 
    0.06287327, 0.06068309, 0.05684181, 0.05502362, 0.05484287, 0.05541428, 
    0.05574714, 0.05534121, 0.05479738, 0.05346734, 0.05056237, 0.04498052, 
    0.04280094, 0.04100163, 0.03921679, 0.03953671, 0.04148877, 0.04177826, 
    0.04181297, 0.04031746, 0.0385203, 0.03728462, 0.03623187, 0.03473642, 
    0.03274352, 0.03092074, 0.0303575, 0.0307982, 0.03234031, 0.03533427, 
    0.03865622, 0.0424513, 0.04638522, 0.04756563, 0.05068956, 0.04835494, 
    0.0383593, 0.03976739, 0.03989594, 0.03449852, 0.03301514, 0.03257196, 
    0.03855477, 0.03789435, 0.03290721, 0.03899308, 0.03666626, 0.0316028, 
    0.02907732, 0.03067148, 0.03143579, 0.03296208, 0.02991068, 0.02501266, 
    0.024991, 0.02408517, 0.02375263, 0.02379674, 0.0262081, 0.02726037, 
    0.0290221, 0.03076881, 0.03374274, 0.03539247, 0.03565591, 0.03639744, 
    0.03842786, 0.04105742, 0.04501266, 0.04766152, 0.05550314, 0.05249427, 
    0.04882639, 0.04893988, 0.0491244, 0.04789237, 0.04683675, 0.04701572, 
    0.04735125, 0.05003987, 0.05333115, 0.05479817, 0.05657042, 0.05868172, 
    0.06124511, 0.06303997, 0.06552113, 0.06992996, 0.0708665, 0.07293587, 
    0.0713136, 0.06377026, 0.06353858, 0.06391053, 0.06386858, 0.06514257, 
    0.0660331, 0.06675749, 0.0672554, 0.0681845, 0.07035859, 0.07161196, 
    0.0732537, 0.07352863, 0.07455348, 0.07610931, 0.07736869, 0.07852015, 
    0.07990509, 0.081081, 0.08197073, 0.08261458, 0.08450457, 0.08439711, 
    0.08408897, 0.08498257, 0.085766, 0.08482853, 0.08477817, 0.08447054, 
    0.08464295, 0.0851474, 0.08643642, 0.08714917, 0.08704732, 0.0873149, 
    0.08766068, 0.08765911, 0.08733951, 0.08692919, 0.08663203, 0.0867197, 
    0.0872838, 0.08811961, 0.08881975, 0.08945148, 0.08948112, 0.08944359, 
    0.08979914, 0.09023596, 0.08970096, 0.08819678, 0.08649889, 0.0860006, 
    0.08567909, 0.08546437, 0.08986323, 0.09343326, 0.1041746, 0.116755, 
    0.09998441, 0.06234347, 0.03949808, 0.04571535, 0.05220936, 0.05390413, 
    0.04962413, 0.04002719, 0.03032448, 0.03155426, 0.03334222, 0.02970444, 
    0.02728639, 0.02738189, 0.02870605, 0.03034722, 0.03166812, 0.03208919, 
    0.0333638, 0.03563824, 0.03734211, 0.03745789, 0.03820922, 0.04061973, 
    0.0421413, 0.04463935, 0.04687842, 0.04874026, 0.05003183, 0.05048791, 
    0.05068677, 0.05087452, 0.05129424, 0.05110363, 0.05192621, 0.05133866, 
    0.05200231, 0.05557698, 0.05936135, 0.06160971, 0.06381829, 0.06515026, 
    0.06574858, 0.06412484, 0.06196699, 0.05883066, 0.05785464, 0.05575331, 
    0.05544157, 0.05581312, 0.0580553, 0.05981291, 0.06192568, 0.06477924, 
    0.06925, 0.07289525, 0.07267942, 0.07303804, 0.07569582, 0.08047771, 
    0.08394434, 0.08772793, 0.09077834, 0.09370327, 0.09761854, 0.1006766, 
    0.1022217, 0.1023719, 0.1023309, 0.10237, 0.1021647, 0.1018277, 
    0.1018995, 0.1016039, 0.1007908, 0.0998919, 0.1003217, 0.10072, 0.100364, 
    0.09933887, 0.09747538, 0.09541938, 0.09443125, 0.09385764, 0.09363377, 
    0.093689, 0.09310623, 0.09229987, 0.0918007, 0.09206451, 0.09216872, 
    0.09210048, 0.09467915, 0.09680217, 0.1030915, 0.09725954, 0.09496678, 
    0.09062847, 0.1027553, 0.1046727, 0.09733707, 0.09196622,
  0.08662438, 0.08343823, 0.08277301, 0.08498958, 0.08770195, 0.08928575, 
    0.09029072, 0.09131797, 0.08925495, 0.08586945, 0.08431756, 0.08401299, 
    0.08647425, 0.08682254, 0.0853757, 0.08503576, 0.08748471, 0.08983606, 
    0.09057964, 0.09173528, 0.09248194, 0.09285863, 0.09242254, 0.09216361, 
    0.09073991, 0.08857426, 0.08696063, 0.08419993, 0.08020745, 0.07651472, 
    0.07425208, 0.07285025, 0.07178843, 0.07136875, 0.06959227, 0.0670794, 
    0.06488683, 0.06196287, 0.05938381, 0.05813063, 0.05838972, 0.05851262, 
    0.05878642, 0.05895633, 0.05840579, 0.05854724, 0.05447232, 0.04861504, 
    0.04427291, 0.04311278, 0.04140373, 0.04137011, 0.0428102, 0.04390264, 
    0.04386538, 0.04235412, 0.04035922, 0.03873773, 0.0370139, 0.03496737, 
    0.03327037, 0.0325953, 0.03284874, 0.03309368, 0.03366138, 0.03414444, 
    0.03517087, 0.03776192, 0.03993244, 0.0426931, 0.04624103, 0.04241036, 
    0.03648819, 0.04191853, 0.0419004, 0.04440048, 0.04491297, 0.03938638, 
    0.03484725, 0.03714945, 0.0376248, 0.0355592, 0.03162374, 0.02993226, 
    0.03009767, 0.0312596, 0.03372844, 0.0355095, 0.03592252, 0.02953893, 
    0.0239402, 0.02521576, 0.02575178, 0.02581447, 0.02565346, 0.02583655, 
    0.02717551, 0.02824247, 0.03021769, 0.03281609, 0.03452361, 0.03604438, 
    0.03744692, 0.04154294, 0.04593484, 0.04507679, 0.04739655, 0.05089669, 
    0.0509946, 0.04933872, 0.0461339, 0.04617912, 0.04568578, 0.04610439, 
    0.04748464, 0.05004674, 0.0528593, 0.05342085, 0.05460681, 0.0563399, 
    0.05824962, 0.0590762, 0.06061428, 0.06527878, 0.06724422, 0.07165834, 
    0.07786047, 0.06515726, 0.06302362, 0.06315927, 0.06354152, 0.06396186, 
    0.0647397, 0.06564789, 0.06599158, 0.06726161, 0.06921557, 0.07050215, 
    0.07139058, 0.07242247, 0.07346106, 0.07455719, 0.0757289, 0.07661734, 
    0.07812262, 0.07935838, 0.08064783, 0.08213413, 0.08311081, 0.0833281, 
    0.08358254, 0.08363952, 0.08497162, 0.08548918, 0.08678573, 0.08111534, 
    0.08174646, 0.082119, 0.08348674, 0.08372728, 0.0834289, 0.08329812, 
    0.08408628, 0.0849376, 0.08462753, 0.08351608, 0.08260053, 0.08249619, 
    0.0827364, 0.08458444, 0.08627845, 0.08662223, 0.0868384, 0.08751638, 
    0.08791707, 0.0879437, 0.08773497, 0.08661957, 0.08481517, 0.08513124, 
    0.08592419, 0.0911928, 0.09597255, 0.1023034, 0.1197709, 0.1086157, 
    0.07942878, 0.04851148, 0.04714495, 0.04924654, 0.05218881, 0.05289641, 
    0.04288738, 0.03010858, 0.03244909, 0.03390051, 0.03173919, 0.0284477, 
    0.02836854, 0.02903652, 0.03173833, 0.0342038, 0.03566636, 0.03580467, 
    0.03595412, 0.03727, 0.03806254, 0.03749017, 0.03879635, 0.04102296, 
    0.04254114, 0.04425936, 0.04604827, 0.04748964, 0.04825762, 0.04839439, 
    0.04839981, 0.04867338, 0.04884669, 0.0490561, 0.04911863, 0.04887104, 
    0.05032561, 0.0546027, 0.05636566, 0.05912283, 0.06127276, 0.06120891, 
    0.06139252, 0.05946634, 0.05813127, 0.05622949, 0.055043, 0.05320476, 
    0.05299846, 0.05363898, 0.05600682, 0.05742682, 0.05898965, 0.0609734, 
    0.06351596, 0.0683551, 0.06957193, 0.07158285, 0.07532343, 0.07860246, 
    0.08276211, 0.08725417, 0.09039044, 0.09252543, 0.09458595, 0.09655324, 
    0.09845379, 0.09979672, 0.09989968, 0.09963857, 0.09915207, 0.09883245, 
    0.09906304, 0.099044, 0.09865096, 0.09803733, 0.0981564, 0.09861125, 
    0.0987471, 0.09792368, 0.09628595, 0.09450492, 0.09305102, 0.0919755, 
    0.09143603, 0.09173883, 0.09124752, 0.09074865, 0.09026342, 0.09044539, 
    0.09051178, 0.09046446, 0.09243742, 0.09690422, 0.1029836, 0.1007763, 
    0.09565762, 0.09178119, 0.09431864, 0.1002519, 0.1013019, 0.09101944,
  0.08410016, 0.08295407, 0.08237162, 0.08413441, 0.0872309, 0.08863794, 
    0.08857597, 0.08800972, 0.08594897, 0.08340227, 0.08253375, 0.08097869, 
    0.08178681, 0.083607, 0.0839863, 0.08437248, 0.08460423, 0.08819577, 
    0.090552, 0.09234463, 0.09219375, 0.09274001, 0.09206109, 0.09108962, 
    0.08898896, 0.08640527, 0.08505262, 0.08287642, 0.07962602, 0.07547119, 
    0.0727073, 0.0714142, 0.07055758, 0.07054801, 0.0700592, 0.06802075, 
    0.06468944, 0.06205563, 0.06000298, 0.05934471, 0.05954609, 0.05966184, 
    0.0599283, 0.06112998, 0.06189848, 0.06260913, 0.05966092, 0.05313564, 
    0.04836529, 0.04568243, 0.04409023, 0.04345505, 0.04443132, 0.04527716, 
    0.04504267, 0.0435337, 0.0415234, 0.03904052, 0.03683173, 0.03518684, 
    0.03465906, 0.0348737, 0.03512063, 0.03547861, 0.03489015, 0.03523616, 
    0.03672665, 0.03831074, 0.03941001, 0.0423148, 0.04676298, 0.04301568, 
    0.03976218, 0.04119166, 0.04498712, 0.04812575, 0.05040729, 0.04427282, 
    0.03824761, 0.03733476, 0.03649988, 0.03227826, 0.0312046, 0.0329106, 
    0.03409342, 0.03271453, 0.03463733, 0.03636846, 0.03867826, 0.03646149, 
    0.02967406, 0.02577897, 0.0265795, 0.02717517, 0.02768504, 0.02778483, 
    0.02916922, 0.03026497, 0.03198135, 0.03296226, 0.03572641, 0.03766595, 
    0.03879857, 0.04124759, 0.04684668, 0.04596091, 0.04646728, 0.04776599, 
    0.04944733, 0.05035359, 0.04873496, 0.0481248, 0.04724671, 0.04673331, 
    0.04740944, 0.04905741, 0.05043606, 0.05107578, 0.05203986, 0.05321522, 
    0.05419946, 0.05444834, 0.0558589, 0.06135982, 0.06022697, 0.06115196, 
    0.06281947, 0.05961887, 0.05911465, 0.06433207, 0.06363026, 0.06371879, 
    0.06315833, 0.06316819, 0.06446795, 0.06564888, 0.06728016, 0.06855917, 
    0.06944329, 0.07060242, 0.07163766, 0.07236886, 0.07345609, 0.07446269, 
    0.07617188, 0.0775779, 0.07848869, 0.07928366, 0.08045989, 0.08108748, 
    0.08096953, 0.08088417, 0.08076733, 0.08055616, 0.0833599, 0.08176793, 
    0.08254059, 0.0806083, 0.08093926, 0.0809895, 0.08166812, 0.08145612, 
    0.0817662, 0.08177903, 0.08218979, 0.0812213, 0.08014445, 0.07964106, 
    0.07982022, 0.0807753, 0.08242497, 0.08315041, 0.08292544, 0.08265502, 
    0.08292814, 0.08314227, 0.08252834, 0.08137669, 0.08273339, 0.08496134, 
    0.08690001, 0.09636553, 0.1021765, 0.11198, 0.1131752, 0.09309145, 
    0.06437001, 0.0518647, 0.04580335, 0.04423377, 0.04321066, 0.04150645, 
    0.03613592, 0.03156669, 0.03458839, 0.03307555, 0.03011916, 0.0294605, 
    0.03146394, 0.03353296, 0.03463323, 0.03758813, 0.03874676, 0.03910189, 
    0.03906491, 0.03917845, 0.03918083, 0.03892726, 0.04019623, 0.04104379, 
    0.04264201, 0.04403429, 0.04500513, 0.04557222, 0.04553023, 0.0452496, 
    0.04490763, 0.04492834, 0.04541081, 0.04633719, 0.04723536, 0.0472804, 
    0.04940872, 0.05243575, 0.05436902, 0.05724909, 0.05861733, 0.058272, 
    0.05688809, 0.05581301, 0.05525374, 0.0542977, 0.05299218, 0.05268736, 
    0.05212404, 0.05194235, 0.05288997, 0.05398608, 0.05482557, 0.05955424, 
    0.06297143, 0.06410087, 0.06651867, 0.07066809, 0.07445951, 0.0783749, 
    0.08276381, 0.08647607, 0.08926824, 0.09122449, 0.09269878, 0.09438657, 
    0.0956856, 0.0964955, 0.09713743, 0.09745255, 0.09648959, 0.09607539, 
    0.0966462, 0.09766664, 0.09754072, 0.0966855, 0.09639155, 0.09680325, 
    0.09663551, 0.09581188, 0.09453332, 0.09313224, 0.09208436, 0.09111498, 
    0.09047984, 0.09047958, 0.09052514, 0.08987416, 0.08904206, 0.08918301, 
    0.08913483, 0.08904751, 0.09042051, 0.09370717, 0.09659341, 0.1009836, 
    0.1016136, 0.1000824, 0.1003438, 0.1039966, 0.106334, 0.08713835,
  0.0827219, 0.08342516, 0.0849273, 0.08594088, 0.08751254, 0.08824693, 
    0.08777242, 0.08795476, 0.08477435, 0.08353663, 0.08461045, 0.08308384, 
    0.08147169, 0.08042289, 0.08216004, 0.08366886, 0.08493175, 0.08935438, 
    0.09054951, 0.0910546, 0.09115615, 0.0903058, 0.08947975, 0.08911202, 
    0.08806015, 0.08646505, 0.08411662, 0.08138409, 0.07861912, 0.07619315, 
    0.07333349, 0.07165474, 0.07061815, 0.06992933, 0.06910644, 0.06759213, 
    0.06483514, 0.06250987, 0.06034542, 0.0596172, 0.05934322, 0.05870036, 
    0.05893403, 0.06107933, 0.06359285, 0.06288293, 0.05997605, 0.05397203, 
    0.05072191, 0.04718325, 0.04563594, 0.04519639, 0.04561509, 0.04532461, 
    0.04531532, 0.04414027, 0.04245427, 0.04077144, 0.03903506, 0.0378213, 
    0.0376568, 0.03786132, 0.03800416, 0.0380311, 0.03732741, 0.03751243, 
    0.03817501, 0.03944135, 0.04121719, 0.04271039, 0.04311774, 0.04236211, 
    0.04068229, 0.04126712, 0.04014562, 0.03957, 0.03959654, 0.04056543, 
    0.03986882, 0.03727537, 0.03317287, 0.03270824, 0.03391391, 0.03775878, 
    0.03807898, 0.03666104, 0.0382354, 0.0383577, 0.03842808, 0.03521816, 
    0.03433055, 0.02970782, 0.02953069, 0.02816545, 0.02938815, 0.03092972, 
    0.03100872, 0.03057728, 0.03161157, 0.03412005, 0.03689267, 0.0378688, 
    0.04116683, 0.042776, 0.04571445, 0.04273506, 0.04446857, 0.04637781, 
    0.04602264, 0.04685693, 0.04486243, 0.046845, 0.04645658, 0.04437067, 
    0.04431996, 0.04499008, 0.04554302, 0.04656665, 0.04812382, 0.04959401, 
    0.05041298, 0.05087869, 0.05331235, 0.05589598, 0.05576911, 0.06275755, 
    0.04816484, 0.05291298, 0.06074607, 0.06404895, 0.06257653, 0.06391029, 
    0.06285334, 0.06243581, 0.06366982, 0.06480759, 0.06602777, 0.06692022, 
    0.06769947, 0.06854475, 0.06948601, 0.07064454, 0.07168838, 0.07276645, 
    0.07418382, 0.07563151, 0.07655057, 0.07693003, 0.07758424, 0.07779239, 
    0.07758192, 0.0775305, 0.07810146, 0.07871127, 0.07909764, 0.07895625, 
    0.08027373, 0.08125998, 0.08712453, 0.08675877, 0.09394397, 0.07827247, 
    0.08075412, 0.08277705, 0.08195405, 0.0805882, 0.07856246, 0.07734416, 
    0.07703792, 0.07727797, 0.07785045, 0.07838608, 0.07801315, 0.07752475, 
    0.07794473, 0.07830957, 0.07825109, 0.08009744, 0.08240737, 0.08647269, 
    0.0957994, 0.1080786, 0.1137527, 0.1142052, 0.1015232, 0.07692423, 
    0.0609814, 0.05071968, 0.04068785, 0.03762452, 0.03425196, 0.03234772, 
    0.02989362, 0.03019405, 0.03054239, 0.03152278, 0.03166796, 0.03401707, 
    0.03579441, 0.03805863, 0.0389029, 0.0390026, 0.03943271, 0.03956197, 
    0.03979852, 0.04046922, 0.04125524, 0.04157991, 0.04251546, 0.04332254, 
    0.04384402, 0.04424089, 0.04442221, 0.04413065, 0.04360219, 0.04336851, 
    0.04340376, 0.04376206, 0.04439146, 0.0456065, 0.04733428, 0.04783321, 
    0.04838997, 0.0495717, 0.05096381, 0.05313159, 0.05433352, 0.05468351, 
    0.05315956, 0.05187672, 0.05083904, 0.05057558, 0.0497628, 0.05062745, 
    0.05068517, 0.05121133, 0.05111219, 0.05326071, 0.05635635, 0.05778505, 
    0.0592852, 0.06175084, 0.06607778, 0.07089826, 0.0755264, 0.0794717, 
    0.08276523, 0.08509122, 0.0871273, 0.08843392, 0.08929934, 0.09033656, 
    0.09132348, 0.0922003, 0.09317959, 0.09331763, 0.09316938, 0.0933079, 
    0.0942397, 0.09546939, 0.09606266, 0.09561586, 0.09562059, 0.09567343, 
    0.09538199, 0.09392607, 0.09265647, 0.09166509, 0.09114792, 0.090875, 
    0.09020635, 0.09013133, 0.08983114, 0.08893208, 0.08825342, 0.08880839, 
    0.08844797, 0.08805986, 0.08868054, 0.09047224, 0.09155463, 0.0966737, 
    0.1001392, 0.1069659, 0.1135684, 0.1057824, 0.09493527, 0.08522883,
  0.08365168, 0.08430514, 0.08721823, 0.08998087, 0.09195295, 0.09197704, 
    0.08896122, 0.08816623, 0.0864739, 0.08387457, 0.08865711, 0.08927332, 
    0.08395755, 0.0800942, 0.0796309, 0.08085202, 0.08253251, 0.08631988, 
    0.08835641, 0.08807475, 0.08817565, 0.08736547, 0.08621577, 0.08496957, 
    0.08461604, 0.08433731, 0.08230599, 0.07937268, 0.07589479, 0.07376089, 
    0.07308403, 0.07262327, 0.07102428, 0.06920511, 0.06805132, 0.06708571, 
    0.06544543, 0.06378289, 0.06215749, 0.06073443, 0.05969592, 0.05869712, 
    0.05835835, 0.05907122, 0.06047271, 0.06106217, 0.06052856, 0.05898015, 
    0.05366692, 0.04935797, 0.04727486, 0.04660411, 0.04681944, 0.04713327, 
    0.04716725, 0.04621249, 0.04518071, 0.04419871, 0.04323571, 0.04217282, 
    0.04182376, 0.04197012, 0.04201901, 0.04172155, 0.04122837, 0.04089439, 
    0.04056475, 0.04077426, 0.04172809, 0.04201537, 0.0428335, 0.04215064, 
    0.04171728, 0.04012547, 0.03859078, 0.03836259, 0.03875721, 0.03699108, 
    0.03615073, 0.03528289, 0.03493268, 0.03440277, 0.03508503, 0.03742724, 
    0.03926964, 0.03909742, 0.04233207, 0.04662257, 0.04223122, 0.04051685, 
    0.04075518, 0.03627176, 0.03628754, 0.03515654, 0.03841696, 0.03679555, 
    0.03282808, 0.0322493, 0.03502285, 0.03616973, 0.03680069, 0.03756227, 
    0.04178157, 0.03950535, 0.03867592, 0.03903386, 0.03847379, 0.03846612, 
    0.04003646, 0.04789359, 0.04876113, 0.04639984, 0.04639016, 0.04566298, 
    0.04336005, 0.04211893, 0.04262556, 0.04407204, 0.04605467, 0.04748367, 
    0.04858796, 0.0496047, 0.05099504, 0.05292621, 0.05078283, 0.04860774, 
    0.05434711, 0.04611393, 0.0538108, 0.05886478, 0.06164727, 0.06489198, 
    0.06338987, 0.06278989, 0.06364128, 0.06454249, 0.06572505, 0.06652691, 
    0.06743696, 0.06843821, 0.06943804, 0.07066406, 0.07199222, 0.07304645, 
    0.07394802, 0.07502431, 0.07586209, 0.07644499, 0.07697222, 0.07688843, 
    0.07578636, 0.07574085, 0.07597166, 0.07596882, 0.07647904, 0.0769223, 
    0.0773813, 0.07816023, 0.07716476, 0.07786743, 0.09378543, 0.08552954, 
    0.08217067, 0.08415969, 0.08422186, 0.08194506, 0.0768324, 0.07554183, 
    0.07427933, 0.07403339, 0.07438883, 0.07418208, 0.07387087, 0.07484207, 
    0.07609538, 0.07632543, 0.0781322, 0.08186264, 0.08738638, 0.09872351, 
    0.104846, 0.1074337, 0.1136272, 0.1031591, 0.07447159, 0.06138768, 
    0.05021227, 0.04047427, 0.03667699, 0.03226856, 0.02752087, 0.02717946, 
    0.02680198, 0.02703477, 0.02836282, 0.03123736, 0.03256366, 0.0346102, 
    0.0372215, 0.03777343, 0.0391139, 0.0396862, 0.03996991, 0.04054135, 
    0.04126171, 0.04162889, 0.04199564, 0.04262089, 0.04345041, 0.04359183, 
    0.04351983, 0.04347296, 0.04330111, 0.04293658, 0.04271108, 0.04296497, 
    0.04346639, 0.04390458, 0.04643488, 0.04748296, 0.04754734, 0.04718763, 
    0.04678156, 0.04660546, 0.04795232, 0.05020675, 0.05269478, 0.05356352, 
    0.05163306, 0.04969106, 0.04835897, 0.04684612, 0.04668814, 0.04829352, 
    0.04957664, 0.05099399, 0.05083265, 0.052944, 0.05594866, 0.0569107, 
    0.06001618, 0.06340085, 0.06764264, 0.07236367, 0.07650927, 0.07947503, 
    0.0816188, 0.08320437, 0.08446012, 0.08520296, 0.08552337, 0.08608185, 
    0.08690329, 0.08769693, 0.08814593, 0.08862491, 0.08936443, 0.09027798, 
    0.09174691, 0.0935267, 0.09428842, 0.0947076, 0.09530242, 0.09551542, 
    0.09480196, 0.09322508, 0.0915833, 0.09062298, 0.08981054, 0.08955371, 
    0.08976399, 0.09006939, 0.08987315, 0.08938418, 0.08906646, 0.08913144, 
    0.08868905, 0.08846391, 0.08828946, 0.08846972, 0.0917911, 0.09650983, 
    0.1014866, 0.1127044, 0.1266951, 0.1064027, 0.08936699, 0.08250239,
  0.08562378, 0.08758283, 0.09318829, 0.0998242, 0.09911515, 0.09897217, 
    0.09612267, 0.09300485, 0.08791348, 0.08671776, 0.09101409, 0.09310657, 
    0.08680589, 0.07996742, 0.07845721, 0.07839964, 0.07925487, 0.08263423, 
    0.08405557, 0.08530058, 0.0859037, 0.08463506, 0.08218162, 0.08076042, 
    0.08076727, 0.08068465, 0.07966419, 0.07763248, 0.07505047, 0.0728408, 
    0.07167406, 0.07163722, 0.07144821, 0.07042163, 0.07000984, 0.06902646, 
    0.06783377, 0.06618361, 0.06487313, 0.06340748, 0.06259175, 0.06127431, 
    0.05934637, 0.05879435, 0.05852916, 0.06019156, 0.06075861, 0.05979059, 
    0.05334986, 0.05125028, 0.04987175, 0.04881473, 0.04865202, 0.0490658, 
    0.0493088, 0.04937941, 0.04905965, 0.04834846, 0.04740369, 0.04656393, 
    0.04645306, 0.04617832, 0.04585339, 0.0452744, 0.04427518, 0.04343327, 
    0.04255681, 0.0419312, 0.04206856, 0.04199616, 0.04213006, 0.042498, 
    0.04177214, 0.04063658, 0.03888347, 0.03769145, 0.03705556, 0.03536364, 
    0.03492532, 0.03494985, 0.03520129, 0.03467779, 0.03480617, 0.03484364, 
    0.03596928, 0.03713947, 0.03789901, 0.04369232, 0.04448531, 0.04372533, 
    0.04037399, 0.03920013, 0.03829302, 0.03805675, 0.04114005, 0.04107433, 
    0.04253273, 0.04113377, 0.03632456, 0.03637088, 0.03942159, 0.03969376, 
    0.04001185, 0.03879601, 0.03657529, 0.03665664, 0.03468282, 0.03587142, 
    0.03568572, 0.03735708, 0.04403064, 0.04955521, 0.04639578, 0.04510501, 
    0.04490339, 0.04336836, 0.04295755, 0.0442978, 0.04641971, 0.04807292, 
    0.04882856, 0.04947671, 0.04995378, 0.05040827, 0.04821119, 0.04672839, 
    0.04584235, 0.04709381, 0.05397152, 0.05648486, 0.05907832, 0.06512892, 
    0.06374393, 0.06341112, 0.06391826, 0.06493519, 0.06619125, 0.06714276, 
    0.06821627, 0.0694103, 0.07013442, 0.07126993, 0.07263187, 0.07377958, 
    0.07433355, 0.07515164, 0.07559361, 0.0759636, 0.07664005, 0.07640751, 
    0.07571682, 0.07500029, 0.07437164, 0.07398989, 0.07400738, 0.07400378, 
    0.07439277, 0.07559496, 0.07864293, 0.07716849, 0.07858066, 0.08329923, 
    0.08593801, 0.08227148, 0.08834177, 0.08797406, 0.07656261, 0.07265282, 
    0.07260532, 0.07191558, 0.07227298, 0.07219737, 0.07315911, 0.07457813, 
    0.07444719, 0.0790397, 0.08773026, 0.09286628, 0.09979159, 0.107024, 
    0.1068859, 0.1055156, 0.09073713, 0.06494183, 0.050569, 0.04610502, 
    0.037193, 0.03355197, 0.03237241, 0.02885335, 0.02834885, 0.02815356, 
    0.027658, 0.02780679, 0.02840477, 0.03033754, 0.03244793, 0.03517756, 
    0.03882682, 0.03973979, 0.04049786, 0.04144144, 0.04162699, 0.04124268, 
    0.0416229, 0.04170623, 0.04206695, 0.04283625, 0.04276646, 0.04252005, 
    0.04229762, 0.0422461, 0.04270325, 0.04214476, 0.04279888, 0.04442137, 
    0.04546875, 0.04559166, 0.04565581, 0.04559125, 0.04526211, 0.04486402, 
    0.04469715, 0.04516589, 0.04666542, 0.04755914, 0.04882264, 0.05070829, 
    0.04942191, 0.04739359, 0.04620005, 0.0443707, 0.04495471, 0.04660884, 
    0.04873542, 0.05373451, 0.05219647, 0.05229774, 0.05430925, 0.05769418, 
    0.06175817, 0.06487915, 0.06915803, 0.07300512, 0.07504269, 0.07675092, 
    0.07833219, 0.07985104, 0.08117236, 0.08172937, 0.08187678, 0.08302386, 
    0.08415179, 0.08502267, 0.08555741, 0.08614171, 0.08655502, 0.08740798, 
    0.08985871, 0.09187958, 0.09307145, 0.09357762, 0.09383868, 0.09359228, 
    0.09263922, 0.09129453, 0.08996075, 0.08886819, 0.08769708, 0.0873823, 
    0.08779816, 0.08848257, 0.08971442, 0.08977333, 0.08911661, 0.08816597, 
    0.08813263, 0.08845073, 0.08841832, 0.08833785, 0.08976734, 0.09232869, 
    0.09572282, 0.1017758, 0.1101114, 0.09530655, 0.08397558, 0.08279845,
  0.08558648, 0.09175688, 0.1010631, 0.1040928, 0.119693, 0.135701, 0.113777, 
    0.1018923, 0.09368405, 0.08990325, 0.0887619, 0.08674294, 0.08410691, 
    0.07973566, 0.07769106, 0.07858468, 0.07935131, 0.08128519, 0.08141237, 
    0.08224797, 0.0820507, 0.08119615, 0.08080779, 0.07961001, 0.07858887, 
    0.07835858, 0.07801755, 0.07698559, 0.07473659, 0.07260929, 0.07179516, 
    0.07198241, 0.07323764, 0.07373431, 0.07328957, 0.0721576, 0.07126103, 
    0.0689496, 0.067011, 0.0658683, 0.06484666, 0.0630135, 0.06102695, 
    0.05980892, 0.05961788, 0.06038874, 0.06086732, 0.0590484, 0.05432776, 
    0.05230161, 0.05165581, 0.05077773, 0.05009368, 0.05066696, 0.05148301, 
    0.05213366, 0.05235663, 0.05118477, 0.05004814, 0.04912392, 0.04870142, 
    0.04838071, 0.04772225, 0.04683938, 0.04577562, 0.0451032, 0.04459753, 
    0.04424093, 0.04369055, 0.04341948, 0.04350606, 0.04387427, 0.0437674, 
    0.04375986, 0.04278571, 0.04014396, 0.03797307, 0.03646974, 0.03399218, 
    0.03371659, 0.03371475, 0.03434135, 0.03515849, 0.03539166, 0.03449024, 
    0.03382475, 0.033662, 0.03501719, 0.0366771, 0.03870984, 0.0402892, 
    0.0443768, 0.0385429, 0.03563951, 0.03792509, 0.03785376, 0.03859876, 
    0.03760115, 0.03713875, 0.03796184, 0.03851716, 0.03775231, 0.03705337, 
    0.03666424, 0.03482605, 0.03510273, 0.03284088, 0.03450232, 0.03426744, 
    0.03375376, 0.03592098, 0.04267115, 0.04572587, 0.04560009, 0.04448095, 
    0.04373016, 0.04410356, 0.04562708, 0.04816113, 0.04993937, 0.04982711, 
    0.04917328, 0.04711872, 0.04709826, 0.0468914, 0.04546307, 0.04232101, 
    0.04468894, 0.05889814, 0.05534876, 0.05602616, 0.05909089, 0.06211195, 
    0.0621469, 0.0628936, 0.06465855, 0.06662976, 0.06857351, 0.06984158, 
    0.07002115, 0.07119081, 0.07241791, 0.0735569, 0.07428706, 0.07488098, 
    0.07517094, 0.07524034, 0.07532034, 0.07545161, 0.07518916, 0.07450244, 
    0.0739916, 0.07334067, 0.07229504, 0.07185654, 0.0719709, 0.07257879, 
    0.07292357, 0.07508315, 0.07954405, 0.07966142, 0.08012272, 0.08359537, 
    0.08409947, 0.08766808, 0.08473628, 0.08009084, 0.07755895, 0.07564667, 
    0.07453518, 0.07431887, 0.07566483, 0.07865876, 0.08152705, 0.08928839, 
    0.09713441, 0.09522455, 0.1026887, 0.1244676, 0.1147518, 0.09381072, 
    0.08094115, 0.05581068, 0.0459457, 0.03679417, 0.03179466, 0.02962499, 
    0.0306377, 0.03073486, 0.02970643, 0.03011046, 0.02684264, 0.02584281, 
    0.02625506, 0.02838892, 0.02936152, 0.03121203, 0.03219897, 0.0344991, 
    0.03713161, 0.03905366, 0.04015863, 0.04137547, 0.04206702, 0.04202829, 
    0.04191324, 0.0417829, 0.0416613, 0.04106035, 0.04063281, 0.04017816, 
    0.03992468, 0.04025884, 0.04146823, 0.04303304, 0.04372934, 0.04397462, 
    0.04370854, 0.0434081, 0.04340984, 0.043527, 0.04331307, 0.04272123, 
    0.04307755, 0.04372053, 0.04394674, 0.04528402, 0.04613563, 0.04533132, 
    0.04441883, 0.04387576, 0.04260878, 0.04354512, 0.04499075, 0.04684846, 
    0.05108273, 0.05301247, 0.05272231, 0.05389598, 0.0599365, 0.06369951, 
    0.0661185, 0.06935084, 0.07188383, 0.07257196, 0.07309544, 0.07398985, 
    0.07495835, 0.0752601, 0.07654075, 0.07931621, 0.08086191, 0.08224866, 
    0.08462037, 0.08529779, 0.08487111, 0.08484517, 0.08582433, 0.08733324, 
    0.08904658, 0.08998866, 0.0904248, 0.09044854, 0.0901621, 0.0897376, 
    0.08907331, 0.08802914, 0.08685966, 0.08601713, 0.08575071, 0.08602415, 
    0.08699869, 0.08851314, 0.08898304, 0.08883537, 0.08846839, 0.08824211, 
    0.0882315, 0.08796182, 0.08764127, 0.08774632, 0.08833382, 0.08794313, 
    0.08679367, 0.08894005, 0.08588564, 0.08316562, 0.08447142,
  0.08579763, 0.09190141, 0.1045918, 0.1020452, 0.1073495, 0.1354327, 
    0.1219357, 0.1044269, 0.09805439, 0.09517749, 0.09213201, 0.0877369, 
    0.08460202, 0.07968778, 0.07619994, 0.07570423, 0.07731857, 0.07845889, 
    0.07887141, 0.07954737, 0.07994957, 0.07866605, 0.07898791, 0.0794599, 
    0.08006764, 0.07928883, 0.07786541, 0.07673792, 0.07563341, 0.07361657, 
    0.07211553, 0.07282047, 0.07371958, 0.07485828, 0.07461796, 0.07381784, 
    0.0723791, 0.07045563, 0.0688714, 0.06748912, 0.06594694, 0.06410242, 
    0.0628672, 0.06213066, 0.06204199, 0.06424289, 0.06296553, 0.06064541, 
    0.05502673, 0.05302062, 0.05354391, 0.05188942, 0.05152141, 0.0516784, 
    0.05242506, 0.05295989, 0.05303005, 0.05254641, 0.05195618, 0.05112348, 
    0.05008917, 0.0490708, 0.04807842, 0.04712879, 0.04642823, 0.04648525, 
    0.04662243, 0.04651346, 0.04646952, 0.04651865, 0.04672555, 0.04616947, 
    0.04743557, 0.04818987, 0.04727231, 0.04419821, 0.04098849, 0.03730411, 
    0.03554272, 0.03430839, 0.03394379, 0.03454677, 0.03521743, 0.03557321, 
    0.03418079, 0.03291707, 0.03155334, 0.03131297, 0.03239631, 0.03412279, 
    0.03650446, 0.04033211, 0.03826057, 0.0334446, 0.03135392, 0.03138521, 
    0.03202926, 0.03208548, 0.03263772, 0.03322353, 0.03352643, 0.03326278, 
    0.03224724, 0.03094042, 0.02953675, 0.03008718, 0.03054264, 0.03294091, 
    0.03443397, 0.0351686, 0.03510936, 0.03698177, 0.04206135, 0.04493257, 
    0.04421223, 0.04242423, 0.04323979, 0.04567983, 0.04821572, 0.04902688, 
    0.04664427, 0.04819018, 0.04992496, 0.04414933, 0.04442672, 0.04527164, 
    0.0448866, 0.04102106, 0.04446936, 0.07107519, 0.05974232, 0.05304184, 
    0.05545702, 0.05684109, 0.05804424, 0.06019339, 0.06283037, 0.06904658, 
    0.07347719, 0.07242344, 0.07260744, 0.07383689, 0.07594796, 0.0757448, 
    0.07558379, 0.0750998, 0.07413114, 0.07351615, 0.07296815, 0.07253122, 
    0.07238296, 0.07240251, 0.07223953, 0.0708513, 0.06962814, 0.07061386, 
    0.0707416, 0.06886382, 0.07778933, 0.08493998, 0.08246389, 0.08059285, 
    0.07851366, 0.08112174, 0.08796142, 0.08718338, 0.08590186, 0.08602128, 
    0.08980578, 0.08700448, 0.084698, 0.08858592, 0.08995815, 0.09409577, 
    0.1041527, 0.1022169, 0.1048325, 0.1184113, 0.105016, 0.07755233, 
    0.0596903, 0.05030539, 0.04309637, 0.03769303, 0.03272565, 0.02903566, 
    0.02920241, 0.02699654, 0.02842303, 0.02633012, 0.02608553, 0.02509334, 
    0.02581707, 0.02675642, 0.02894744, 0.03085936, 0.03161269, 0.03295973, 
    0.03409513, 0.03526117, 0.03659362, 0.03879008, 0.04002408, 0.04117637, 
    0.04212991, 0.04162557, 0.0408729, 0.04014869, 0.03980584, 0.03949006, 
    0.03931708, 0.03951633, 0.0406525, 0.04192229, 0.042611, 0.04307819, 
    0.0431451, 0.04284005, 0.04249625, 0.04225438, 0.04217429, 0.04216972, 
    0.04185603, 0.04189344, 0.04256396, 0.04233571, 0.04223815, 0.04285237, 
    0.0423962, 0.04261095, 0.04141372, 0.04062106, 0.04136092, 0.04251155, 
    0.04438798, 0.04956654, 0.05634846, 0.05226425, 0.05562858, 0.06209279, 
    0.0641919, 0.06545441, 0.06718324, 0.06854383, 0.06909496, 0.06928568, 
    0.068751, 0.06870313, 0.07276489, 0.07754636, 0.07730529, 0.07831036, 
    0.07973778, 0.08307061, 0.08680768, 0.08743113, 0.08481865, 0.08333779, 
    0.08387157, 0.08490714, 0.08556342, 0.08599351, 0.08647905, 0.08661082, 
    0.08658588, 0.08634859, 0.08598751, 0.08570654, 0.08498614, 0.08487671, 
    0.08576049, 0.08699384, 0.08818888, 0.08819494, 0.08806932, 0.08805011, 
    0.08818515, 0.08793181, 0.08768754, 0.08741749, 0.08715526, 0.08711404, 
    0.08681499, 0.08639284, 0.08659893, 0.08616436, 0.08560626, 0.08445191,
  0.08604755, 0.09208687, 0.09786369, 0.1001682, 0.1103092, 0.1149185, 
    0.106521, 0.09204811, 0.08836354, 0.09228321, 0.08836335, 0.08515882, 
    0.08259666, 0.0768797, 0.0714236, 0.07190995, 0.07280969, 0.07462578, 
    0.07664615, 0.07826348, 0.07837456, 0.07700759, 0.07798015, 0.07894084, 
    0.07911665, 0.07879774, 0.07764971, 0.07668155, 0.07554661, 0.07374921, 
    0.07277532, 0.07380851, 0.07326879, 0.07316894, 0.07240896, 0.07206938, 
    0.07106446, 0.07004848, 0.06947776, 0.06813847, 0.06687611, 0.06527664, 
    0.06438496, 0.06401616, 0.06369431, 0.06451348, 0.0650862, 0.06001518, 
    0.05615514, 0.05470467, 0.05441802, 0.05402888, 0.05344193, 0.05332354, 
    0.0535529, 0.05406542, 0.05407446, 0.05381628, 0.05407435, 0.05331329, 
    0.05204628, 0.05100887, 0.0498174, 0.04893711, 0.04897201, 0.04900488, 
    0.04893345, 0.04872476, 0.0483546, 0.04799618, 0.04765088, 0.04834883, 
    0.04877393, 0.04886268, 0.0479292, 0.04531169, 0.04122766, 0.03916386, 
    0.03748133, 0.03485052, 0.034276, 0.03429897, 0.03459584, 0.03422556, 
    0.0331522, 0.03221153, 0.03131799, 0.03093211, 0.03109434, 0.03140159, 
    0.03213762, 0.03207031, 0.03147631, 0.03159342, 0.03000731, 0.02875398, 
    0.0288296, 0.02952066, 0.02981286, 0.03020441, 0.03016905, 0.02980084, 
    0.02955409, 0.0284533, 0.0276441, 0.02832793, 0.02948979, 0.03182672, 
    0.03415667, 0.03595638, 0.03621944, 0.03571916, 0.0362818, 0.03657279, 
    0.03874461, 0.03892171, 0.03998116, 0.04165545, 0.04245552, 0.04188934, 
    0.04110327, 0.04294147, 0.04653703, 0.04886871, 0.05027917, 0.0479701, 
    0.04627058, 0.0412309, 0.04167829, 0.04219695, 0.04535179, 0.04816968, 
    0.05255916, 0.05327318, 0.05158917, 0.0515308, 0.0565945, 0.06148452, 
    0.0658388, 0.07342126, 0.07398283, 0.07391366, 0.07416803, 0.07440881, 
    0.07420359, 0.07316867, 0.0720138, 0.07113113, 0.07075661, 0.07023805, 
    0.06991053, 0.07011246, 0.06946612, 0.06793065, 0.06776943, 0.06761704, 
    0.06900021, 0.06626223, 0.06315162, 0.07392654, 0.07763883, 0.07559026, 
    0.07083101, 0.07620506, 0.08579976, 0.08680556, 0.08379246, 0.08687434, 
    0.09214094, 0.0911025, 0.1011508, 0.1070404, 0.1003658, 0.1045804, 
    0.1194907, 0.09127211, 0.09191798, 0.06338777, 0.03725251, 0.03780603, 
    0.03717464, 0.03843465, 0.03880139, 0.03386495, 0.03280997, 0.02765657, 
    0.03094194, 0.02871471, 0.02601019, 0.0259132, 0.02510386, 0.02563847, 
    0.02716287, 0.02732719, 0.0290197, 0.03130858, 0.03206987, 0.03260285, 
    0.03350024, 0.03495579, 0.03682096, 0.03874719, 0.0398743, 0.04027304, 
    0.04016327, 0.03993576, 0.03892247, 0.0379497, 0.0375245, 0.03765819, 
    0.0378487, 0.03767802, 0.039207, 0.04092869, 0.04205471, 0.04302962, 
    0.0432505, 0.04277006, 0.04191747, 0.04118442, 0.04087693, 0.04091565, 
    0.04103026, 0.04097597, 0.04096926, 0.04038828, 0.04082871, 0.04057906, 
    0.04024175, 0.03995979, 0.03872767, 0.03994888, 0.04137748, 0.04253466, 
    0.0426458, 0.04355485, 0.04599809, 0.04866658, 0.05487301, 0.06058154, 
    0.06169, 0.06262103, 0.06342182, 0.06348541, 0.06261426, 0.06128397, 
    0.06258118, 0.06798871, 0.07156651, 0.06861465, 0.06408431, 0.05615124, 
    0.06621058, 0.07820566, 0.07582357, 0.08825218, 0.08666583, 0.08185729, 
    0.0815944, 0.08207753, 0.082158, 0.08229721, 0.08264332, 0.08326839, 
    0.08373971, 0.08396468, 0.08439706, 0.08460865, 0.08401398, 0.08452795, 
    0.08588892, 0.08691567, 0.08817252, 0.08930773, 0.08944788, 0.08971369, 
    0.08987305, 0.08972759, 0.08970872, 0.08943818, 0.08854781, 0.08801632, 
    0.08769902, 0.08753661, 0.08728472, 0.08672567, 0.08599417, 0.08472349,
  0.08439524, 0.08888623, 0.09094735, 0.08883715, 0.09608783, 0.09908669, 
    0.08728772, 0.07670029, 0.07560642, 0.07840592, 0.07787655, 0.07714932, 
    0.07493254, 0.070466, 0.06821316, 0.06870396, 0.06943255, 0.07130225, 
    0.07492372, 0.07664397, 0.07684621, 0.07714295, 0.07726534, 0.07688913, 
    0.07630344, 0.07510915, 0.07435262, 0.07238164, 0.07120032, 0.07117874, 
    0.07069957, 0.07151338, 0.0690706, 0.06934364, 0.06877082, 0.06829192, 
    0.06815477, 0.06788244, 0.06793621, 0.06654698, 0.06494452, 0.06335771, 
    0.06261551, 0.06323349, 0.06306957, 0.06340025, 0.06251818, 0.05900085, 
    0.05557974, 0.05414993, 0.05571654, 0.05528421, 0.05434933, 0.05407233, 
    0.05330013, 0.05266232, 0.0526869, 0.05266153, 0.05272333, 0.05250924, 
    0.05208331, 0.05122886, 0.05070908, 0.05047109, 0.05104497, 0.0509399, 
    0.05049094, 0.04944846, 0.0487497, 0.04819376, 0.04771777, 0.04733318, 
    0.04688849, 0.04758571, 0.04690794, 0.0440882, 0.04235945, 0.04060721, 
    0.0363448, 0.03468459, 0.03405022, 0.03398647, 0.0339699, 0.03316217, 
    0.03262268, 0.03163863, 0.03139687, 0.03119254, 0.03059204, 0.03027602, 
    0.02979166, 0.02938226, 0.02884289, 0.02857928, 0.02831707, 0.02791335, 
    0.0283146, 0.02843664, 0.02850596, 0.02795138, 0.02751096, 0.02727094, 
    0.02689286, 0.02683681, 0.02582788, 0.02663152, 0.02799639, 0.0301951, 
    0.03328249, 0.0356807, 0.03592872, 0.03502915, 0.03334503, 0.0335698, 
    0.03435908, 0.03125382, 0.03085737, 0.03094676, 0.03306959, 0.03500614, 
    0.03578799, 0.03686289, 0.03601272, 0.04025441, 0.04545437, 0.04844015, 
    0.04532269, 0.04227245, 0.04599345, 0.04770447, 0.04155795, 0.04166285, 
    0.04214517, 0.04009159, 0.04015297, 0.04303702, 0.05418851, 0.0569884, 
    0.05818513, 0.06098365, 0.063978, 0.06654793, 0.06689403, 0.06858564, 
    0.07063617, 0.07034048, 0.06926829, 0.06777068, 0.06723235, 0.06699743, 
    0.06704821, 0.06642877, 0.06556418, 0.06371395, 0.06185032, 0.05959666, 
    0.06035709, 0.06316435, 0.05991089, 0.05675553, 0.06110293, 0.06172698, 
    0.05411451, 0.05450759, 0.06610275, 0.07617877, 0.07390898, 0.06653704, 
    0.07594068, 0.08061948, 0.08922125, 0.07808331, 0.06099841, 0.05374635, 
    0.04469845, 0.03927993, 0.02936066, 0.02668611, 0.02756302, 0.02798375, 
    0.03086649, 0.03350539, 0.03614622, 0.03399591, 0.0360977, 0.03546283, 
    0.03287987, 0.02905139, 0.02693708, 0.02953096, 0.0286474, 0.02730638, 
    0.02705675, 0.02871732, 0.02963488, 0.03207326, 0.03389055, 0.03313336, 
    0.03320203, 0.03386888, 0.0354853, 0.036913, 0.03764101, 0.03787781, 
    0.03765232, 0.03666316, 0.03611556, 0.03580904, 0.03604289, 0.03646883, 
    0.03692846, 0.03682113, 0.03758292, 0.03874991, 0.04070726, 0.04162624, 
    0.04154054, 0.04071584, 0.0395892, 0.03888797, 0.03828472, 0.03809507, 
    0.03889006, 0.03936432, 0.03881705, 0.03853027, 0.03872822, 0.03849889, 
    0.03973296, 0.04215915, 0.04231895, 0.04117234, 0.04051291, 0.03964286, 
    0.04051375, 0.03978566, 0.04164639, 0.04520528, 0.05005578, 0.05383458, 
    0.05670063, 0.05850337, 0.05862606, 0.05668507, 0.05528459, 0.05763457, 
    0.06123639, 0.05955897, 0.05571868, 0.04983721, 0.04199096, 0.04428343, 
    0.06546114, 0.08531494, 0.07401775, 0.08551242, 0.08830746, 0.08236137, 
    0.07888826, 0.07990149, 0.08021481, 0.08050486, 0.08069827, 0.08110084, 
    0.08173072, 0.08233505, 0.08330457, 0.08343285, 0.08345245, 0.08373243, 
    0.08516522, 0.08687933, 0.08862387, 0.0895211, 0.08944977, 0.09012172, 
    0.09061608, 0.09164152, 0.09195022, 0.0919906, 0.09070679, 0.09012187, 
    0.08974434, 0.09016192, 0.08925841, 0.08764072, 0.08589526, 0.08445893,
  0.08088534, 0.08155236, 0.08262568, 0.07669964, 0.07554161, 0.08658136, 
    0.07828043, 0.06846619, 0.06835095, 0.06651165, 0.06730387, 0.06678574, 
    0.06866708, 0.06812835, 0.06499805, 0.06518961, 0.0661348, 0.06822845, 
    0.07125522, 0.07220364, 0.07235163, 0.07389797, 0.07457123, 0.07401767, 
    0.07359235, 0.07186878, 0.07047423, 0.0691903, 0.06888448, 0.06877051, 
    0.0676337, 0.06799804, 0.06731205, 0.0672249, 0.0670701, 0.06656917, 
    0.06710285, 0.06705946, 0.06595335, 0.06438436, 0.06274964, 0.06135891, 
    0.06071176, 0.06070487, 0.05972904, 0.05920021, 0.05942304, 0.05686341, 
    0.05366427, 0.05132617, 0.05128859, 0.05340114, 0.0533214, 0.05281517, 
    0.05264669, 0.05196649, 0.05164631, 0.05133895, 0.05104425, 0.05084036, 
    0.0508742, 0.0513003, 0.05102575, 0.05082669, 0.05155335, 0.05063171, 
    0.04909182, 0.04831803, 0.04739433, 0.04663837, 0.04704896, 0.04731228, 
    0.0466488, 0.04622943, 0.04555472, 0.04360212, 0.04140373, 0.03790807, 
    0.03582267, 0.03438799, 0.03347123, 0.03286509, 0.03180633, 0.03133985, 
    0.03145159, 0.03114435, 0.03148961, 0.03084903, 0.03039118, 0.02958667, 
    0.02857717, 0.02846972, 0.02730952, 0.0269728, 0.02663392, 0.02693294, 
    0.02786127, 0.02757532, 0.02794809, 0.02785213, 0.02762985, 0.02728592, 
    0.02629156, 0.02640706, 0.02582649, 0.02610164, 0.02734424, 0.02926454, 
    0.03205512, 0.03377454, 0.03318868, 0.03223801, 0.03014093, 0.02563937, 
    0.02558883, 0.02435955, 0.02547524, 0.02703436, 0.02680949, 0.03058432, 
    0.03281584, 0.03320323, 0.03351056, 0.03140032, 0.0335235, 0.0382416, 
    0.04108281, 0.04153366, 0.041728, 0.04167894, 0.04071781, 0.04012886, 
    0.03920161, 0.03769974, 0.03594168, 0.03716585, 0.04429357, 0.04700583, 
    0.04836314, 0.04994839, 0.05171809, 0.05316331, 0.05703557, 0.0608279, 
    0.06521863, 0.06582829, 0.06484938, 0.06389871, 0.06371436, 0.06408351, 
    0.06409429, 0.06263873, 0.06134838, 0.05961275, 0.0580522, 0.05625703, 
    0.05372042, 0.05505926, 0.05864367, 0.05596445, 0.05140118, 0.05150389, 
    0.05152627, 0.04630208, 0.03975448, 0.05583578, 0.067235, 0.05998649, 
    0.05396952, 0.04922492, 0.04097929, 0.04381253, 0.04500191, 0.03921821, 
    0.03372251, 0.0329853, 0.0331371, 0.0323691, 0.02864796, 0.0283848, 
    0.03015561, 0.0331745, 0.03417487, 0.03404937, 0.0371771, 0.03822235, 
    0.02995933, 0.02834184, 0.03307089, 0.03320139, 0.02905111, 0.02777226, 
    0.02715327, 0.02911817, 0.03141113, 0.03191134, 0.03264838, 0.03250641, 
    0.03308794, 0.0333656, 0.03377771, 0.03442809, 0.03499329, 0.03436126, 
    0.03396839, 0.03405505, 0.03390051, 0.03412619, 0.03533686, 0.0354869, 
    0.03540492, 0.03636329, 0.03669744, 0.03667853, 0.03798339, 0.03888614, 
    0.03898042, 0.03837125, 0.0374435, 0.03699133, 0.03654094, 0.03537004, 
    0.03648787, 0.03843666, 0.03819082, 0.0378961, 0.03863829, 0.03908739, 
    0.03958932, 0.04029399, 0.03954601, 0.03973993, 0.03966825, 0.04100934, 
    0.04214347, 0.03868571, 0.03916759, 0.04126995, 0.04501457, 0.04895753, 
    0.05183424, 0.05363773, 0.05337472, 0.05238552, 0.05295597, 0.05357144, 
    0.0510021, 0.04589442, 0.04261533, 0.03509408, 0.02835687, 0.03106749, 
    0.04193233, 0.06648725, 0.07186922, 0.07995006, 0.08779731, 0.08413155, 
    0.07959067, 0.07890189, 0.07998231, 0.08015718, 0.07984896, 0.08029684, 
    0.08077141, 0.08121984, 0.08114294, 0.08080872, 0.08195854, 0.08391593, 
    0.08656358, 0.08966542, 0.09318583, 0.09500329, 0.0963825, 0.09654339, 
    0.09598068, 0.0936446, 0.09202027, 0.09066532, 0.09090634, 0.0909244, 
    0.09108223, 0.09029825, 0.08895508, 0.08687542, 0.08515044, 0.08336937,
  0.07714528, 0.07486928, 0.073012, 0.07005376, 0.06890542, 0.06759936, 
    0.06638341, 0.06767563, 0.06837054, 0.06906851, 0.06961418, 0.0641094, 
    0.06224274, 0.06715725, 0.06704681, 0.06407525, 0.06289926, 0.06198476, 
    0.06322701, 0.0657798, 0.06746743, 0.06984863, 0.07039534, 0.0701285, 
    0.06956661, 0.06766102, 0.06612472, 0.06492005, 0.06478649, 0.06497411, 
    0.06404266, 0.06472215, 0.06480155, 0.06516827, 0.06589131, 0.0660599, 
    0.06608306, 0.06550714, 0.0646221, 0.0635292, 0.06193755, 0.06087011, 
    0.05969432, 0.05850101, 0.05817851, 0.05872908, 0.05669674, 0.05173114, 
    0.05067281, 0.04848887, 0.0474103, 0.04833949, 0.04932999, 0.04985448, 
    0.05045441, 0.05062689, 0.05018133, 0.04977418, 0.04972154, 0.05057926, 
    0.05082271, 0.05080741, 0.05047674, 0.05008745, 0.04937004, 0.04849729, 
    0.04722569, 0.04548788, 0.04468081, 0.04533511, 0.04639949, 0.04791699, 
    0.04649972, 0.04425439, 0.04267384, 0.0407418, 0.03844415, 0.03659356, 
    0.03533278, 0.03410202, 0.03325966, 0.03273102, 0.03219555, 0.03149249, 
    0.03144566, 0.03192099, 0.03189684, 0.03116123, 0.03088151, 0.02992753, 
    0.02928753, 0.0287048, 0.02747762, 0.02691023, 0.02590007, 0.02522811, 
    0.02512459, 0.02517613, 0.02657392, 0.02714409, 0.02762795, 0.02790901, 
    0.02747058, 0.02711675, 0.02790486, 0.02852745, 0.02901538, 0.03170155, 
    0.03152168, 0.03072975, 0.02972811, 0.02762686, 0.02729893, 0.0229717, 
    0.02107132, 0.02171957, 0.02230509, 0.02644411, 0.02852863, 0.03093486, 
    0.03205273, 0.03092459, 0.03059251, 0.03053252, 0.02765059, 0.02928953, 
    0.0348529, 0.03554954, 0.03573732, 0.03713875, 0.03797406, 0.0366955, 
    0.03627749, 0.03592337, 0.03712511, 0.03874188, 0.03896369, 0.03989819, 
    0.04036982, 0.04240716, 0.0447114, 0.04830306, 0.05125204, 0.05463101, 
    0.05776411, 0.05952377, 0.05867409, 0.05809473, 0.05780536, 0.06032344, 
    0.06250122, 0.06148784, 0.05994404, 0.05715864, 0.05484803, 0.05380626, 
    0.05184059, 0.0482565, 0.04914838, 0.05319357, 0.04990446, 0.04331117, 
    0.04323855, 0.04541555, 0.04070402, 0.03877646, 0.04045317, 0.03937929, 
    0.03502274, 0.03472319, 0.03305394, 0.03552528, 0.03290956, 0.02736111, 
    0.03085301, 0.0286726, 0.02910682, 0.02701264, 0.02627807, 0.03207596, 
    0.03350706, 0.03384845, 0.03579052, 0.04076302, 0.03872814, 0.0303163, 
    0.02763651, 0.03318188, 0.03464359, 0.03328022, 0.03058686, 0.02775629, 
    0.02916921, 0.03079964, 0.0314947, 0.03222731, 0.0332045, 0.03324487, 
    0.03318778, 0.03296166, 0.03250789, 0.03228376, 0.03201336, 0.03215086, 
    0.03203204, 0.03200472, 0.03310538, 0.03422953, 0.03492715, 0.03565378, 
    0.03621732, 0.03627022, 0.03635175, 0.03639812, 0.03649227, 0.03670857, 
    0.03713662, 0.03705144, 0.03560825, 0.03469545, 0.03378327, 0.03477919, 
    0.03560569, 0.03714581, 0.03758901, 0.03619974, 0.03558463, 0.03628272, 
    0.03698931, 0.03807738, 0.03822871, 0.03661765, 0.03421087, 0.03372652, 
    0.03612661, 0.03899596, 0.03863847, 0.03797546, 0.04001775, 0.04384126, 
    0.04671722, 0.04836739, 0.04864896, 0.04892801, 0.04964976, 0.04886829, 
    0.04436172, 0.03889043, 0.0326017, 0.02225773, 0.01479694, 0.01718678, 
    0.02489968, 0.04965189, 0.06674615, 0.07134541, 0.08293698, 0.08485703, 
    0.08259621, 0.08083567, 0.08128904, 0.08191489, 0.08176041, 0.0813206, 
    0.08003905, 0.07948279, 0.07933379, 0.0795627, 0.08108171, 0.0823883, 
    0.08468495, 0.09202263, 0.09936297, 0.103266, 0.102314, 0.1012097, 
    0.09863207, 0.09772138, 0.09285755, 0.08981015, 0.08909407, 0.08876652, 
    0.08882106, 0.08871631, 0.08761463, 0.08522984, 0.08292863, 0.08031828,
  0.07466579, 0.07199614, 0.06826572, 0.06435532, 0.06249203, 0.06172044, 
    0.06241614, 0.06354471, 0.06534534, 0.06950305, 0.08179868, 0.07998825, 
    0.06546767, 0.06164889, 0.06444418, 0.06414521, 0.06123744, 0.0588983, 
    0.0583323, 0.05943865, 0.06269305, 0.06605916, 0.06723712, 0.06691801, 
    0.06575745, 0.06378788, 0.06197444, 0.06011444, 0.05896351, 0.05909976, 
    0.0600214, 0.06147471, 0.06249935, 0.06354398, 0.06346282, 0.06328206, 
    0.06292841, 0.06290415, 0.06263024, 0.06197727, 0.06041531, 0.05888411, 
    0.05747889, 0.05692065, 0.05688982, 0.05771067, 0.06340821, 0.05747756, 
    0.05017471, 0.04901661, 0.04582186, 0.04583762, 0.04797497, 0.04858575, 
    0.04917919, 0.0500399, 0.04991178, 0.04884206, 0.04885247, 0.04943431, 
    0.04927581, 0.04877929, 0.04779652, 0.04713246, 0.0474745, 0.04653137, 
    0.04499393, 0.04448266, 0.04429571, 0.04390718, 0.04458665, 0.04668245, 
    0.04565112, 0.0429249, 0.04115882, 0.0394443, 0.03735498, 0.03552664, 
    0.0341961, 0.03285095, 0.03332748, 0.03377249, 0.03351667, 0.03324479, 
    0.03301628, 0.03297171, 0.0322369, 0.03166175, 0.03138614, 0.03078583, 
    0.02978641, 0.02863679, 0.02740285, 0.02641885, 0.02541035, 0.02494698, 
    0.0244588, 0.02407279, 0.02533709, 0.02655781, 0.02805652, 0.02956552, 
    0.03048518, 0.03000933, 0.03050557, 0.03123454, 0.03063148, 0.02936673, 
    0.02607374, 0.02415486, 0.02336616, 0.02225936, 0.02130949, 0.0202105, 
    0.02062487, 0.02213648, 0.02397598, 0.02702244, 0.03019634, 0.03093623, 
    0.03031215, 0.02903854, 0.02671269, 0.02651405, 0.02711762, 0.0284317, 
    0.03012913, 0.02895842, 0.02853259, 0.02983967, 0.03046342, 0.03138154, 
    0.03266563, 0.0341456, 0.03509402, 0.03595066, 0.03734058, 0.03749907, 
    0.03724762, 0.03736774, 0.03851265, 0.04056077, 0.04359913, 0.04801191, 
    0.05107658, 0.05250508, 0.05188876, 0.05073769, 0.0533943, 0.05628093, 
    0.05808975, 0.05817187, 0.05799473, 0.05610912, 0.05082159, 0.05019572, 
    0.05271691, 0.05181671, 0.04477418, 0.0446963, 0.0458964, 0.04293454, 
    0.04170727, 0.03986649, 0.03946519, 0.04045679, 0.03780753, 0.0371401, 
    0.03571195, 0.03266769, 0.03007543, 0.02987947, 0.02973434, 0.02921538, 
    0.03026021, 0.02563193, 0.02527563, 0.03042585, 0.03325181, 0.03388709, 
    0.03437655, 0.03655742, 0.03844488, 0.04014847, 0.03186434, 0.02746959, 
    0.03343137, 0.03493676, 0.03093353, 0.02855094, 0.02819615, 0.0286851, 
    0.03189426, 0.03321308, 0.03292923, 0.03357024, 0.03400248, 0.03367162, 
    0.03310145, 0.03290046, 0.03250065, 0.03229649, 0.03191491, 0.03128563, 
    0.03156894, 0.03226718, 0.03242202, 0.03308809, 0.03505212, 0.03556526, 
    0.03554741, 0.03622794, 0.03668181, 0.03629386, 0.03611883, 0.03615921, 
    0.0360781, 0.0355815, 0.03454723, 0.03405995, 0.03621414, 0.0375283, 
    0.03563237, 0.03523015, 0.03527018, 0.03436362, 0.0324747, 0.03208241, 
    0.03288581, 0.03329537, 0.0328011, 0.03238965, 0.03307611, 0.03771835, 
    0.04474813, 0.04242894, 0.03752517, 0.03817422, 0.03728204, 0.03895957, 
    0.04166593, 0.04479254, 0.04711805, 0.04695205, 0.04288969, 0.03874482, 
    0.03702407, 0.03520407, 0.02915335, 0.0206094, 0.01422705, 0.01518632, 
    0.02110503, 0.03575141, 0.05999089, 0.06551054, 0.07398786, 0.08046754, 
    0.08092867, 0.08118497, 0.08281176, 0.08368181, 0.08288341, 0.08214873, 
    0.07983064, 0.07819336, 0.0759264, 0.0716237, 0.06949329, 0.07147475, 
    0.07484376, 0.0838448, 0.09318634, 0.1098116, 0.1171719, 0.1162677, 
    0.1057948, 0.09231445, 0.08982077, 0.08830678, 0.0847308, 0.08488902, 
    0.08644539, 0.08672751, 0.08597522, 0.08414465, 0.08158863, 0.07778782,
  0.07515094, 0.07190193, 0.06854692, 0.06474854, 0.06249017, 0.06063208, 
    0.06107197, 0.06241978, 0.0642035, 0.06668378, 0.0738993, 0.08484171, 
    0.08012901, 0.06384908, 0.05815141, 0.06134326, 0.06179832, 0.05881931, 
    0.05748689, 0.05834016, 0.06129178, 0.06480528, 0.06615417, 0.065078, 
    0.0632062, 0.06147988, 0.05914079, 0.05732634, 0.05654537, 0.05677679, 
    0.05824682, 0.05915895, 0.06093127, 0.06273947, 0.06219807, 0.06110924, 
    0.0607421, 0.06135043, 0.06061595, 0.05933013, 0.0574337, 0.05479594, 
    0.05418881, 0.05516608, 0.05608748, 0.05420412, 0.0550118, 0.05540431, 
    0.05068976, 0.04988905, 0.04993208, 0.04702329, 0.0467562, 0.04717379, 
    0.04830427, 0.05002109, 0.04961582, 0.04845868, 0.04834647, 0.04839715, 
    0.04757644, 0.04668387, 0.04571214, 0.04520339, 0.04474206, 0.04447166, 
    0.04432261, 0.04346389, 0.04266635, 0.04274802, 0.04326703, 0.04430836, 
    0.04431098, 0.04298086, 0.04127045, 0.03894376, 0.03697016, 0.03539176, 
    0.03389699, 0.03236476, 0.03256072, 0.03266007, 0.03265626, 0.03274334, 
    0.03215038, 0.03210622, 0.03164178, 0.03095135, 0.03098116, 0.03085282, 
    0.03003929, 0.02905791, 0.02779979, 0.02682158, 0.02611572, 0.02564784, 
    0.02542529, 0.02549166, 0.02599556, 0.02689727, 0.02807588, 0.02991519, 
    0.033119, 0.03153165, 0.0295399, 0.02928684, 0.02703273, 0.02482794, 
    0.0235962, 0.02276509, 0.02156097, 0.02191235, 0.02237141, 0.0199551, 
    0.02099155, 0.02388912, 0.02527251, 0.03210498, 0.03376069, 0.02907337, 
    0.02750238, 0.02616215, 0.02493191, 0.02518519, 0.02583569, 0.02701042, 
    0.02729725, 0.02675945, 0.02733205, 0.02858368, 0.02855211, 0.02886212, 
    0.03075052, 0.03242201, 0.03253079, 0.03304981, 0.03320952, 0.03346574, 
    0.03342772, 0.03426619, 0.03596795, 0.03776629, 0.04010667, 0.04222878, 
    0.04418299, 0.04631133, 0.04741469, 0.04588372, 0.04729645, 0.05218226, 
    0.05474847, 0.05339008, 0.05224685, 0.05104471, 0.04900008, 0.04719947, 
    0.04621209, 0.0455007, 0.0429537, 0.0441308, 0.04272894, 0.04186291, 
    0.04220659, 0.03956069, 0.039458, 0.04021677, 0.03847475, 0.03774134, 
    0.03568916, 0.03333073, 0.03262447, 0.03258034, 0.03113344, 0.02865505, 
    0.02842424, 0.02782005, 0.03029271, 0.03375601, 0.03137391, 0.03040732, 
    0.03329055, 0.03457023, 0.03606956, 0.03607589, 0.03424032, 0.03408358, 
    0.03363966, 0.03074547, 0.02927219, 0.02905336, 0.02935356, 0.03113125, 
    0.0318099, 0.03123691, 0.03191271, 0.03366264, 0.03425059, 0.03386221, 
    0.03377577, 0.03368718, 0.03313811, 0.03250282, 0.03239784, 0.03256402, 
    0.03241561, 0.03257478, 0.0333125, 0.0339784, 0.03456654, 0.03511818, 
    0.03562162, 0.03632259, 0.03684083, 0.03655569, 0.03569448, 0.03520609, 
    0.03458034, 0.0332095, 0.03211156, 0.03152682, 0.03169451, 0.03270938, 
    0.03285985, 0.03282871, 0.03240599, 0.03065584, 0.02961497, 0.02940361, 
    0.03004286, 0.03034222, 0.03083571, 0.0323006, 0.03328381, 0.03339016, 
    0.03186524, 0.03169617, 0.03665783, 0.03876168, 0.03369986, 0.0329053, 
    0.03755975, 0.04274218, 0.04474514, 0.0402841, 0.03633397, 0.03329741, 
    0.02939975, 0.02724483, 0.02475763, 0.02041882, 0.01423569, 0.01374065, 
    0.02004217, 0.02964237, 0.04152318, 0.04775349, 0.05330804, 0.055888, 
    0.06014508, 0.06396496, 0.07245217, 0.08331298, 0.08714131, 0.08245636, 
    0.08123185, 0.07980842, 0.07855628, 0.07010143, 0.07060368, 0.08069997, 
    0.0766516, 0.06805718, 0.07077263, 0.07540306, 0.0840954, 0.09009045, 
    0.08898032, 0.08573845, 0.08272601, 0.0814623, 0.08119459, 0.08194327, 
    0.08375277, 0.08470691, 0.08484425, 0.08433843, 0.08244129, 0.07884102,
  0.07647, 0.07325453, 0.07007048, 0.06716159, 0.06513029, 0.0644237, 
    0.06509975, 0.06531065, 0.06567465, 0.06683441, 0.06969291, 0.07414152, 
    0.08211958, 0.07815298, 0.06100625, 0.0540256, 0.05762003, 0.05969595, 
    0.05942144, 0.05999215, 0.06141796, 0.06397236, 0.06511876, 0.06327953, 
    0.06196959, 0.06062083, 0.05881366, 0.057911, 0.05767747, 0.05849554, 
    0.0605534, 0.05996621, 0.05742459, 0.05516423, 0.05638669, 0.05827819, 
    0.05877448, 0.0590709, 0.05868427, 0.05759325, 0.05502316, 0.05337385, 
    0.05273528, 0.05262631, 0.05338847, 0.05365457, 0.05274529, 0.05252274, 
    0.05066567, 0.04819648, 0.04689124, 0.04549727, 0.04746982, 0.04849543, 
    0.04662612, 0.04615655, 0.04644456, 0.04600979, 0.04521969, 0.04470146, 
    0.04430655, 0.04392502, 0.0433706, 0.04324618, 0.0440363, 0.04382088, 
    0.04289912, 0.04242519, 0.04210466, 0.04238034, 0.04327296, 0.04368648, 
    0.04330581, 0.04230146, 0.04068436, 0.03835407, 0.03582943, 0.03462465, 
    0.0338625, 0.03276784, 0.03166439, 0.03138441, 0.03220832, 0.03120513, 
    0.03034023, 0.03054235, 0.02993405, 0.02959585, 0.02995029, 0.02936881, 
    0.02918276, 0.02959445, 0.02896515, 0.02822209, 0.02775882, 0.02700258, 
    0.02687173, 0.02701962, 0.02709385, 0.02805334, 0.02857648, 0.02886418, 
    0.02891761, 0.02807601, 0.02705943, 0.02749649, 0.0260952, 0.02458864, 
    0.02338076, 0.02201027, 0.0214192, 0.02257839, 0.02753951, 0.02759324, 
    0.02558053, 0.02752545, 0.02785732, 0.02696699, 0.02800018, 0.02656724, 
    0.02513862, 0.02517872, 0.02472601, 0.0242722, 0.02518246, 0.02589147, 
    0.02572676, 0.02561498, 0.02606531, 0.02644567, 0.02580492, 0.02583895, 
    0.02662289, 0.0279153, 0.02947139, 0.03021456, 0.031691, 0.03170508, 
    0.03131109, 0.03186141, 0.03256793, 0.03386538, 0.03531628, 0.0377609, 
    0.04196574, 0.04615902, 0.05015508, 0.05007522, 0.04854121, 0.05161134, 
    0.05361538, 0.05069338, 0.04744218, 0.04555333, 0.04366317, 0.0415886, 
    0.03957843, 0.03975213, 0.04106024, 0.0414267, 0.04068735, 0.0433699, 
    0.04495497, 0.04464851, 0.04710948, 0.04410309, 0.04098567, 0.04276112, 
    0.03935646, 0.03714932, 0.03707227, 0.03414968, 0.03152542, 0.0306228, 
    0.03234515, 0.0320298, 0.03088516, 0.03176436, 0.0320027, 0.03488329, 
    0.03787276, 0.03416247, 0.03247162, 0.03212782, 0.02885671, 0.02849543, 
    0.0287798, 0.02808772, 0.02886846, 0.02972808, 0.03006048, 0.03076752, 
    0.03012271, 0.02980489, 0.03115243, 0.03229458, 0.03299179, 0.03327889, 
    0.03422078, 0.03409687, 0.03240773, 0.0316016, 0.03178613, 0.03206017, 
    0.03219026, 0.03239439, 0.03256169, 0.03288956, 0.03296899, 0.0333917, 
    0.03391179, 0.03465982, 0.0357413, 0.03547937, 0.03436621, 0.03383106, 
    0.03281124, 0.03140079, 0.02972259, 0.02880655, 0.02841536, 0.02877907, 
    0.02907551, 0.0293388, 0.02984849, 0.02942053, 0.02895694, 0.0286091, 
    0.02872317, 0.0285835, 0.02923845, 0.02950164, 0.02907367, 0.02903883, 
    0.02877302, 0.02985292, 0.03281068, 0.03403958, 0.03193923, 0.03039101, 
    0.03363305, 0.03838896, 0.04055615, 0.03759882, 0.0338425, 0.03059661, 
    0.02394015, 0.02100247, 0.01995345, 0.01695195, 0.01356213, 0.01249788, 
    0.01513374, 0.01671397, 0.01940475, 0.02323519, 0.02869279, 0.03170567, 
    0.03273294, 0.04359007, 0.05623981, 0.05584399, 0.0734312, 0.07866289, 
    0.07995783, 0.0782982, 0.07690234, 0.0751481, 0.07499284, 0.07633841, 
    0.07464331, 0.06976904, 0.06933443, 0.07102117, 0.07361378, 0.07542875, 
    0.07523154, 0.07445539, 0.0748485, 0.07516793, 0.0772235, 0.07862075, 
    0.08073819, 0.08219187, 0.08355621, 0.08379861, 0.08290367, 0.08039959,
  0.07816631, 0.0758271, 0.07329971, 0.07101642, 0.06831919, 0.06677577, 
    0.06660675, 0.06641231, 0.06600301, 0.06660631, 0.0651484, 0.06354662, 
    0.06967019, 0.07935978, 0.07623563, 0.06196807, 0.05282186, 0.05226465, 
    0.0557522, 0.05691714, 0.05831437, 0.06042136, 0.06147178, 0.06088474, 
    0.06094139, 0.06087163, 0.06066509, 0.06087829, 0.06100773, 0.06065496, 
    0.05960479, 0.05857185, 0.05772122, 0.05539118, 0.05509563, 0.05617448, 
    0.05655626, 0.05684303, 0.05693755, 0.05685977, 0.05580056, 0.05369237, 
    0.05259147, 0.05201103, 0.05171136, 0.05232505, 0.05214824, 0.0509063, 
    0.04983708, 0.04905768, 0.04986421, 0.04881146, 0.04499288, 0.04479497, 
    0.04472816, 0.04388012, 0.04390633, 0.04320433, 0.04164066, 0.04097526, 
    0.0409653, 0.04091748, 0.04128503, 0.04147342, 0.04214004, 0.04207291, 
    0.04117862, 0.04107446, 0.04168257, 0.04200903, 0.04280426, 0.04243101, 
    0.04115473, 0.03983688, 0.03808878, 0.03613143, 0.03432626, 0.03254168, 
    0.0314143, 0.0309217, 0.03022629, 0.03005962, 0.02938562, 0.02840061, 
    0.02849342, 0.02825216, 0.02739976, 0.02767518, 0.02779502, 0.02751913, 
    0.02837397, 0.02889958, 0.02896538, 0.02874231, 0.02820807, 0.02754833, 
    0.02706044, 0.02691967, 0.02723618, 0.02800351, 0.02991675, 0.03120035, 
    0.02831326, 0.02584938, 0.02528581, 0.02474035, 0.02433464, 0.02351516, 
    0.0220412, 0.02184678, 0.02335676, 0.02421947, 0.02658778, 0.0300422, 
    0.02867601, 0.02786089, 0.02886842, 0.0255979, 0.02345114, 0.02382657, 
    0.02346285, 0.02320176, 0.02406921, 0.02433776, 0.02459214, 0.02471838, 
    0.02448778, 0.02430592, 0.02393304, 0.02395754, 0.02375208, 0.02440103, 
    0.02504519, 0.02604774, 0.02971165, 0.03037926, 0.02825238, 0.02807247, 
    0.02701313, 0.02791552, 0.03166509, 0.03385802, 0.03336487, 0.03534729, 
    0.04127279, 0.04418164, 0.04334873, 0.04273765, 0.04522385, 0.04626827, 
    0.0460494, 0.04547763, 0.04465275, 0.04339487, 0.04163367, 0.03984542, 
    0.03935418, 0.04374051, 0.04648782, 0.04186712, 0.04034907, 0.04327684, 
    0.04272393, 0.04398372, 0.0479342, 0.04630484, 0.04539721, 0.0492172, 
    0.04697399, 0.04323059, 0.04154687, 0.03998497, 0.03709694, 0.033679, 
    0.0330492, 0.0319389, 0.03107175, 0.03226798, 0.03294397, 0.03197416, 
    0.02933336, 0.02751192, 0.02647365, 0.02632798, 0.0262305, 0.02636981, 
    0.02740828, 0.02873669, 0.02913847, 0.02841087, 0.02852151, 0.03009037, 
    0.03054732, 0.03128125, 0.03232146, 0.03219781, 0.03210745, 0.03148669, 
    0.03068465, 0.03034901, 0.02897712, 0.02870594, 0.02928253, 0.02955638, 
    0.02990114, 0.03015989, 0.03040924, 0.03068706, 0.03106275, 0.03144329, 
    0.03192828, 0.03248222, 0.03352187, 0.03346547, 0.03300007, 0.03221, 
    0.03099508, 0.02996059, 0.02850163, 0.02781407, 0.02766452, 0.02732809, 
    0.0263789, 0.02606515, 0.02665425, 0.02700929, 0.02659191, 0.02598628, 
    0.02622142, 0.02687633, 0.02725113, 0.02584471, 0.02667968, 0.02961284, 
    0.03578807, 0.03678761, 0.03049076, 0.02850749, 0.02822836, 0.02937653, 
    0.03102282, 0.03312102, 0.03401207, 0.03331856, 0.03104873, 0.02799021, 
    0.02441118, 0.02188916, 0.01963213, 0.01731311, 0.01388163, 0.01121303, 
    0.01145755, 0.01081989, 0.009366368, 0.009567187, 0.01059177, 0.01430051, 
    0.02158946, 0.04910821, 0.07323223, 0.06313359, 0.05699631, 0.06309833, 
    0.06945479, 0.07342558, 0.07947934, 0.08521953, 0.08902189, 0.08721576, 
    0.08040167, 0.07809604, 0.07348003, 0.07277366, 0.07154131, 0.0717627, 
    0.0730435, 0.0733472, 0.07315012, 0.07385633, 0.07572162, 0.07718313, 
    0.07937149, 0.08066833, 0.08201855, 0.08222319, 0.08204854, 0.08057863,
  0.07873114, 0.07672868, 0.07461166, 0.07237664, 0.07007594, 0.06769417, 
    0.06626792, 0.06507272, 0.06407732, 0.06365796, 0.06310718, 0.06252772, 
    0.06266493, 0.06536513, 0.06992372, 0.06761996, 0.05885042, 0.05261236, 
    0.05352956, 0.05415037, 0.05420695, 0.05583033, 0.05683599, 0.05728946, 
    0.05890498, 0.06019505, 0.06084538, 0.06060511, 0.05986686, 0.05891549, 
    0.05779193, 0.0568568, 0.05655031, 0.05635472, 0.05705487, 0.05815373, 
    0.05770369, 0.05652278, 0.05595837, 0.05551159, 0.05488726, 0.05353102, 
    0.05203341, 0.05139324, 0.05087355, 0.05022735, 0.04977517, 0.04907461, 
    0.04911305, 0.04846355, 0.04717395, 0.04887899, 0.04839175, 0.04398822, 
    0.04206485, 0.04211409, 0.04195174, 0.04070457, 0.03923687, 0.0387269, 
    0.03889868, 0.03905632, 0.03970861, 0.03994003, 0.03998163, 0.04005637, 
    0.04015533, 0.04033318, 0.04068866, 0.04079781, 0.04060031, 0.04002025, 
    0.03890444, 0.03716739, 0.0361176, 0.03528728, 0.03300394, 0.02980207, 
    0.02896176, 0.02941579, 0.02908968, 0.02844514, 0.02759291, 0.02756376, 
    0.02790538, 0.027624, 0.02684567, 0.02634742, 0.02632922, 0.02648536, 
    0.02682778, 0.02746032, 0.02766355, 0.02757827, 0.02738137, 0.02695206, 
    0.02621077, 0.02557562, 0.02561588, 0.0262224, 0.02816372, 0.02963969, 
    0.02751117, 0.02603594, 0.0280522, 0.02639355, 0.02350129, 0.02188088, 
    0.0221827, 0.02421699, 0.02544022, 0.02616247, 0.02703941, 0.02769399, 
    0.02576338, 0.02390386, 0.02334316, 0.0229534, 0.02177924, 0.02180761, 
    0.02203628, 0.02197285, 0.02214832, 0.02233516, 0.02252105, 0.02243051, 
    0.0224128, 0.0223194, 0.02232305, 0.02272257, 0.02334236, 0.02458903, 
    0.02677136, 0.02698965, 0.02511621, 0.02506905, 0.0264199, 0.02640045, 
    0.02480992, 0.02614863, 0.03116264, 0.03362343, 0.03412579, 0.03604475, 
    0.03808641, 0.03901889, 0.04073444, 0.04373121, 0.04452685, 0.04363913, 
    0.04391403, 0.0442642, 0.04406595, 0.04295344, 0.04121091, 0.03892479, 
    0.03698439, 0.03791415, 0.03850619, 0.03576517, 0.03734009, 0.03693707, 
    0.03478121, 0.03490009, 0.03575553, 0.0370979, 0.03410457, 0.03260975, 
    0.03735568, 0.03785444, 0.03627019, 0.0378451, 0.03836473, 0.036393, 
    0.03407591, 0.03097649, 0.02762468, 0.02785429, 0.02862238, 0.02768057, 
    0.02677861, 0.02550061, 0.02499428, 0.02552613, 0.0271173, 0.02806626, 
    0.02989082, 0.03075447, 0.03157552, 0.03288659, 0.03453517, 0.03628442, 
    0.03490613, 0.03351854, 0.03331061, 0.03099495, 0.02955083, 0.02876339, 
    0.02793001, 0.02721407, 0.02685157, 0.02683352, 0.02720258, 0.02731327, 
    0.02732125, 0.02741747, 0.02774389, 0.02782268, 0.02839163, 0.02862638, 
    0.02924299, 0.02947491, 0.02947125, 0.02938329, 0.02937513, 0.02899492, 
    0.02814756, 0.02708828, 0.02673028, 0.02705816, 0.02656298, 0.02542915, 
    0.02476166, 0.0245474, 0.02503898, 0.02549217, 0.0256796, 0.02569043, 
    0.02582492, 0.02662027, 0.02780735, 0.02868283, 0.03005808, 0.02981545, 
    0.03031554, 0.02923189, 0.02779323, 0.02673974, 0.02657877, 0.02733322, 
    0.02818532, 0.0296277, 0.0302605, 0.02982838, 0.02695538, 0.02315756, 
    0.02169999, 0.02076101, 0.01947187, 0.0175058, 0.01467937, 0.01129012, 
    0.009375268, 0.008023321, 0.006558553, 0.006050877, 0.006710421, 
    0.008259483, 0.01086476, 0.0147399, 0.01834062, 0.02235366, 0.03105876, 
    0.04011358, 0.04482698, 0.04620742, 0.05154724, 0.05747419, 0.06203266, 
    0.07309817, 0.07727819, 0.07942119, 0.07886332, 0.07669158, 0.07421526, 
    0.07404453, 0.07492635, 0.07521494, 0.07528429, 0.07582343, 0.07708799, 
    0.07810953, 0.07919502, 0.0800932, 0.08093521, 0.08118773, 0.08117595, 
    0.08008865,
  0.07768919, 0.07554206, 0.0737023, 0.07176733, 0.06999295, 0.06833351, 
    0.06668395, 0.06495223, 0.06320789, 0.06201337, 0.06040352, 0.05910799, 
    0.05861343, 0.05803754, 0.05890278, 0.06326994, 0.06571101, 0.06204385, 
    0.05723322, 0.05544841, 0.05434893, 0.05434602, 0.05464275, 0.05579132, 
    0.05705366, 0.05641558, 0.05528197, 0.05472291, 0.05580209, 0.05816532, 
    0.05866247, 0.05890012, 0.05985839, 0.06039279, 0.06013373, 0.05950841, 
    0.05874392, 0.05814527, 0.05738957, 0.05606829, 0.05461574, 0.05292803, 
    0.05167108, 0.0512886, 0.05055075, 0.04940281, 0.04832081, 0.04760833, 
    0.04837432, 0.04859166, 0.04625651, 0.04312668, 0.04266547, 0.04273549, 
    0.04156103, 0.04077167, 0.039999, 0.03837514, 0.03731224, 0.0370335, 
    0.03731035, 0.03736845, 0.03761739, 0.03770217, 0.03803758, 0.03809512, 
    0.03829624, 0.03850147, 0.0389515, 0.03947994, 0.03962248, 0.03946622, 
    0.03918635, 0.04022418, 0.03962657, 0.03541735, 0.03255858, 0.03107763, 
    0.03025746, 0.02968857, 0.02893635, 0.02851862, 0.02781157, 0.02798916, 
    0.02911262, 0.0310249, 0.03175189, 0.0300547, 0.02782516, 0.02715142, 
    0.02649185, 0.02595901, 0.02581332, 0.02583654, 0.02579243, 0.02557342, 
    0.02516803, 0.02489459, 0.02463938, 0.02435884, 0.02533076, 0.02786485, 
    0.02579253, 0.0246864, 0.02695077, 0.02674785, 0.02533631, 0.02429943, 
    0.02409448, 0.0244565, 0.02398274, 0.02339467, 0.02413672, 0.02457207, 
    0.02395379, 0.0229615, 0.02224562, 0.02177445, 0.02124358, 0.02090095, 
    0.02086456, 0.02095672, 0.02099901, 0.02118484, 0.02139076, 0.02162287, 
    0.02183623, 0.02215732, 0.02260116, 0.02353919, 0.02447397, 0.02563369, 
    0.02655403, 0.02629391, 0.02466409, 0.02429927, 0.02370453, 0.02405192, 
    0.02548897, 0.02668775, 0.02725594, 0.02850596, 0.03076424, 0.03349753, 
    0.03501784, 0.03696248, 0.03875736, 0.03978417, 0.04053137, 0.04141973, 
    0.04201964, 0.04271904, 0.0434599, 0.04287471, 0.04071439, 0.03854943, 
    0.03690622, 0.03435127, 0.03269254, 0.03236729, 0.03282562, 0.03145489, 
    0.03022536, 0.03178171, 0.03359599, 0.03435627, 0.03364596, 0.03172676, 
    0.03205172, 0.03065893, 0.02882762, 0.02904134, 0.02945499, 0.03054245, 
    0.03158356, 0.03155157, 0.0289182, 0.0268324, 0.02528455, 0.02428974, 
    0.02396807, 0.02405898, 0.02410095, 0.02471066, 0.02649096, 0.02868468, 
    0.03008812, 0.02981091, 0.02975967, 0.03167387, 0.03463423, 0.035418, 
    0.03257479, 0.03089223, 0.03131111, 0.03189364, 0.03062163, 0.02847177, 
    0.02812526, 0.02888196, 0.02883126, 0.02858212, 0.02843282, 0.02850473, 
    0.02842148, 0.02804871, 0.02759782, 0.0271977, 0.02621585, 0.02623853, 
    0.02641133, 0.02655361, 0.02653029, 0.02609668, 0.02589104, 0.02577394, 
    0.02508505, 0.02383278, 0.02352828, 0.02443551, 0.02469974, 0.02402055, 
    0.02331734, 0.02346846, 0.02380019, 0.02392782, 0.02430208, 0.02506841, 
    0.0261967, 0.02733576, 0.02825361, 0.03122513, 0.03338202, 0.03035862, 
    0.02656237, 0.026208, 0.02554003, 0.02490136, 0.02435707, 0.02481622, 
    0.02624217, 0.02731048, 0.02772763, 0.02619075, 0.02512277, 0.02416274, 
    0.02039198, 0.01713113, 0.0170642, 0.01636393, 0.01453459, 0.01156246, 
    0.008967145, 0.007414438, 0.005938448, 0.005098359, 0.005544522, 
    0.006266736, 0.00678795, 0.006614801, 0.007778181, 0.009145586, 
    0.01368443, 0.01886699, 0.02372731, 0.03044033, 0.04531545, 0.06182382, 
    0.06416893, 0.05845626, 0.0640235, 0.07332256, 0.07705264, 0.07622689, 
    0.07574272, 0.07662349, 0.07754695, 0.07785132, 0.07710268, 0.0774627, 
    0.07785557, 0.07838996, 0.0787987, 0.0792411, 0.08017164, 0.08058896, 
    0.08025787, 0.07901227,
  0.07532079, 0.07382081, 0.07233258, 0.07102875, 0.07001527, 0.06873608, 
    0.06712169, 0.06555105, 0.06412903, 0.0629675, 0.0618379, 0.06068347, 
    0.05949382, 0.05813692, 0.05577151, 0.05483348, 0.05518692, 0.0560238, 
    0.05517038, 0.05488824, 0.05838092, 0.05883541, 0.05560172, 0.05504824, 
    0.05540246, 0.05509807, 0.05573762, 0.0584477, 0.06048043, 0.06126414, 
    0.06174668, 0.06207805, 0.06249248, 0.06243891, 0.06170559, 0.06145976, 
    0.06152978, 0.06125708, 0.06018861, 0.05830569, 0.05610401, 0.05380544, 
    0.05204227, 0.05076406, 0.04877821, 0.04686442, 0.04586866, 0.04546357, 
    0.04483923, 0.04444857, 0.04394983, 0.04301258, 0.04175475, 0.04092558, 
    0.04013955, 0.03928045, 0.03842145, 0.03730923, 0.03674746, 0.03663461, 
    0.03662207, 0.0363897, 0.03606433, 0.03591034, 0.03561623, 0.0354424, 
    0.0352358, 0.03527007, 0.03574803, 0.03648287, 0.03632266, 0.03562952, 
    0.03492743, 0.03455549, 0.03320169, 0.03174165, 0.03156535, 0.03060937, 
    0.03007757, 0.02965453, 0.02910342, 0.02849957, 0.02880783, 0.03003605, 
    0.03151736, 0.03263177, 0.03313217, 0.03156812, 0.02992231, 0.02867645, 
    0.02699676, 0.02547965, 0.02495405, 0.02460429, 0.02460892, 0.02462261, 
    0.02451968, 0.02461322, 0.02480833, 0.02484659, 0.02588782, 0.02750434, 
    0.0268202, 0.02582232, 0.02619378, 0.02618632, 0.02551821, 0.02464281, 
    0.02314764, 0.02320427, 0.02340532, 0.02293769, 0.02279694, 0.02278701, 
    0.02235705, 0.02200178, 0.02184573, 0.02174807, 0.02176534, 0.02189826, 
    0.02206661, 0.02220291, 0.02207203, 0.02204465, 0.02213241, 0.02241139, 
    0.02300596, 0.02367938, 0.02418039, 0.02504881, 0.02521673, 0.02488068, 
    0.02444912, 0.02399456, 0.02344429, 0.02316098, 0.02351902, 0.0238319, 
    0.02394908, 0.02459658, 0.02526057, 0.02611285, 0.02737298, 0.02955504, 
    0.0312744, 0.03282308, 0.03396519, 0.03549844, 0.03785863, 0.03901367, 
    0.04001971, 0.04053262, 0.04083597, 0.04023276, 0.03919508, 0.0382815, 
    0.03708502, 0.03495918, 0.03211592, 0.03092235, 0.03011182, 0.02926932, 
    0.02844947, 0.02810078, 0.02725387, 0.02686895, 0.02782505, 0.02716692, 
    0.02576183, 0.02520981, 0.02537185, 0.0264732, 0.02700306, 0.0266965, 
    0.02758083, 0.02800351, 0.02710811, 0.02540872, 0.02441249, 0.0238331, 
    0.0235452, 0.02389656, 0.02457597, 0.02610927, 0.02725893, 0.02769595, 
    0.0281842, 0.02897275, 0.02968618, 0.03022568, 0.03033661, 0.02901181, 
    0.02870229, 0.02909661, 0.02993291, 0.03002668, 0.02829501, 0.02810514, 
    0.02928428, 0.03057715, 0.03079383, 0.03068089, 0.03027897, 0.0300836, 
    0.02957916, 0.02856343, 0.02711849, 0.0263773, 0.02507382, 0.02513172, 
    0.02652802, 0.02736506, 0.02691344, 0.02533015, 0.02482907, 0.02399908, 
    0.02349229, 0.02297611, 0.02297671, 0.02333686, 0.02434851, 0.02461073, 
    0.02430632, 0.02382429, 0.02361149, 0.02310613, 0.02362913, 0.02598175, 
    0.02788982, 0.02828196, 0.02734189, 0.02652535, 0.02561034, 0.02431893, 
    0.02412746, 0.0243885, 0.02335976, 0.02318701, 0.02342547, 0.02544079, 
    0.02750099, 0.02795658, 0.02746206, 0.02660611, 0.0255562, 0.02351936, 
    0.01910261, 0.01529045, 0.01516617, 0.01580991, 0.01443174, 0.01229022, 
    0.009127212, 0.007467016, 0.006486935, 0.00598706, 0.005758731, 
    0.005566111, 0.004824356, 0.004562692, 0.00517362, 0.006137937, 
    0.006853093, 0.007517867, 0.01007144, 0.01374787, 0.0180661, 0.02378243, 
    0.0331375, 0.04029418, 0.05007716, 0.05974958, 0.06515863, 0.06743486, 
    0.07038803, 0.0739492, 0.07616682, 0.0770917, 0.07665848, 0.07721134, 
    0.07795975, 0.07822353, 0.07792936, 0.07770623, 0.07797809, 0.07820761, 
    0.07776581, 0.07659764,
  0.07321498, 0.07231235, 0.07106166, 0.07017588, 0.0697015, 0.06931753, 
    0.06828535, 0.06680828, 0.06552214, 0.06437367, 0.06282438, 0.06152888, 
    0.06082416, 0.06007583, 0.05899305, 0.05742379, 0.05810114, 0.05799884, 
    0.05606181, 0.05582031, 0.05700281, 0.05638947, 0.05535655, 0.05702337, 
    0.05938769, 0.06031386, 0.06111062, 0.06223692, 0.06301501, 0.06341934, 
    0.06370621, 0.06381591, 0.06363056, 0.06349549, 0.06350258, 0.06360988, 
    0.06347319, 0.06317495, 0.06194834, 0.05995687, 0.05656002, 0.05377707, 
    0.05218172, 0.05013973, 0.04704945, 0.04506429, 0.04387571, 0.04289512, 
    0.04241841, 0.04250549, 0.04197424, 0.04146837, 0.04080922, 0.0400121, 
    0.03894648, 0.03821737, 0.03734285, 0.03675804, 0.03638293, 0.03641893, 
    0.0362442, 0.03581608, 0.03538685, 0.0351792, 0.0348609, 0.03444463, 
    0.03365564, 0.03279203, 0.03230618, 0.03279662, 0.03253339, 0.03201514, 
    0.03153999, 0.03102978, 0.03081327, 0.03035807, 0.02950971, 0.02838353, 
    0.02767571, 0.0272013, 0.02682164, 0.02670045, 0.02783166, 0.02871037, 
    0.02994816, 0.03104508, 0.03106167, 0.03074255, 0.03137869, 0.03057442, 
    0.02767491, 0.02624477, 0.02581416, 0.02527674, 0.02476829, 0.02482498, 
    0.02507692, 0.02537015, 0.02569882, 0.02597951, 0.02662434, 0.02720487, 
    0.02664232, 0.02511539, 0.02434206, 0.02367312, 0.02312106, 0.02236184, 
    0.02169015, 0.02145859, 0.02154061, 0.02154372, 0.02166753, 0.02174613, 
    0.02173684, 0.02185179, 0.02202329, 0.02228274, 0.02273957, 0.02324812, 
    0.02388684, 0.02471257, 0.02490663, 0.02498656, 0.02505026, 0.02507438, 
    0.02535148, 0.02548999, 0.02539687, 0.02531586, 0.02522675, 0.02436613, 
    0.02398944, 0.02343522, 0.02295379, 0.02278671, 0.02239344, 0.0227198, 
    0.0236264, 0.0245764, 0.02503745, 0.02487742, 0.02560033, 0.02638676, 
    0.02733773, 0.0284135, 0.03085878, 0.03243892, 0.03398112, 0.03512834, 
    0.03592054, 0.03665483, 0.03688686, 0.03675419, 0.03590118, 0.03516051, 
    0.034644, 0.03411798, 0.03312331, 0.0318897, 0.03095377, 0.03002732, 
    0.02846464, 0.02785728, 0.02775203, 0.02730319, 0.02653007, 0.0264612, 
    0.02603526, 0.02586664, 0.02573031, 0.02600085, 0.02620409, 0.02614226, 
    0.0259436, 0.02555865, 0.0244954, 0.02396803, 0.0244603, 0.02492319, 
    0.02493287, 0.02533483, 0.02639032, 0.02690493, 0.0272432, 0.0267404, 
    0.02651701, 0.02649103, 0.02683182, 0.02721827, 0.02702665, 0.02656852, 
    0.02630297, 0.02737177, 0.02825152, 0.03055356, 0.03194531, 0.03226659, 
    0.0330571, 0.03298099, 0.03197491, 0.03083082, 0.03017515, 0.02887676, 
    0.0280604, 0.02690003, 0.02587569, 0.02527296, 0.0247226, 0.02489418, 
    0.02604853, 0.0267165, 0.02640067, 0.0249141, 0.02440484, 0.02412853, 
    0.02427949, 0.02409364, 0.02336787, 0.02334593, 0.02415909, 0.02531108, 
    0.02544841, 0.02486683, 0.02494738, 0.02518779, 0.02776507, 0.02900337, 
    0.02838044, 0.02691935, 0.02595807, 0.02441302, 0.02449745, 0.02422944, 
    0.02406776, 0.0237199, 0.02340946, 0.02337769, 0.02402013, 0.02494124, 
    0.02616634, 0.02618774, 0.02496065, 0.02256017, 0.01916056, 0.0161104, 
    0.01603108, 0.01766545, 0.01772529, 0.01565126, 0.01270081, 0.009761089, 
    0.007999327, 0.007062942, 0.006438474, 0.005974101, 0.005889356, 
    0.00552346, 0.00510462, 0.004328318, 0.004031623, 0.004408936, 
    0.004970905, 0.006231547, 0.007942936, 0.01102824, 0.015247, 0.02050471, 
    0.02668369, 0.03238354, 0.03971014, 0.0465562, 0.05312081, 0.05837479, 
    0.06310268, 0.06843967, 0.07169368, 0.07409635, 0.07501157, 0.07613444, 
    0.07650819, 0.07666469, 0.07632632, 0.07585414, 0.07573035, 0.07555694, 
    0.07505252, 0.07427611,
  0.0716515, 0.07114205, 0.07072167, 0.07057973, 0.07026485, 0.0697326, 
    0.06916229, 0.0686037, 0.06782378, 0.06703173, 0.06625294, 0.06527971, 
    0.06437442, 0.06321036, 0.06172949, 0.06077273, 0.06042036, 0.06070016, 
    0.06117566, 0.06148342, 0.06209234, 0.06323446, 0.06407146, 0.06453139, 
    0.06490777, 0.06501992, 0.0649533, 0.0648941, 0.06459203, 0.06419096, 
    0.06394003, 0.06378628, 0.06345497, 0.06319887, 0.06326984, 0.06365986, 
    0.06424341, 0.06391578, 0.06257138, 0.05999684, 0.05740041, 0.05512261, 
    0.05764661, 0.05804508, 0.05332979, 0.04414141, 0.04165712, 0.04113063, 
    0.04139572, 0.04045692, 0.03941821, 0.03810478, 0.03760882, 0.03827464, 
    0.03816478, 0.03754553, 0.03614831, 0.03593131, 0.03618224, 0.03690046, 
    0.03678609, 0.03608803, 0.03570805, 0.0356339, 0.03741486, 0.03691045, 
    0.03549926, 0.03321507, 0.03245912, 0.03202721, 0.03136527, 0.03069661, 
    0.0293358, 0.02845589, 0.02774722, 0.02722095, 0.02655129, 0.02595406, 
    0.02542104, 0.0250682, 0.0249687, 0.0253529, 0.02587297, 0.02656859, 
    0.02702351, 0.02762955, 0.02821356, 0.02857487, 0.0289049, 0.02796262, 
    0.02722455, 0.02696254, 0.02682922, 0.02623923, 0.02592008, 0.0257476, 
    0.02571783, 0.02567172, 0.02579743, 0.02600529, 0.02594901, 0.02560663, 
    0.02529556, 0.0252144, 0.02511409, 0.02485706, 0.02425002, 0.02350938, 
    0.02312056, 0.02271377, 0.02228501, 0.02194047, 0.02189642, 0.02193935, 
    0.02208427, 0.02233772, 0.02278459, 0.023486, 0.02398021, 0.02452121, 
    0.0254391, 0.0257862, 0.02566946, 0.02516502, 0.02524677, 0.02560522, 
    0.02578747, 0.0258834, 0.02554784, 0.02525041, 0.02491697, 0.02438462, 
    0.02411388, 0.02404262, 0.02410616, 0.02408024, 0.02439978, 0.02466997, 
    0.02490556, 0.02520878, 0.02558434, 0.02567445, 0.0261748, 0.02667916, 
    0.02729371, 0.02826278, 0.02921245, 0.02969336, 0.03050659, 0.03118634, 
    0.03180361, 0.03252169, 0.03335154, 0.03354247, 0.03358857, 0.03359148, 
    0.03343683, 0.03313394, 0.03278888, 0.03223304, 0.03164789, 0.0308545, 
    0.03025319, 0.02973441, 0.02941871, 0.02899722, 0.02865238, 0.02835715, 
    0.02818183, 0.02800854, 0.02767906, 0.02712104, 0.02695845, 0.02712285, 
    0.02676598, 0.02608365, 0.02604715, 0.02639735, 0.02629085, 0.02601592, 
    0.02580052, 0.02587141, 0.02610608, 0.0265776, 0.02668392, 0.02662529, 
    0.02563712, 0.02534956, 0.02614839, 0.02804467, 0.02822759, 0.02795706, 
    0.02695742, 0.02692086, 0.02771896, 0.0294071, 0.03002028, 0.03047071, 
    0.03067435, 0.03074735, 0.03005661, 0.02944076, 0.02888677, 0.02799915, 
    0.02734267, 0.02618691, 0.02559994, 0.02533597, 0.02643732, 0.02659426, 
    0.02659332, 0.02632346, 0.02614408, 0.02529771, 0.0248842, 0.02502706, 
    0.0267412, 0.0268635, 0.02591123, 0.02376986, 0.02388046, 0.02511271, 
    0.02662981, 0.02745312, 0.02745163, 0.02701587, 0.02695171, 0.02457293, 
    0.0230551, 0.02280791, 0.02302415, 0.02324978, 0.02355501, 0.02301681, 
    0.02254128, 0.02224328, 0.02232282, 0.02305818, 0.02348554, 0.02429155, 
    0.02387987, 0.0218843, 0.01985661, 0.01811943, 0.01688941, 0.01625716, 
    0.01673881, 0.01715123, 0.01526397, 0.01209552, 0.009996142, 0.008188894, 
    0.007274842, 0.006708029, 0.00621935, 0.006078088, 0.005834338, 
    0.005442473, 0.004797427, 0.004465941, 0.004225201, 0.004166346, 
    0.004476589, 0.005008305, 0.00550219, 0.007538688, 0.01015518, 
    0.01437498, 0.0190718, 0.02538258, 0.03155753, 0.0373242, 0.04429582, 
    0.05023464, 0.0562041, 0.06182294, 0.0661669, 0.07012841, 0.07231586, 
    0.07420425, 0.07324021, 0.0735345, 0.07384813, 0.07380714, 0.07363079, 
    0.07335463, 0.07290087, 0.07243475,
  0.06995843, 0.06971903, 0.06954571, 0.06997277, 0.07023616, 0.07007417, 
    0.06982622, 0.06946035, 0.06903684, 0.06882011, 0.06846148, 0.06780808, 
    0.06667479, 0.06557599, 0.06456295, 0.06338915, 0.06286516, 0.0631145, 
    0.06376053, 0.06488501, 0.06579453, 0.06670932, 0.067418, 0.06758419, 
    0.06771711, 0.06770959, 0.06733772, 0.06670057, 0.06591909, 0.06479404, 
    0.06351959, 0.06242353, 0.06184577, 0.06174333, 0.06204331, 0.0622499, 
    0.06266511, 0.06300687, 0.06209459, 0.0604929, 0.05778232, 0.05427063, 
    0.05221109, 0.05448817, 0.05570566, 0.05186343, 0.04425945, 0.04094512, 
    0.03989077, 0.03907079, 0.03861762, 0.03824374, 0.03738391, 0.03693515, 
    0.03667821, 0.03614437, 0.0355373, 0.03541291, 0.03624534, 0.03688378, 
    0.0369001, 0.03627821, 0.03602277, 0.03595395, 0.03760932, 0.03697685, 
    0.03586545, 0.03310149, 0.03224058, 0.03162207, 0.03189063, 0.03137121, 
    0.02969624, 0.02775085, 0.02690645, 0.02732633, 0.02763126, 0.02703842, 
    0.02595033, 0.02597862, 0.02603989, 0.02618942, 0.02621274, 0.02631832, 
    0.02650009, 0.02640741, 0.02612824, 0.02605934, 0.02701043, 0.02706303, 
    0.02710922, 0.02723499, 0.0269794, 0.02665246, 0.02629592, 0.0260545, 
    0.02597923, 0.02610774, 0.02571991, 0.02496145, 0.02500696, 0.02573284, 
    0.0265083, 0.02696012, 0.02681152, 0.02601358, 0.02523287, 0.024764, 
    0.02434635, 0.02408105, 0.02369528, 0.02320039, 0.02279741, 0.02292452, 
    0.02322088, 0.02404527, 0.02505039, 0.02532251, 0.02548372, 0.02563658, 
    0.0256919, 0.02558042, 0.02518543, 0.02502054, 0.02490012, 0.02494505, 
    0.02502435, 0.0252688, 0.0254614, 0.02545662, 0.02532086, 0.0251864, 
    0.02509789, 0.02497759, 0.02502603, 0.0250948, 0.0253287, 0.0255507, 
    0.02579163, 0.02608731, 0.02633488, 0.02662324, 0.02691586, 0.02717742, 
    0.02734016, 0.02757417, 0.02790286, 0.02824757, 0.02881138, 0.02931834, 
    0.02999287, 0.03053636, 0.03097985, 0.03129262, 0.03144456, 0.03156294, 
    0.03158088, 0.03149864, 0.03132695, 0.03122736, 0.03105297, 0.03075176, 
    0.03038586, 0.03002739, 0.02970902, 0.0294616, 0.02921621, 0.02893725, 
    0.02864235, 0.02840935, 0.02812074, 0.02779524, 0.0275897, 0.02752963, 
    0.02732197, 0.02696303, 0.02674676, 0.0266101, 0.02634119, 0.02605795, 
    0.02582797, 0.02547947, 0.02542585, 0.02549438, 0.02556108, 0.02559538, 
    0.0258468, 0.02591234, 0.02649277, 0.02742237, 0.02878091, 0.02920609, 
    0.02920336, 0.0288418, 0.02906226, 0.02901587, 0.02773065, 0.02603296, 
    0.02588897, 0.02599956, 0.0262332, 0.02622184, 0.02659456, 0.02669973, 
    0.02651389, 0.02611022, 0.02600607, 0.02600229, 0.02701527, 0.02710623, 
    0.02717807, 0.02672178, 0.02639175, 0.02565377, 0.02505727, 0.02510011, 
    0.02608714, 0.02661652, 0.02626046, 0.02565621, 0.02565602, 0.02534589, 
    0.02722478, 0.02748403, 0.02631264, 0.02438251, 0.02375854, 0.02258071, 
    0.02198613, 0.02190516, 0.02126441, 0.02120463, 0.02153905, 0.02137556, 
    0.0210371, 0.02104384, 0.02147021, 0.02206657, 0.02378896, 0.0251573, 
    0.02395374, 0.02041001, 0.01746817, 0.01602948, 0.01479469, 0.01429639, 
    0.01351729, 0.01205294, 0.01052873, 0.008801954, 0.007283441, 
    0.006454876, 0.005991087, 0.005697061, 0.005441713, 0.005072094, 
    0.004502845, 0.004109027, 0.00395073, 0.003677051, 0.003529439, 
    0.003755657, 0.003998119, 0.004400206, 0.005577939, 0.006755748, 
    0.008617328, 0.01137299, 0.01389324, 0.01775103, 0.02232414, 0.02738857, 
    0.03356162, 0.03956424, 0.04755144, 0.05414337, 0.05954709, 0.06484763, 
    0.06806769, 0.0710214, 0.07111079, 0.07185957, 0.07238013, 0.07123333, 
    0.07107074, 0.07087259, 0.07055632, 0.07025856,
  0.06860585, 0.0679152, 0.06767669, 0.06760912, 0.0680648, 0.0682332, 
    0.06835718, 0.0686151, 0.0687924, 0.06872766, 0.06902124, 0.06895952, 
    0.06839614, 0.0673642, 0.06596942, 0.06522409, 0.06497288, 0.06534933, 
    0.06646522, 0.06745658, 0.06809426, 0.06893092, 0.06951698, 0.06995811, 
    0.0696229, 0.06881596, 0.06785072, 0.06696228, 0.06561156, 0.06417858, 
    0.06282271, 0.06197508, 0.06136118, 0.06084052, 0.06090802, 0.06105288, 
    0.06093502, 0.06063446, 0.06026086, 0.05872482, 0.05701832, 0.05472481, 
    0.04963505, 0.04878585, 0.05057, 0.05969097, 0.05441413, 0.04934599, 
    0.04242193, 0.03873405, 0.03567766, 0.0342678, 0.03650482, 0.03598983, 
    0.03559697, 0.03618647, 0.03594671, 0.03570315, 0.03570046, 0.03563562, 
    0.03554761, 0.03530339, 0.03510294, 0.03490796, 0.03439229, 0.03388243, 
    0.03332987, 0.03171022, 0.03144216, 0.03137548, 0.03352065, 0.03338575, 
    0.03307549, 0.0322211, 0.03184291, 0.03135757, 0.02795969, 0.02656442, 
    0.02636201, 0.02746601, 0.02687748, 0.02654685, 0.02621358, 0.0269463, 
    0.02720447, 0.02668254, 0.02567985, 0.02675913, 0.02818105, 0.02882439, 
    0.02700737, 0.02659855, 0.026433, 0.02639678, 0.02644876, 0.02650891, 
    0.02668386, 0.02683403, 0.02693472, 0.0268591, 0.02689664, 0.02699601, 
    0.02691695, 0.02659495, 0.02609085, 0.02557739, 0.02488226, 0.0240929, 
    0.02350729, 0.02321108, 0.02298912, 0.02265106, 0.02276352, 0.02312436, 
    0.02402099, 0.02470217, 0.02510645, 0.02485054, 0.02492519, 0.02527567, 
    0.02567634, 0.02559711, 0.0254907, 0.025202, 0.02448165, 0.02442461, 
    0.02445076, 0.02484203, 0.02500097, 0.02514615, 0.02532849, 0.02533088, 
    0.02531772, 0.02511624, 0.02518584, 0.02525788, 0.02561892, 0.02581329, 
    0.02600533, 0.02626335, 0.02644554, 0.02660513, 0.02656939, 0.02672388, 
    0.02686163, 0.02701602, 0.02729995, 0.02756663, 0.02777386, 0.02804107, 
    0.02835126, 0.02875283, 0.02901522, 0.02924801, 0.0294526, 0.02977613, 
    0.02990433, 0.02991262, 0.0297745, 0.0297386, 0.02975706, 0.02979157, 
    0.02960207, 0.02942497, 0.02927241, 0.0291239, 0.02883588, 0.02856097, 
    0.02821341, 0.02789077, 0.02764175, 0.02746816, 0.02731748, 0.02713767, 
    0.02695164, 0.02674195, 0.02659124, 0.02646847, 0.0264651, 0.02646467, 
    0.02634759, 0.02600281, 0.02543504, 0.02501723, 0.02482243, 0.0247076, 
    0.02483181, 0.02509283, 0.02534917, 0.02575554, 0.02690014, 0.02732264, 
    0.02709609, 0.0251817, 0.02493822, 0.02511739, 0.02526407, 0.02486522, 
    0.02451025, 0.02433394, 0.02420167, 0.0241403, 0.02493142, 0.02491825, 
    0.02482454, 0.02433514, 0.02444223, 0.02453986, 0.02543429, 0.02550861, 
    0.02555325, 0.0250467, 0.02502095, 0.02500268, 0.02581846, 0.02613081, 
    0.02641031, 0.02610648, 0.02616096, 0.02630528, 0.02261735, 0.02192587, 
    0.02370172, 0.02507663, 0.0216291, 0.02030361, 0.01976717, 0.02079959, 
    0.02075086, 0.02016018, 0.01903439, 0.0192485, 0.01989795, 0.02104243, 
    0.02184767, 0.02230509, 0.0221509, 0.0217892, 0.022538, 0.02243686, 
    0.02067275, 0.01811668, 0.01694342, 0.01640356, 0.01562476, 0.01417996, 
    0.0124939, 0.01113252, 0.009438115, 0.007765074, 0.006206553, 
    0.005957027, 0.005807415, 0.00525811, 0.004780693, 0.004063783, 
    0.003461306, 0.002975318, 0.002939825, 0.002949929, 0.002926055, 
    0.002936252, 0.00302452, 0.003513828, 0.003914488, 0.00475063, 
    0.006280338, 0.007806127, 0.009636582, 0.01237219, 0.01511784, 
    0.01784706, 0.02280116, 0.02811974, 0.03725653, 0.0431083, 0.04881833, 
    0.05541631, 0.05955453, 0.06362621, 0.06756366, 0.06922874, 0.07085758, 
    0.06865379, 0.0686811, 0.06886096, 0.06871319, 0.06863483,
  0.06906155, 0.06905086, 0.06778993, 0.06792921, 0.06816265, 0.06878117, 
    0.06910409, 0.06937351, 0.06972189, 0.06944497, 0.06902441, 0.06857014, 
    0.06838539, 0.06760088, 0.06641274, 0.06416091, 0.06294224, 0.06283221, 
    0.0631353, 0.0645586, 0.06627919, 0.06697454, 0.0672665, 0.0674204, 
    0.06687175, 0.06614332, 0.06523693, 0.06395661, 0.06224014, 0.06032036, 
    0.05936491, 0.05901978, 0.05935646, 0.05965585, 0.05969779, 0.05942998, 
    0.05865393, 0.05792413, 0.05710139, 0.05594477, 0.05419512, 0.05287353, 
    0.05189728, 0.04953757, 0.05060234, 0.05654273, 0.0584041, 0.05704285, 
    0.04971304, 0.04786418, 0.04500623, 0.03921092, 0.03762286, 0.03647476, 
    0.03532252, 0.03498979, 0.03467847, 0.03487593, 0.03481441, 0.03451808, 
    0.034206, 0.03380798, 0.03349958, 0.03319376, 0.03348376, 0.03312125, 
    0.03276103, 0.03243785, 0.03226949, 0.03206782, 0.03223987, 0.03202584, 
    0.03167276, 0.03162428, 0.03221103, 0.03150687, 0.03076635, 0.03071606, 
    0.03001334, 0.02897911, 0.0265644, 0.02656667, 0.02699287, 0.02790735, 
    0.02919536, 0.02981171, 0.03007143, 0.03061955, 0.03024368, 0.02871665, 
    0.02680931, 0.02561735, 0.02587348, 0.02586571, 0.02600816, 0.02637961, 
    0.02615706, 0.02604487, 0.02621678, 0.02667904, 0.02686583, 0.02667502, 
    0.02644554, 0.02624159, 0.0258648, 0.02515222, 0.02442869, 0.02380515, 
    0.02320628, 0.02261026, 0.02226955, 0.02210234, 0.02199776, 0.02192179, 
    0.02223871, 0.02292555, 0.02356791, 0.02354748, 0.02372797, 0.02430849, 
    0.02510223, 0.02517246, 0.02509832, 0.02439606, 0.02424094, 0.02418122, 
    0.02447434, 0.02472221, 0.02487859, 0.02513312, 0.02538963, 0.02547397, 
    0.02549038, 0.02529731, 0.02536462, 0.02543187, 0.02572295, 0.02586068, 
    0.02599671, 0.02621225, 0.02630375, 0.02637247, 0.02633025, 0.02632991, 
    0.02640205, 0.02647437, 0.02656366, 0.02666533, 0.0267504, 0.02683249, 
    0.02695211, 0.02708202, 0.02717488, 0.0274182, 0.02765569, 0.02795221, 
    0.02825606, 0.02839766, 0.02850961, 0.02859934, 0.02859268, 0.02851046, 
    0.0284206, 0.02837529, 0.02831149, 0.02812171, 0.02787323, 0.0275677, 
    0.02719239, 0.02689797, 0.02667989, 0.02655853, 0.02639343, 0.0261851, 
    0.02607602, 0.02600028, 0.026008, 0.02617115, 0.02627809, 0.02627046, 
    0.02617423, 0.02590658, 0.02557145, 0.02525766, 0.02489455, 0.02467175, 
    0.02455931, 0.02449275, 0.02450888, 0.02453307, 0.02459612, 0.02483084, 
    0.02486059, 0.02511474, 0.02623406, 0.03023517, 0.03015434, 0.02956975, 
    0.02620683, 0.0251792, 0.02479104, 0.02506609, 0.02560471, 0.02556583, 
    0.02535087, 0.0245111, 0.02458004, 0.02464797, 0.02594036, 0.02599082, 
    0.02603985, 0.02524315, 0.02487746, 0.02485324, 0.02549416, 0.02598452, 
    0.0259098, 0.02524095, 0.02294581, 0.02340407, 0.02530049, 0.0399317, 
    0.04140109, 0.03904266, 0.02728312, 0.02151632, 0.02023672, 0.01984457, 
    0.02056283, 0.02083076, 0.02077018, 0.02050735, 0.02063506, 0.02091173, 
    0.02119783, 0.02145026, 0.02114641, 0.02053298, 0.0197803, 0.01904102, 
    0.01817104, 0.01705482, 0.01626826, 0.01603821, 0.01462446, 0.01207999, 
    0.01044199, 0.009481807, 0.008856134, 0.007322167, 0.006057046, 
    0.00525279, 0.005118116, 0.005049787, 0.004552295, 0.004055561, 
    0.003395126, 0.002861722, 0.002695991, 0.002723149, 0.003067741, 
    0.003220465, 0.003417081, 0.003443871, 0.003685042, 0.004577696, 
    0.005623404, 0.007433737, 0.009283212, 0.01118699, 0.01243959, 
    0.01523424, 0.01884098, 0.0236217, 0.02934659, 0.03391828, 0.03847452, 
    0.04317874, 0.04757936, 0.05198327, 0.06054934, 0.06333452, 0.06614561, 
    0.06599283, 0.06629453, 0.06729189, 0.068198, 0.06861148,
  0.06882598, 0.06985036, 0.07051083, 0.07112386, 0.07142413, 0.07176729, 
    0.07184929, 0.07120672, 0.07040163, 0.06899095, 0.06877276, 0.06847911, 
    0.06757903, 0.06460532, 0.05874953, 0.05660474, 0.05569747, 0.05641018, 
    0.05688203, 0.05698099, 0.05733994, 0.05835455, 0.05932573, 0.05970312, 
    0.05943254, 0.05897551, 0.05829562, 0.05778976, 0.05719838, 0.05665848, 
    0.05620642, 0.05601691, 0.05577558, 0.05566112, 0.05555588, 0.05524463, 
    0.05457676, 0.05361711, 0.05229278, 0.05111519, 0.05008731, 0.04926247, 
    0.04937037, 0.04698649, 0.04524105, 0.04366818, 0.04272166, 0.04161859, 
    0.03989152, 0.03926619, 0.04122804, 0.04046742, 0.03942104, 0.03881732, 
    0.037892, 0.03702758, 0.03607796, 0.03494533, 0.03456369, 0.03407518, 
    0.03359029, 0.03307641, 0.03264979, 0.03222634, 0.03164573, 0.03134445, 
    0.03104048, 0.0309989, 0.03099278, 0.030763, 0.0304634, 0.02997745, 
    0.02970167, 0.02939898, 0.02905082, 0.0278537, 0.02711466, 0.02629759, 
    0.02519517, 0.02487958, 0.02477598, 0.02563985, 0.0274914, 0.02784764, 
    0.02793775, 0.02787535, 0.02671755, 0.02618263, 0.02595566, 0.02537079, 
    0.02508019, 0.02523289, 0.02560559, 0.02599081, 0.02621368, 0.02635677, 
    0.02642361, 0.02639764, 0.02667468, 0.02684776, 0.02702997, 0.02712127, 
    0.02701193, 0.02670459, 0.02621626, 0.02557106, 0.02500891, 0.02441639, 
    0.02393628, 0.02356515, 0.02340942, 0.02337448, 0.02334602, 0.02337006, 
    0.02363008, 0.02403815, 0.02413991, 0.02423525, 0.0244665, 0.02468429, 
    0.02473371, 0.02469207, 0.02437409, 0.02427253, 0.02420623, 0.02420394, 
    0.02439966, 0.02454147, 0.02469581, 0.02498435, 0.02512201, 0.02524301, 
    0.02533116, 0.02536448, 0.02543043, 0.02549639, 0.02560828, 0.02566217, 
    0.02571471, 0.02567494, 0.02561215, 0.02561927, 0.02561187, 0.02561389, 
    0.02565558, 0.02569153, 0.02578519, 0.02594505, 0.02600771, 0.0260297, 
    0.025804, 0.02581672, 0.02591908, 0.0261005, 0.02630051, 0.02645301, 
    0.02659717, 0.02684402, 0.0271444, 0.02725339, 0.02730256, 0.02721789, 
    0.0272064, 0.02716805, 0.02705535, 0.02685971, 0.02656531, 0.02620257, 
    0.02587715, 0.02555849, 0.02542251, 0.02536, 0.02526684, 0.02512138, 
    0.0250079, 0.02494641, 0.0249252, 0.02489402, 0.0248666, 0.02491378, 
    0.02501648, 0.02510058, 0.02508252, 0.02489679, 0.02478112, 0.02462011, 
    0.02433841, 0.02421473, 0.02423466, 0.02431131, 0.0245937, 0.02491335, 
    0.02521273, 0.02534077, 0.02516544, 0.02552866, 0.02588125, 0.02553756, 
    0.02400223, 0.02371067, 0.02345643, 0.02425906, 0.02445094, 0.0245203, 
    0.02431289, 0.02426579, 0.02446692, 0.02466582, 0.02574264, 0.02570372, 
    0.0256646, 0.02458168, 0.02382922, 0.02384226, 0.02396953, 0.02550958, 
    0.02572503, 0.02584598, 0.02487706, 0.02464721, 0.02526651, 0.02575096, 
    0.02412141, 0.02290771, 0.02215732, 0.02143294, 0.02143291, 0.02101452, 
    0.02066664, 0.02037749, 0.01870454, 0.0186965, 0.01906431, 0.02013641, 
    0.02394161, 0.02688285, 0.02832414, 0.02573709, 0.02113718, 0.01805269, 
    0.01717715, 0.01665929, 0.01615642, 0.01544068, 0.01437015, 0.01272929, 
    0.01074145, 0.009609379, 0.008556479, 0.007466472, 0.006302336, 
    0.005434135, 0.004866909, 0.004393699, 0.003876376, 0.003291233, 
    0.002999067, 0.002735035, 0.002622703, 0.002827166, 0.003034141, 
    0.003208597, 0.003258205, 0.003797312, 0.004629524, 0.005489939, 
    0.006688516, 0.008302335, 0.009947208, 0.01123536, 0.01326224, 
    0.01621752, 0.01935857, 0.02437663, 0.02770725, 0.03098375, 0.03268769, 
    0.03439434, 0.03793161, 0.04149189, 0.04987805, 0.05329436, 0.05671964, 
    0.05980025, 0.06213039, 0.06423856, 0.06651532, 0.06792332,
  0.06754619, 0.06901011, 0.07052105, 0.07250084, 0.07317252, 0.07269854, 
    0.07193017, 0.06814124, 0.06486051, 0.06325093, 0.06187822, 0.06214299, 
    0.06048862, 0.05807293, 0.05530138, 0.05326088, 0.05246096, 0.05152563, 
    0.050584, 0.05001541, 0.04975102, 0.04957113, 0.04951182, 0.0496801, 
    0.05034476, 0.05070013, 0.05031003, 0.04991456, 0.04987581, 0.05015263, 
    0.05040077, 0.05046925, 0.05039139, 0.05025173, 0.05024201, 0.05018639, 
    0.04956372, 0.04853476, 0.04771434, 0.0468066, 0.04579133, 0.04520971, 
    0.0451209, 0.04487876, 0.04472185, 0.04417371, 0.04364455, 0.04312055, 
    0.04188428, 0.03998457, 0.03933341, 0.03875482, 0.03817626, 0.03804146, 
    0.03758141, 0.03710939, 0.03658048, 0.03549708, 0.03492251, 0.03434598, 
    0.03386521, 0.03340612, 0.03290759, 0.03241, 0.03145873, 0.03107864, 
    0.03069717, 0.03036531, 0.03009453, 0.02980048, 0.02950426, 0.02923569, 
    0.02898544, 0.02860078, 0.02821183, 0.02729381, 0.02697922, 0.02682372, 
    0.02663558, 0.02587292, 0.02611782, 0.02669621, 0.02734478, 0.02819265, 
    0.02691229, 0.02647226, 0.02592054, 0.02580617, 0.02607857, 0.02602792, 
    0.02589624, 0.02580715, 0.02563419, 0.02545389, 0.02548789, 0.0256283, 
    0.02596074, 0.0264041, 0.02688691, 0.02718298, 0.02727945, 0.0272108, 
    0.02685509, 0.02637222, 0.02583938, 0.02547011, 0.02515875, 0.02489456, 
    0.02471253, 0.02463353, 0.0245773, 0.02448732, 0.0243098, 0.02430666, 
    0.02438246, 0.02448451, 0.02463452, 0.02451052, 0.02446442, 0.02443596, 
    0.02424257, 0.02393654, 0.02389609, 0.02387558, 0.02390629, 0.02399435, 
    0.02409219, 0.02419362, 0.02438867, 0.02457893, 0.02469357, 0.02481015, 
    0.02499556, 0.02507175, 0.02512661, 0.02518191, 0.02512187, 0.02513179, 
    0.02514151, 0.02512396, 0.02509641, 0.02509474, 0.02509254, 0.02504757, 
    0.02493788, 0.02494274, 0.02494425, 0.02502898, 0.02506929, 0.02507411, 
    0.02507956, 0.02510817, 0.02514768, 0.02520655, 0.02525907, 0.0252763, 
    0.02532068, 0.02541765, 0.02551991, 0.02574091, 0.0259082, 0.02598036, 
    0.0260196, 0.02601862, 0.0258229, 0.02548225, 0.02522106, 0.02502916, 
    0.02485531, 0.02467266, 0.02448116, 0.02435733, 0.02424393, 0.02414224, 
    0.0240377, 0.02391729, 0.02379143, 0.02375047, 0.02377704, 0.02387065, 
    0.02399197, 0.02409325, 0.0240986, 0.0240751, 0.02397824, 0.0238321, 
    0.02379128, 0.02378373, 0.02384057, 0.02397133, 0.0240153, 0.02405418, 
    0.02406369, 0.02397059, 0.02382755, 0.0236851, 0.02365163, 0.02328233, 
    0.02289636, 0.02250803, 0.02160847, 0.0215038, 0.02153222, 0.02156028, 
    0.02176996, 0.02180492, 0.02197122, 0.02213881, 0.02353822, 0.02353702, 
    0.0235366, 0.02333925, 0.02230904, 0.02222032, 0.02212896, 0.02278108, 
    0.02319631, 0.0230052, 0.02279502, 0.02242705, 0.02271876, 0.02257772, 
    0.02235473, 0.02183738, 0.02164681, 0.02155683, 0.02158505, 0.02205621, 
    0.02099702, 0.02033324, 0.01956575, 0.01830898, 0.01749018, 0.01743846, 
    0.01747232, 0.01985799, 0.02231269, 0.02320748, 0.02213136, 0.02072568, 
    0.01719876, 0.014407, 0.0143607, 0.01379747, 0.01265461, 0.01098657, 
    0.008992876, 0.007778152, 0.006947781, 0.006146738, 0.005373012, 
    0.004839631, 0.004400796, 0.003953747, 0.003566006, 0.00316559, 
    0.002813326, 0.002580114, 0.002542072, 0.002555315, 0.002654122, 
    0.00262689, 0.003091748, 0.003648863, 0.004359953, 0.005450838, 
    0.006936263, 0.008444613, 0.01021706, 0.01233847, 0.01485038, 0.01738786, 
    0.02163834, 0.0256655, 0.02824337, 0.03083261, 0.03061048, 0.03194663, 
    0.03427361, 0.03661764, 0.03907908, 0.04241159, 0.04573719, 0.05000557, 
    0.05650171, 0.05956403, 0.06268977, 0.06574261,
  0.06432424, 0.06720491, 0.06865314, 0.07009163, 0.06906261, 0.06573682, 
    0.06420355, 0.06269938, 0.06010622, 0.05749011, 0.05705084, 0.05648764, 
    0.05606746, 0.0540185, 0.04943351, 0.04764833, 0.04609482, 0.04499478, 
    0.04460786, 0.04394945, 0.04330729, 0.04277757, 0.04267951, 0.04350043, 
    0.04416487, 0.04447359, 0.04465724, 0.04458719, 0.04459614, 0.04470744, 
    0.0446789, 0.04478458, 0.0450909, 0.04538969, 0.04577741, 0.04585421, 
    0.04574833, 0.04569335, 0.04551088, 0.04495698, 0.04418568, 0.04338865, 
    0.04253808, 0.04199865, 0.04135152, 0.04059326, 0.03983339, 0.03981707, 
    0.0395984, 0.0388812, 0.03815413, 0.03741755, 0.03670983, 0.03616117, 
    0.03561321, 0.03502479, 0.03496, 0.03457513, 0.03417066, 0.03375838, 
    0.03332137, 0.0328866, 0.03245031, 0.032012, 0.03095711, 0.0306032, 
    0.03025145, 0.02989952, 0.02954273, 0.02938975, 0.02923563, 0.0290976, 
    0.02867073, 0.02817049, 0.02795925, 0.02777134, 0.02769539, 0.0276113, 
    0.02754459, 0.0275075, 0.02890138, 0.03064916, 0.03020357, 0.02958504, 
    0.02831351, 0.02628637, 0.02589808, 0.02561687, 0.02534497, 0.02519784, 
    0.02524357, 0.02531031, 0.02525844, 0.02521731, 0.02523206, 0.02551545, 
    0.0257601, 0.02593312, 0.02608918, 0.02631093, 0.02630857, 0.02606014, 
    0.02585778, 0.02570037, 0.02559861, 0.02544191, 0.02523595, 0.02504476, 
    0.024862, 0.02466411, 0.02448723, 0.02438392, 0.02429424, 0.02423028, 
    0.02420283, 0.02422597, 0.02423158, 0.02421767, 0.02419012, 0.02403514, 
    0.02391403, 0.02390384, 0.02388651, 0.02398344, 0.02409387, 0.02413217, 
    0.02417239, 0.0242055, 0.02427921, 0.02432758, 0.02437907, 0.02443222, 
    0.02453103, 0.02456001, 0.02458817, 0.02461706, 0.02459419, 0.0245918, 
    0.02458906, 0.02458745, 0.0246784, 0.02466207, 0.02464037, 0.02461468, 
    0.02448489, 0.02450892, 0.02451549, 0.02452158, 0.02448556, 0.02441995, 
    0.02442939, 0.02443746, 0.02447433, 0.02451899, 0.02456662, 0.02460827, 
    0.0246182, 0.02464297, 0.02481709, 0.02492521, 0.02501816, 0.02510063, 
    0.02510072, 0.02502368, 0.02491734, 0.02476969, 0.02456302, 0.02458281, 
    0.0245419, 0.02440611, 0.02420726, 0.02395662, 0.02378269, 0.02369505, 
    0.02362235, 0.02358981, 0.0236392, 0.02367647, 0.02369788, 0.02363636, 
    0.02356213, 0.02347887, 0.02340558, 0.02334896, 0.02332875, 0.0233229, 
    0.02348228, 0.02352866, 0.02343919, 0.02333887, 0.02320386, 0.02295638, 
    0.02282476, 0.0228116, 0.02280006, 0.02310486, 0.02332492, 0.02312779, 
    0.02291564, 0.02234265, 0.02098214, 0.02095618, 0.02094866, 0.02122315, 
    0.02329466, 0.02336278, 0.02341668, 0.02347468, 0.02171832, 0.02175779, 
    0.02180169, 0.02182678, 0.02277332, 0.02344465, 0.02354606, 0.02364339, 
    0.02215734, 0.02084525, 0.02053693, 0.02018147, 0.0215186, 0.02320549, 
    0.02330038, 0.02332532, 0.02279756, 0.02167057, 0.02045985, 0.0194148, 
    0.01811194, 0.01778897, 0.01976434, 0.0197164, 0.01942237, 0.01733086, 
    0.01424232, 0.01313419, 0.01334077, 0.0136545, 0.01414917, 0.01134213, 
    0.009285202, 0.008344252, 0.008146929, 0.008697787, 0.008336323, 
    0.007005626, 0.006153633, 0.005477738, 0.005028244, 0.004716283, 
    0.004559075, 0.004458565, 0.004349956, 0.004444494, 0.004747784, 
    0.004772285, 0.004495458, 0.00415651, 0.003259225, 0.002972451, 
    0.003299899, 0.003723026, 0.004234046, 0.005251154, 0.00652604, 
    0.007628124, 0.008722969, 0.009755683, 0.01145298, 0.01350412, 
    0.01559616, 0.0179244, 0.02171761, 0.0241202, 0.02649052, 0.02900192, 
    0.03038733, 0.03197798, 0.0335915, 0.03520909, 0.03321731, 0.03590465, 
    0.03857788, 0.04129177, 0.049008, 0.05279956, 0.05611916, 0.05945197,
  0.05142672, 0.05920278, 0.06141463, 0.0622282, 0.06300874, 0.06075977, 
    0.0553074, 0.05345191, 0.05210589, 0.05132248, 0.05386798, 0.05425352, 
    0.05134512, 0.04870514, 0.04520807, 0.04128564, 0.04181827, 0.04178377, 
    0.04111006, 0.04023947, 0.03932558, 0.03883706, 0.0384794, 0.03852906, 
    0.03875386, 0.03921781, 0.03965253, 0.04022895, 0.04068463, 0.04089744, 
    0.04108803, 0.04128277, 0.04152212, 0.04172226, 0.04197689, 0.04243679, 
    0.04276121, 0.04274582, 0.04264693, 0.04237675, 0.0417175, 0.04128184, 
    0.04093931, 0.04054832, 0.04018831, 0.0392455, 0.03774492, 0.03692814, 
    0.03632194, 0.03572971, 0.03489355, 0.03429188, 0.03386806, 0.03345235, 
    0.03322707, 0.03320328, 0.03283455, 0.03250579, 0.03217603, 0.03187186, 
    0.0316067, 0.0313035, 0.03099774, 0.03068944, 0.03047019, 0.03024465, 
    0.03002128, 0.0298001, 0.02967314, 0.02949551, 0.02949749, 0.02951889, 
    0.02947464, 0.03068146, 0.03133865, 0.03148464, 0.03163507, 0.03152752, 
    0.03056686, 0.03018831, 0.02979763, 0.02911287, 0.02761961, 0.02664849, 
    0.02637933, 0.02604283, 0.02575476, 0.02538298, 0.02472305, 0.02437621, 
    0.0242152, 0.02415049, 0.0243496, 0.0246248, 0.02485169, 0.02501227, 
    0.02516272, 0.02533815, 0.02544728, 0.0254701, 0.02547989, 0.02548377, 
    0.02541151, 0.02532491, 0.02527188, 0.02519128, 0.02506397, 0.02495582, 
    0.02485378, 0.02473575, 0.0245966, 0.02440971, 0.02418746, 0.02405391, 
    0.02399399, 0.02394454, 0.02390796, 0.02386922, 0.02380542, 0.02381938, 
    0.02385229, 0.02391174, 0.02422279, 0.02439162, 0.02441444, 0.02443916, 
    0.02442291, 0.02426982, 0.0242569, 0.02425548, 0.02425635, 0.02422152, 
    0.02416373, 0.02415838, 0.02415345, 0.02414897, 0.02414539, 0.02412532, 
    0.02410459, 0.02408318, 0.02403929, 0.0239858, 0.02396541, 0.02394398, 
    0.02393445, 0.02405082, 0.02406725, 0.0240599, 0.02405355, 0.02401606, 
    0.02400397, 0.02400069, 0.02399432, 0.0239898, 0.02400042, 0.02395798, 
    0.02393268, 0.02391512, 0.02390527, 0.02395472, 0.02403563, 0.02403854, 
    0.02402249, 0.02401772, 0.02399438, 0.02394043, 0.02389758, 0.02387101, 
    0.02385632, 0.0237856, 0.0236926, 0.02360301, 0.02363611, 0.02376689, 
    0.02387559, 0.02392997, 0.02386214, 0.02377312, 0.02361907, 0.02348783, 
    0.02338585, 0.02331846, 0.02324537, 0.02318658, 0.02319645, 0.02330789, 
    0.02328128, 0.02319433, 0.02308184, 0.02265408, 0.0221947, 0.02208385, 
    0.02202542, 0.0220153, 0.0223986, 0.02266765, 0.02260782, 0.02253484, 
    0.02238298, 0.02162528, 0.02151209, 0.02152872, 0.02154703, 0.02240017, 
    0.02345835, 0.02342098, 0.02338395, 0.02334724, 0.01948638, 0.01974499, 
    0.02000492, 0.02026617, 0.02402579, 0.02713908, 0.026878, 0.02659769, 
    0.02576854, 0.02002352, 0.01827106, 0.01750703, 0.01671127, 0.01708778, 
    0.01817402, 0.01786245, 0.01749505, 0.01717026, 0.01550131, 0.01442018, 
    0.01471775, 0.01505959, 0.01611498, 0.01785584, 0.01678555, 0.01580269, 
    0.01515849, 0.01466577, 0.01402383, 0.01318063, 0.01235935, 0.01155246, 
    0.0106912, 0.01004441, 0.009551477, 0.009150258, 0.008737398, 
    0.008259049, 0.007821096, 0.007220573, 0.006595217, 0.005971406, 
    0.005338598, 0.005047597, 0.004816298, 0.004677254, 0.004684474, 
    0.004967692, 0.0054119, 0.004893904, 0.004601351, 0.004570424, 
    0.004538418, 0.00470324, 0.005391238, 0.006174739, 0.006993258, 
    0.007841218, 0.008657712, 0.009936516, 0.01161329, 0.01331492, 
    0.01524387, 0.01772006, 0.01964409, 0.02156868, 0.02351143, 0.02616604, 
    0.02861498, 0.02996917, 0.03132657, 0.03268716, 0.03037516, 0.0322583, 
    0.03412825, 0.03598497, 0.03928004, 0.04279252, 0.04556112, 0.04828117,
  0.03847485, 0.04110792, 0.0463425, 0.04708233, 0.04722502, 0.04734449, 
    0.04663682, 0.04521867, 0.04446444, 0.04363136, 0.04277644, 0.04172786, 
    0.03899615, 0.03665823, 0.03585437, 0.03558077, 0.03544636, 0.03656268, 
    0.03704237, 0.0373954, 0.03758242, 0.03745729, 0.03718186, 0.03657988, 
    0.03609538, 0.03643814, 0.03694521, 0.03726755, 0.03742443, 0.03753565, 
    0.03758099, 0.03766956, 0.03802517, 0.03837276, 0.03860105, 0.03875348, 
    0.03896593, 0.03924499, 0.03933499, 0.03897729, 0.03865741, 0.0383017, 
    0.03772256, 0.03788979, 0.03836227, 0.03814375, 0.03767982, 0.03704932, 
    0.03597499, 0.03464642, 0.03393264, 0.03332953, 0.0327286, 0.03206329, 
    0.03183177, 0.03165711, 0.03135238, 0.03104898, 0.03074714, 0.03047037, 
    0.03026807, 0.03007289, 0.02987692, 0.02968017, 0.02996774, 0.02983464, 
    0.02970255, 0.02957147, 0.02936604, 0.02862445, 0.02877274, 0.02897118, 
    0.02917012, 0.02983122, 0.03282897, 0.03333935, 0.03315891, 0.03295919, 
    0.03233284, 0.02878195, 0.02597831, 0.02515129, 0.02458025, 0.02437049, 
    0.02526468, 0.02602575, 0.0258207, 0.02563463, 0.02546612, 0.02514837, 
    0.02491471, 0.02473765, 0.0246012, 0.02454823, 0.02451207, 0.02457316, 
    0.02465742, 0.02466741, 0.02463405, 0.02460752, 0.02460324, 0.02462778, 
    0.02466348, 0.02465892, 0.0246341, 0.02457983, 0.02452167, 0.02445335, 
    0.02434844, 0.02420719, 0.02404888, 0.02394062, 0.02391276, 0.02388391, 
    0.02389306, 0.02396999, 0.02406373, 0.02410857, 0.02413633, 0.02414607, 
    0.02412653, 0.02418358, 0.02425126, 0.02427566, 0.02430324, 0.02433939, 
    0.02424937, 0.024189, 0.02416567, 0.02414254, 0.02412357, 0.02413685, 
    0.02412067, 0.02410273, 0.02408481, 0.02406692, 0.02403193, 0.02399306, 
    0.0239539, 0.02391443, 0.02386231, 0.02365194, 0.02361446, 0.02358967, 
    0.02356347, 0.02355598, 0.02359611, 0.02359209, 0.02359021, 0.02358788, 
    0.0235854, 0.02363809, 0.02367395, 0.02366176, 0.02364326, 0.02360535, 
    0.02344638, 0.02332524, 0.02334658, 0.02337011, 0.02338911, 0.02343551, 
    0.02344085, 0.02342413, 0.02339716, 0.02336846, 0.02332518, 0.02327531, 
    0.02322437, 0.02317701, 0.02314566, 0.02313109, 0.02312331, 0.02316744, 
    0.02327546, 0.02335058, 0.02322653, 0.02307801, 0.0229938, 0.02292365, 
    0.02285389, 0.02277903, 0.02271721, 0.02270082, 0.02264287, 0.02258112, 
    0.02251349, 0.02223296, 0.02187829, 0.02172385, 0.02162528, 0.02152955, 
    0.02157162, 0.02178386, 0.02184639, 0.02182862, 0.02180997, 0.02178352, 
    0.02157007, 0.02150659, 0.02151114, 0.02151847, 0.02154171, 0.02192056, 
    0.0219329, 0.02190264, 0.0218706, 0.02183678, 0.02120878, 0.02138775, 
    0.02156175, 0.02173076, 0.02223435, 0.02467864, 0.02413959, 0.02357619, 
    0.02301096, 0.02148155, 0.01737393, 0.01663348, 0.01618449, 0.01575332, 
    0.01573002, 0.01742921, 0.01856386, 0.01852477, 0.01824982, 0.01758686, 
    0.0167116, 0.01636652, 0.01652502, 0.01621999, 0.01591862, 0.01529026, 
    0.01478525, 0.01436477, 0.01405271, 0.01388597, 0.01393804, 0.01394395, 
    0.01394991, 0.01394801, 0.01389513, 0.01361674, 0.01316657, 0.01245308, 
    0.01138401, 0.01034814, 0.0096088, 0.009030087, 0.008653787, 0.00834544, 
    0.008293367, 0.008495761, 0.008771778, 0.008844472, 0.008647338, 
    0.008458749, 0.008063747, 0.007497886, 0.007230874, 0.007433236, 
    0.007721988, 0.00803464, 0.00838044, 0.00915941, 0.0102584, 0.01147027, 
    0.01271104, 0.01472694, 0.01830762, 0.01980571, 0.02116246, 0.02253879, 
    0.02371128, 0.02381615, 0.0249101, 0.02598137, 0.02705609, 0.02813425, 
    0.02873634, 0.02993014, 0.03111479, 0.03229026, 0.0333678, 0.03323612, 
    0.03497387, 0.03675913,
  0.03116049, 0.03204077, 0.03302708, 0.03437229, 0.03448213, 0.03474777, 
    0.03498875, 0.03520464, 0.0355476, 0.03694298, 0.03785599, 0.03761312, 
    0.03719803, 0.03671156, 0.03564195, 0.03440396, 0.03391142, 0.03371207, 
    0.0335525, 0.03344369, 0.03350204, 0.03332509, 0.03328286, 0.03333006, 
    0.03353621, 0.03373927, 0.03394285, 0.03426212, 0.03439821, 0.03431451, 
    0.03428658, 0.03425782, 0.03423139, 0.03428612, 0.03430551, 0.03436903, 
    0.03458771, 0.03473, 0.03485247, 0.03495925, 0.0348521, 0.03424698, 
    0.03371175, 0.03346899, 0.0332273, 0.03301802, 0.03299476, 0.0327994, 
    0.03241185, 0.03214288, 0.03185623, 0.03155228, 0.03125309, 0.03071684, 
    0.03041974, 0.03015713, 0.0298926, 0.02962616, 0.02932123, 0.02911573, 
    0.02896508, 0.02881453, 0.02866407, 0.02851371, 0.02868327, 0.02859416, 
    0.02850572, 0.02841794, 0.02833083, 0.02796548, 0.02783911, 0.02796154, 
    0.02807241, 0.02817158, 0.02848624, 0.0297063, 0.02904859, 0.02854112, 
    0.02803332, 0.02752514, 0.02640178, 0.02648288, 0.0268433, 0.0266249, 
    0.02634661, 0.02606642, 0.025818, 0.02568057, 0.02550518, 0.02531768, 
    0.02515131, 0.0249916, 0.02479877, 0.02468389, 0.02460416, 0.02457203, 
    0.02453166, 0.02449766, 0.02446728, 0.02443814, 0.02442476, 0.02440995, 
    0.02437034, 0.0243282, 0.02431938, 0.02434644, 0.02436131, 0.02435008, 
    0.02425975, 0.02417608, 0.0240905, 0.02401143, 0.02397412, 0.0240233, 
    0.02405497, 0.02403535, 0.02402383, 0.02402208, 0.02405592, 0.0241215, 
    0.02410318, 0.02407618, 0.02405373, 0.02403571, 0.02396271, 0.02391146, 
    0.02389381, 0.02387626, 0.02385977, 0.02384435, 0.02388673, 0.02390014, 
    0.02388497, 0.02386995, 0.0238551, 0.02384041, 0.02387333, 0.02382571, 
    0.02377821, 0.02373084, 0.02368361, 0.0235422, 0.0233867, 0.02334577, 
    0.0233049, 0.02326409, 0.02322299, 0.02320797, 0.02322595, 0.02321521, 
    0.02320211, 0.02318662, 0.02319611, 0.02323866, 0.02324452, 0.0232096, 
    0.02316408, 0.02311037, 0.02304645, 0.02297177, 0.02289794, 0.02283024, 
    0.02276568, 0.02269837, 0.02262384, 0.02256597, 0.0225352, 0.02251011, 
    0.02251753, 0.02251802, 0.02251898, 0.02253085, 0.02256727, 0.02259557, 
    0.02258491, 0.02256269, 0.0225152, 0.02243883, 0.02234364, 0.02222181, 
    0.02214615, 0.02208401, 0.02201715, 0.02195895, 0.02190297, 0.02183429, 
    0.02174501, 0.02164074, 0.02153732, 0.02143166, 0.0212357, 0.02104066, 
    0.0210075, 0.02096822, 0.02093331, 0.02090266, 0.02087508, 0.02079993, 
    0.02077456, 0.02075839, 0.02074461, 0.02073319, 0.02072529, 0.02081923, 
    0.02085892, 0.02089808, 0.02093668, 0.02097476, 0.02110649, 0.02108732, 
    0.02106537, 0.02104061, 0.02101305, 0.02086075, 0.02012085, 0.01976513, 
    0.01942058, 0.01908734, 0.01866866, 0.0184662, 0.01933246, 0.01922651, 
    0.01913789, 0.01906716, 0.0187754, 0.01542789, 0.01266247, 0.01230219, 
    0.01237057, 0.01265488, 0.01385176, 0.01553888, 0.01572488, 0.01554793, 
    0.01560835, 0.01567926, 0.01584596, 0.01633905, 0.01663085, 0.01684009, 
    0.01679426, 0.01652745, 0.01624988, 0.01588551, 0.01521437, 0.01444091, 
    0.01390708, 0.01338342, 0.01293249, 0.01276066, 0.01271481, 0.01281016, 
    0.01288809, 0.01279734, 0.01271731, 0.01269621, 0.01248421, 0.01166357, 
    0.0111081, 0.01097474, 0.01090065, 0.01089953, 0.01091591, 0.01126785, 
    0.01166741, 0.01224464, 0.01288472, 0.01358629, 0.01408686, 0.01667548, 
    0.01815899, 0.01939648, 0.02065189, 0.02192501, 0.02277315, 0.0224607, 
    0.02327758, 0.02409551, 0.02491448, 0.02573448, 0.02695155, 0.02766889, 
    0.02838088, 0.02908748, 0.02978868, 0.02942163, 0.02928225, 0.03024083,
  0.02859143, 0.02903524, 0.02946824, 0.02989028, 0.02982533, 0.02976386, 
    0.03001019, 0.03031216, 0.03058665, 0.0308331, 0.03124301, 0.03121706, 
    0.03098491, 0.03083301, 0.03083541, 0.03086166, 0.0308911, 0.0309304, 
    0.03098739, 0.03102908, 0.03106244, 0.0311223, 0.03121781, 0.03131116, 
    0.03138568, 0.03151457, 0.03161928, 0.03169376, 0.03174987, 0.03177935, 
    0.03175284, 0.03166381, 0.03159254, 0.03150043, 0.03138501, 0.03120656, 
    0.03097204, 0.0308803, 0.03094928, 0.03091267, 0.03081788, 0.03070948, 
    0.030594, 0.03060874, 0.03062937, 0.030535, 0.03039948, 0.03021037, 
    0.03000532, 0.0297847, 0.0294951, 0.02918697, 0.02908205, 0.02888669, 
    0.02868752, 0.02848461, 0.02827799, 0.02809713, 0.0279123, 0.02777556, 
    0.02763867, 0.02750145, 0.02736391, 0.02722606, 0.02699281, 0.02694565, 
    0.02689898, 0.02685278, 0.02680707, 0.02676224, 0.0268905, 0.02703815, 
    0.02702926, 0.02701657, 0.02700004, 0.02697962, 0.02665484, 0.02640632, 
    0.02631169, 0.0262231, 0.02614234, 0.02606959, 0.02609469, 0.02586549, 
    0.02558313, 0.02539865, 0.02527869, 0.02515909, 0.02504683, 0.02493678, 
    0.02485375, 0.02486958, 0.02496212, 0.02504189, 0.02506961, 0.0250862, 
    0.02502397, 0.02489922, 0.02476062, 0.02462827, 0.02453638, 0.02448257, 
    0.0244413, 0.02441808, 0.02438545, 0.02435529, 0.02433126, 0.02431214, 
    0.0243024, 0.0242924, 0.02427809, 0.0242639, 0.02424501, 0.02422864, 
    0.02420845, 0.02413483, 0.02402755, 0.0239309, 0.02388595, 0.02384694, 
    0.02381076, 0.02377734, 0.02373599, 0.0236322, 0.0235069, 0.02346364, 
    0.02342222, 0.0233826, 0.02334476, 0.02334335, 0.02337215, 0.02334566, 
    0.02331956, 0.02329403, 0.02326905, 0.02324462, 0.02323907, 0.02320355, 
    0.02316824, 0.02313315, 0.02309828, 0.02306346, 0.02299701, 0.02299331, 
    0.02296448, 0.02293571, 0.02290698, 0.0228783, 0.02287595, 0.02286288, 
    0.02282701, 0.02278919, 0.02274726, 0.02270113, 0.02265471, 0.02257812, 
    0.02248123, 0.02239686, 0.02233675, 0.02227514, 0.02221344, 0.02214542, 
    0.02207125, 0.02199381, 0.02191495, 0.02184869, 0.02180183, 0.02176351, 
    0.02176051, 0.0218004, 0.02185111, 0.0218986, 0.02193968, 0.02196672, 
    0.02196698, 0.02193509, 0.02189965, 0.02185949, 0.02180972, 0.0217272, 
    0.02160693, 0.02153746, 0.02154571, 0.02151259, 0.02144836, 0.02137868, 
    0.02130117, 0.02114937, 0.02091761, 0.02066304, 0.02055749, 0.020499, 
    0.02044032, 0.02038143, 0.02039977, 0.02047405, 0.02038639, 0.02031608, 
    0.02024709, 0.0201794, 0.02011298, 0.01982136, 0.01955123, 0.01958281, 
    0.01961564, 0.01964925, 0.01968365, 0.01971883, 0.02115854, 0.0210537, 
    0.02094954, 0.02084604, 0.02074323, 0.02063869, 0.01938718, 0.01850805, 
    0.01831384, 0.01812056, 0.01792825, 0.01773691, 0.01859528, 0.01943923, 
    0.01932642, 0.01897024, 0.01862333, 0.01828592, 0.01758219, 0.01802312, 
    0.01869873, 0.01891641, 0.01862711, 0.01826352, 0.01789658, 0.01729777, 
    0.01653061, 0.01615849, 0.01603849, 0.01587961, 0.01567883, 0.01548344, 
    0.01542173, 0.01553988, 0.01564997, 0.01575314, 0.01564885, 0.01536343, 
    0.01512172, 0.01488975, 0.01480602, 0.01480463, 0.01482557, 0.01486891, 
    0.01497113, 0.01510017, 0.01524004, 0.01540487, 0.01555213, 0.01569225, 
    0.01580384, 0.01600369, 0.01629865, 0.01649805, 0.01648684, 0.0165364, 
    0.01662303, 0.01674592, 0.01660145, 0.01585042, 0.01569869, 0.01627078, 
    0.01686135, 0.01747017, 0.01809698, 0.01963639, 0.02230195, 0.02296397, 
    0.02362408, 0.02428721, 0.02495335, 0.02562247, 0.02494939, 0.02539795, 
    0.02584403, 0.02628764, 0.02672875, 0.0271674, 0.02754664, 0.02813695,
  0.02717811, 0.02745047, 0.02771812, 0.027981, 0.02823903, 0.02848559, 
    0.02841942, 0.02843807, 0.02854226, 0.02867414, 0.02879724, 0.0289079, 
    0.02900582, 0.02905509, 0.02908667, 0.02908042, 0.02905222, 0.02907562, 
    0.02911664, 0.02915362, 0.02918636, 0.02920832, 0.02921126, 0.02921506, 
    0.02920486, 0.02916411, 0.02910391, 0.02905493, 0.02903215, 0.0290106, 
    0.0289863, 0.02896134, 0.02890602, 0.02881371, 0.02868465, 0.02859144, 
    0.02852503, 0.02845393, 0.02837832, 0.02833907, 0.02835862, 0.0283575, 
    0.0283306, 0.02832827, 0.02828818, 0.02823856, 0.02817963, 0.02811412, 
    0.02807366, 0.02797669, 0.02778792, 0.02765483, 0.02752141, 0.02738539, 
    0.02724682, 0.02710573, 0.02690324, 0.02687751, 0.02678707, 0.02669388, 
    0.02659996, 0.02650531, 0.02640994, 0.02631384, 0.02602003, 0.02600457, 
    0.02598961, 0.02597512, 0.02596113, 0.02594764, 0.025945, 0.02632624, 
    0.02642482, 0.02636954, 0.0263139, 0.02625789, 0.02620149, 0.02614421, 
    0.02604792, 0.02578103, 0.02550464, 0.02534323, 0.02518759, 0.02503152, 
    0.02487502, 0.02471315, 0.02462389, 0.02457304, 0.02455387, 0.02450513, 
    0.0244495, 0.02439671, 0.02434689, 0.0243525, 0.02445825, 0.02449498, 
    0.02447568, 0.02446241, 0.02447649, 0.02447688, 0.02444846, 0.02441919, 
    0.02438645, 0.02434386, 0.02430547, 0.02426161, 0.02420967, 0.02416421, 
    0.02412029, 0.0240767, 0.02403347, 0.0239949, 0.02398207, 0.02397056, 
    0.02396527, 0.02391934, 0.02386473, 0.02381058, 0.02375689, 0.02370491, 
    0.023678, 0.02363296, 0.0235372, 0.02347076, 0.02340562, 0.02334103, 
    0.02327698, 0.02321348, 0.02306662, 0.02300966, 0.0229676, 0.02292475, 
    0.02288218, 0.02283988, 0.02279785, 0.0227561, 0.0226821, 0.02265812, 
    0.02263406, 0.02260992, 0.02258569, 0.02256137, 0.02253959, 0.02263227, 
    0.02271273, 0.0226818, 0.02265005, 0.02261747, 0.02258404, 0.02254926, 
    0.02248003, 0.02231489, 0.02215576, 0.02208263, 0.02201247, 0.02194069, 
    0.02186724, 0.02180281, 0.02179069, 0.02178371, 0.02178303, 0.02177245, 
    0.02175355, 0.02173632, 0.02172085, 0.02169665, 0.02165644, 0.0216426, 
    0.0216418, 0.02163127, 0.02159807, 0.02156734, 0.02155049, 0.02155191, 
    0.02156621, 0.02158276, 0.0215824, 0.02154743, 0.02146771, 0.02138873, 
    0.02131587, 0.02124014, 0.02116166, 0.02110255, 0.02110001, 0.02109305, 
    0.02107784, 0.02100828, 0.02093466, 0.02085889, 0.02078101, 0.02070319, 
    0.02066383, 0.02070422, 0.02082928, 0.02077783, 0.02072036, 0.02066133, 
    0.02060078, 0.02053873, 0.02036004, 0.01978816, 0.01974849, 0.01972397, 
    0.0197004, 0.01967779, 0.01965612, 0.01963539, 0.02068012, 0.02061231, 
    0.0205454, 0.02047937, 0.02041425, 0.02035004, 0.02025324, 0.01910129, 
    0.01925078, 0.01923904, 0.01922829, 0.01921853, 0.01920977, 0.01921535, 
    0.01965753, 0.01896068, 0.01803057, 0.01777232, 0.01754469, 0.01731339, 
    0.01707836, 0.01693979, 0.01684237, 0.01675878, 0.01666615, 0.01657382, 
    0.01649376, 0.01641222, 0.01632918, 0.01625288, 0.01618451, 0.01600101, 
    0.01574976, 0.0155245, 0.01533473, 0.01521139, 0.01516333, 0.01513699, 
    0.01515533, 0.01526198, 0.01541175, 0.01552237, 0.01558393, 0.01571513, 
    0.01587524, 0.01604595, 0.01622677, 0.01642071, 0.01658149, 0.01676876, 
    0.01701759, 0.01735488, 0.01765667, 0.01795467, 0.01824903, 0.01853977, 
    0.0188448, 0.01884787, 0.01839853, 0.01873756, 0.01910364, 0.0194774, 
    0.01985876, 0.02024758, 0.02103092, 0.02238796, 0.02286304, 0.02331248, 
    0.02376502, 0.02422064, 0.02467932, 0.02514105, 0.02389812, 0.0242088, 
    0.02451838, 0.02482683, 0.02513416, 0.02544035, 0.02576137, 0.02662579,
  0.02539306, 0.02580472, 0.02600617, 0.02616375, 0.02631673, 0.02646505, 
    0.0266086, 0.02674729, 0.02684037, 0.02681888, 0.02686017, 0.02687976, 
    0.02690562, 0.02694103, 0.02697397, 0.02700437, 0.02704024, 0.02709822, 
    0.02716078, 0.02719978, 0.02722083, 0.02724023, 0.02731203, 0.02735891, 
    0.02737266, 0.02738256, 0.0273884, 0.02736278, 0.02730842, 0.027252, 
    0.02718284, 0.02710781, 0.02702727, 0.02691575, 0.0267965, 0.02681736, 
    0.02685829, 0.0268898, 0.02690483, 0.02689122, 0.02684634, 0.02679516, 
    0.0267409, 0.02668366, 0.02662068, 0.02653915, 0.02645349, 0.02647696, 
    0.02643422, 0.02636134, 0.02628595, 0.0262081, 0.02612784, 0.02604521, 
    0.02593403, 0.025692, 0.02547832, 0.02542201, 0.02536515, 0.02530776, 
    0.02524982, 0.02519135, 0.02513235, 0.02507282, 0.02541345, 0.02541435, 
    0.02541548, 0.02541685, 0.02541845, 0.02542029, 0.02542237, 0.02542469, 
    0.025477, 0.02556708, 0.02555138, 0.02551201, 0.02547355, 0.02543601, 
    0.0253994, 0.02536375, 0.02526916, 0.02504913, 0.02492274, 0.02482124, 
    0.02475525, 0.02470464, 0.02465708, 0.02461269, 0.02455763, 0.02445954, 
    0.02434112, 0.02423465, 0.02413918, 0.02405652, 0.02400018, 0.02395958, 
    0.02393107, 0.02389992, 0.02386598, 0.02385329, 0.02386178, 0.02386174, 
    0.02386332, 0.02386531, 0.0238676, 0.02386963, 0.02386434, 0.02382522, 
    0.02377779, 0.02372495, 0.02366222, 0.0236119, 0.02358283, 0.02355783, 
    0.02353251, 0.02350688, 0.02346825, 0.02339616, 0.02332191, 0.0233189, 
    0.0233028, 0.0232748, 0.02324592, 0.02321615, 0.02318553, 0.02315406, 
    0.02314165, 0.02300687, 0.02282071, 0.02277466, 0.02272842, 0.02268197, 
    0.02263532, 0.02258848, 0.02254144, 0.0224942, 0.022419, 0.02239885, 
    0.0223784, 0.02235767, 0.02233664, 0.02231531, 0.02229369, 0.02227176, 
    0.02235897, 0.02242925, 0.02238572, 0.02234555, 0.02230469, 0.0222631, 
    0.0222208, 0.02217776, 0.02209124, 0.02192558, 0.02189083, 0.0218773, 
    0.02186411, 0.02185129, 0.02184041, 0.02183155, 0.0218164, 0.02179614, 
    0.02178237, 0.02177127, 0.02176252, 0.02176198, 0.02179664, 0.02181777, 
    0.02181897, 0.02181827, 0.02181553, 0.02179761, 0.02177572, 0.02174324, 
    0.02169149, 0.02163909, 0.0215861, 0.02150916, 0.02141402, 0.02135178, 
    0.02129625, 0.02124001, 0.02117952, 0.02112804, 0.02108838, 0.02105081, 
    0.02101387, 0.02097754, 0.02093164, 0.02086716, 0.02081974, 0.02086162, 
    0.020869, 0.02085653, 0.02084299, 0.02082839, 0.02081276, 0.02079611, 
    0.0207967, 0.02085665, 0.02086829, 0.02083556, 0.02080264, 0.02076952, 
    0.02073622, 0.02070273, 0.02066905, 0.02063518, 0.02000062, 0.01998312, 
    0.01996545, 0.01994762, 0.0199296, 0.01991142, 0.01989306, 0.01987452, 
    0.0206457, 0.02140724, 0.0212262, 0.02104669, 0.02086812, 0.02069051, 
    0.02051389, 0.02033829, 0.01985445, 0.01885293, 0.01894321, 0.01915168, 
    0.0191827, 0.01913303, 0.0190811, 0.0190268, 0.01892328, 0.01870414, 
    0.01844307, 0.01816091, 0.01788518, 0.01761113, 0.01725871, 0.0169591, 
    0.01672583, 0.01650317, 0.01629192, 0.01603704, 0.01589859, 0.01595049, 
    0.01601915, 0.01610876, 0.01621806, 0.01642554, 0.01670913, 0.01687301, 
    0.01704338, 0.01725248, 0.0175016, 0.01772255, 0.01788648, 0.01804625, 
    0.01820799, 0.01837164, 0.01852101, 0.01865856, 0.01883444, 0.01902856, 
    0.01927267, 0.0195291, 0.01979032, 0.02005626, 0.02032682, 0.02060191, 
    0.02090525, 0.02143117, 0.02200879, 0.02228693, 0.02256631, 0.0228469, 
    0.02312871, 0.02341173, 0.02369595, 0.02398136, 0.02348747, 0.02370198, 
    0.02391558, 0.02412825, 0.02434, 0.02455081, 0.02476068, 0.02496961,
  0.02380959, 0.02395286, 0.02417563, 0.02430808, 0.02439949, 0.02447919, 
    0.0245555, 0.02462821, 0.02469724, 0.02476249, 0.0248239, 0.02487991, 
    0.02488024, 0.02487102, 0.02492943, 0.02496924, 0.02498761, 0.02499224, 
    0.0250035, 0.02502368, 0.02504705, 0.02507042, 0.02509343, 0.02514011, 
    0.02520607, 0.02525605, 0.02529051, 0.02530995, 0.02530492, 0.02527776, 
    0.02524086, 0.02519419, 0.02513772, 0.0251027, 0.02508971, 0.02507613, 
    0.02506256, 0.02505353, 0.02505743, 0.02506727, 0.02506958, 0.02505994, 
    0.02503893, 0.0250296, 0.02501448, 0.02499554, 0.0249738, 0.02494917, 
    0.02492172, 0.02489152, 0.02485863, 0.02482293, 0.02477246, 0.02469183, 
    0.02458003, 0.02454804, 0.02452326, 0.02449802, 0.02447232, 0.02444616, 
    0.02441955, 0.02439249, 0.02436498, 0.02433704, 0.02445546, 0.02446228, 
    0.02446923, 0.02447632, 0.02448354, 0.0244909, 0.02449839, 0.02450602, 
    0.02451379, 0.02452919, 0.02463974, 0.02476134, 0.02479288, 0.0247653, 
    0.02473724, 0.02471057, 0.02468535, 0.0246616, 0.02463937, 0.02461749, 
    0.02456331, 0.02451364, 0.0244801, 0.02444355, 0.02440335, 0.02436033, 
    0.02431241, 0.02426445, 0.02421634, 0.02416824, 0.02412108, 0.02406446, 
    0.02399418, 0.02392711, 0.02386312, 0.02380207, 0.02374662, 0.02369389, 
    0.02363885, 0.02358127, 0.02352092, 0.02346071, 0.02341652, 0.02337524, 
    0.02333397, 0.02329539, 0.02326593, 0.02325418, 0.02324951, 0.023247, 
    0.02324409, 0.0231854, 0.02310937, 0.02306359, 0.02301937, 0.02297559, 
    0.02293223, 0.02288927, 0.02284672, 0.02280529, 0.02279416, 0.0228718, 
    0.02293611, 0.02291098, 0.02287931, 0.02284769, 0.02281612, 0.0227846, 
    0.02275313, 0.02272171, 0.02269033, 0.022659, 0.02264987, 0.0226219, 
    0.02259387, 0.0225658, 0.02253768, 0.0225095, 0.02248128, 0.022453, 
    0.02242467, 0.02239412, 0.02232754, 0.02224698, 0.02218978, 0.02215664, 
    0.02212382, 0.02209056, 0.02205685, 0.02202267, 0.02198802, 0.02195305, 
    0.02192337, 0.02189809, 0.02187175, 0.02184221, 0.02180934, 0.02177506, 
    0.02174372, 0.02171289, 0.0216823, 0.02165171, 0.02162021, 0.02160208, 
    0.0216006, 0.02159411, 0.02158254, 0.02156585, 0.02151912, 0.02144313, 
    0.02136369, 0.02128058, 0.02119363, 0.02113103, 0.02109244, 0.02105376, 
    0.02101508, 0.02097855, 0.02094954, 0.0209365, 0.02092971, 0.0209254, 
    0.02092114, 0.02086803, 0.02081007, 0.02078638, 0.02076398, 0.02074176, 
    0.02071973, 0.02069787, 0.02067619, 0.02065419, 0.02062103, 0.02069191, 
    0.02077038, 0.02075995, 0.02074274, 0.02072507, 0.02070696, 0.02068839, 
    0.02066939, 0.02064995, 0.02063007, 0.02060976, 0.02037484, 0.02036062, 
    0.02034642, 0.02033222, 0.02031803, 0.02030385, 0.02028967, 0.02027551, 
    0.02026135, 0.0202447, 0.02017898, 0.02009189, 0.02002157, 0.01997428, 
    0.01992866, 0.01988403, 0.01984042, 0.01979785, 0.01975635, 0.01972283, 
    0.01988046, 0.0199814, 0.01973484, 0.01948096, 0.01923447, 0.01901403, 
    0.01885238, 0.0187478, 0.01866054, 0.01857328, 0.01849212, 0.01839458, 
    0.01826256, 0.01815988, 0.01808599, 0.01804026, 0.01803964, 0.01808859, 
    0.01817596, 0.01830316, 0.01847148, 0.0185875, 0.01865206, 0.01871985, 
    0.01878765, 0.01885546, 0.01892291, 0.0189396, 0.0189597, 0.01900746, 
    0.01908122, 0.01912441, 0.01920605, 0.019353, 0.01950708, 0.0196664, 
    0.01983082, 0.02000022, 0.02017448, 0.02035678, 0.02065312, 0.02086492, 
    0.02109631, 0.02127643, 0.02145086, 0.02162619, 0.02180243, 0.02197955, 
    0.02215756, 0.02233644, 0.02251619, 0.0226968, 0.02270785, 0.02284887, 
    0.02298895, 0.02312811, 0.02326632, 0.02340358, 0.02353989, 0.02367522,
  0.02296175, 0.02303322, 0.02310404, 0.02317419, 0.023235, 0.02324219, 
    0.02319674, 0.02321286, 0.02325384, 0.0232955, 0.02333735, 0.02337689, 
    0.02341405, 0.02344877, 0.02348097, 0.02351059, 0.02353754, 0.02355427, 
    0.02353743, 0.02353961, 0.02356087, 0.02357097, 0.02357064, 0.0235636, 
    0.02355159, 0.02353487, 0.02351377, 0.02349691, 0.02350158, 0.02351793, 
    0.02353545, 0.02354971, 0.02356051, 0.02356803, 0.02357224, 0.02356854, 
    0.02355607, 0.02356588, 0.02360185, 0.02361656, 0.02362437, 0.02363018, 
    0.02363405, 0.02363603, 0.02363617, 0.02363452, 0.02363113, 0.02363053, 
    0.02364127, 0.02366301, 0.02370658, 0.02372177, 0.02371952, 0.02371752, 
    0.02371515, 0.02371241, 0.02370931, 0.02370584, 0.02370202, 0.02369784, 
    0.02369331, 0.02368844, 0.02368322, 0.02367767, 0.02350264, 0.02352058, 
    0.02353864, 0.02355682, 0.02357513, 0.02359356, 0.02361211, 0.02363079, 
    0.0236496, 0.02366854, 0.0236876, 0.0237068, 0.02376038, 0.02388405, 
    0.02400278, 0.02407632, 0.02412697, 0.02414577, 0.02415584, 0.02416614, 
    0.02417669, 0.02418747, 0.0241985, 0.02420977, 0.0242213, 0.02423405, 
    0.024249, 0.02424379, 0.02422059, 0.02419478, 0.02416545, 0.02412729, 
    0.02408566, 0.02404187, 0.02399619, 0.0239526, 0.02391693, 0.02387834, 
    0.02383877, 0.0237996, 0.02376081, 0.02371909, 0.02365683, 0.02359169, 
    0.02352736, 0.02348196, 0.02345889, 0.02341795, 0.02337154, 0.02332631, 
    0.02328222, 0.02323925, 0.02319736, 0.02315652, 0.0231167, 0.02306872, 
    0.02299196, 0.02292753, 0.02290579, 0.02290237, 0.02288714, 0.02286202, 
    0.02283716, 0.02281257, 0.02278824, 0.02276416, 0.02274035, 0.02271678, 
    0.02269346, 0.02267039, 0.02264756, 0.02262497, 0.02265855, 0.02263175, 
    0.02260494, 0.02257812, 0.0225513, 0.02252447, 0.02249764, 0.02247079, 
    0.02244394, 0.02241709, 0.02239022, 0.02236335, 0.02232134, 0.02225115, 
    0.02218869, 0.02219563, 0.02222345, 0.02221383, 0.02219337, 0.0221727, 
    0.02215181, 0.02213067, 0.02210928, 0.02208761, 0.02206566, 0.02204107, 
    0.02200809, 0.02194874, 0.02186848, 0.02178624, 0.02170317, 0.02162539, 
    0.02154909, 0.0214734, 0.02139835, 0.02133339, 0.02129481, 0.02126016, 
    0.02122675, 0.02119425, 0.02116277, 0.02113249, 0.02110399, 0.02107664, 
    0.02105043, 0.02103825, 0.0210416, 0.021029, 0.02101135, 0.0209943, 
    0.02097783, 0.02096191, 0.02094653, 0.02093165, 0.02091727, 0.02090504, 
    0.02090156, 0.02089821, 0.02088035, 0.02085562, 0.02084553, 0.02084445, 
    0.02084332, 0.02084214, 0.0208409, 0.02083961, 0.02083826, 0.02083687, 
    0.02083542, 0.02083393, 0.02083238, 0.02083079, 0.02128302, 0.02126604, 
    0.0212492, 0.02123248, 0.02121589, 0.02119943, 0.02118311, 0.02116692, 
    0.02115086, 0.02113494, 0.02111916, 0.02110352, 0.021073, 0.02101692, 
    0.02096648, 0.02088434, 0.02079703, 0.02074048, 0.02069322, 0.02064737, 
    0.02060298, 0.0205601, 0.02051877, 0.02047906, 0.020441, 0.02038233, 
    0.0202623, 0.02022121, 0.02025391, 0.02030596, 0.02036887, 0.02040422, 
    0.02044041, 0.02048311, 0.02053183, 0.02057018, 0.02056491, 0.02052167, 
    0.02047145, 0.02042931, 0.02039597, 0.02036922, 0.02033865, 0.02032622, 
    0.02033692, 0.02029454, 0.02018903, 0.02018268, 0.02020964, 0.02024082, 
    0.02027611, 0.02031539, 0.02035856, 0.02040549, 0.02045608, 0.02051658, 
    0.02061012, 0.02072856, 0.02089396, 0.0211239, 0.02127616, 0.02137254, 
    0.0214697, 0.02156763, 0.02166632, 0.02176577, 0.02186597, 0.0219669, 
    0.02206857, 0.02217096, 0.02227407, 0.02237788, 0.02236713, 0.02244362, 
    0.0225195, 0.02259477, 0.02266942, 0.02274345, 0.02281686, 0.02288962,
  0.02249446, 0.02252353, 0.02255239, 0.02258102, 0.02260943, 0.02263761, 
    0.02266555, 0.02269325, 0.02271961, 0.02272766, 0.02271944, 0.0226999, 
    0.02267082, 0.02264931, 0.02266161, 0.02267358, 0.02268357, 0.02269164, 
    0.02269794, 0.02270621, 0.02271526, 0.02272325, 0.02273014, 0.0227359, 
    0.02274049, 0.02274387, 0.02274601, 0.0227355, 0.02273005, 0.02274426, 
    0.02275163, 0.02275806, 0.02276359, 0.02276824, 0.02277205, 0.02277505, 
    0.02277728, 0.0227798, 0.0227836, 0.02278672, 0.02278915, 0.0227909, 
    0.02279379, 0.02283451, 0.02288858, 0.02293901, 0.02298516, 0.02302043, 
    0.02303272, 0.02304321, 0.02305359, 0.02306387, 0.02307406, 0.02308414, 
    0.02309412, 0.023104, 0.02311379, 0.02312349, 0.0231331, 0.02314261, 
    0.02315203, 0.02316136, 0.02317061, 0.02317977, 0.02325458, 0.02326852, 
    0.02328238, 0.02329616, 0.02330984, 0.02332343, 0.02333693, 0.02335034, 
    0.02336365, 0.02337687, 0.02338999, 0.02340301, 0.02341593, 0.02342875, 
    0.02344147, 0.02345407, 0.02346982, 0.02352423, 0.02358506, 0.02363979, 
    0.02368903, 0.02372519, 0.02373727, 0.02374477, 0.02374856, 0.02374877, 
    0.02374547, 0.02373362, 0.02371722, 0.02369954, 0.02368051, 0.02366008, 
    0.02363817, 0.02361473, 0.02358969, 0.0235582, 0.0235239, 0.023504, 
    0.02348503, 0.02346516, 0.02344442, 0.02342287, 0.02340055, 0.02337751, 
    0.02335378, 0.02333001, 0.0233062, 0.02328072, 0.02325348, 0.02322442, 
    0.02319147, 0.0231119, 0.02301279, 0.0229144, 0.02281731, 0.02273463, 
    0.02269854, 0.02266611, 0.02263372, 0.02260136, 0.02256904, 0.02253676, 
    0.02250452, 0.02247231, 0.02244014, 0.022408, 0.02237591, 0.02234384, 
    0.02231182, 0.02227983, 0.02224787, 0.02221595, 0.02234372, 0.02232531, 
    0.02230681, 0.02228824, 0.02226959, 0.02225085, 0.02223203, 0.02221312, 
    0.02219413, 0.02217504, 0.02215587, 0.0221366, 0.02211724, 0.02209778, 
    0.02207823, 0.02205858, 0.02204257, 0.02207112, 0.02210874, 0.02214021, 
    0.02216603, 0.02217163, 0.0221361, 0.0220986, 0.02206087, 0.02202294, 
    0.02198483, 0.02194524, 0.02190482, 0.02186438, 0.02182392, 0.02178345, 
    0.02174299, 0.02170253, 0.0216621, 0.02160871, 0.02155155, 0.02152231, 
    0.02149309, 0.02146462, 0.02143689, 0.02140986, 0.0213835, 0.0213578, 
    0.02133271, 0.02130934, 0.02128921, 0.02127096, 0.02125474, 0.02124065, 
    0.02122829, 0.02121083, 0.02119395, 0.02118263, 0.02117792, 0.02117778, 
    0.02117565, 0.02117327, 0.02117105, 0.02116896, 0.02116702, 0.02116522, 
    0.02116355, 0.02116202, 0.02116063, 0.02115936, 0.02115823, 0.02115722, 
    0.02115634, 0.02115558, 0.02115494, 0.02115442, 0.02145357, 0.02144551, 
    0.0214375, 0.02142955, 0.02142165, 0.02141382, 0.02140604, 0.02139833, 
    0.02139068, 0.02138309, 0.02137557, 0.02136811, 0.02136072, 0.0213534, 
    0.02134615, 0.02133896, 0.02132892, 0.02128437, 0.02123719, 0.02119794, 
    0.02116606, 0.02113703, 0.02110222, 0.02107099, 0.02104391, 0.02102097, 
    0.02100218, 0.02099103, 0.02098465, 0.02098086, 0.02097977, 0.02098151, 
    0.02098619, 0.02099394, 0.02100488, 0.02104109, 0.02105641, 0.02104436, 
    0.02105472, 0.02106776, 0.02108336, 0.02110144, 0.02112189, 0.02114464, 
    0.02116957, 0.02119711, 0.02122875, 0.02126458, 0.0213047, 0.02134921, 
    0.0213965, 0.02141491, 0.0214331, 0.02146836, 0.02152319, 0.02159078, 
    0.02163924, 0.02168602, 0.02173319, 0.02178074, 0.02182867, 0.02187698, 
    0.02192565, 0.02197468, 0.02202407, 0.02207381, 0.02212389, 0.02217431, 
    0.02222506, 0.02227614, 0.02232754, 0.02237925, 0.02225429, 0.02228502, 
    0.02231555, 0.02234588, 0.02237601, 0.02240594, 0.02243565, 0.02246516,
  0.02209185, 0.02210473, 0.02211759, 0.02213043, 0.02214323, 0.022156, 
    0.02216874, 0.02218144, 0.02219411, 0.02220674, 0.02221933, 0.02223188, 
    0.02224439, 0.02225686, 0.02226928, 0.02228166, 0.02229398, 0.02230626, 
    0.02231834, 0.02232417, 0.02232568, 0.02232591, 0.02232499, 0.02232302, 
    0.02232013, 0.02231642, 0.022312, 0.02230697, 0.0223114, 0.0223257, 
    0.02233989, 0.02235396, 0.02236791, 0.02238172, 0.02239539, 0.02240892, 
    0.02242232, 0.02243399, 0.02244245, 0.02245079, 0.02245908, 0.02246732, 
    0.02247551, 0.02248366, 0.02249177, 0.02249983, 0.02250785, 0.02251583, 
    0.02252378, 0.02253168, 0.02253955, 0.02254738, 0.02255518, 0.02256295, 
    0.02257068, 0.02257838, 0.02258605, 0.02259369, 0.02260131, 0.02260889, 
    0.02261645, 0.02262399, 0.0226315, 0.02263898, 0.02264009, 0.02264642, 
    0.02265265, 0.02265878, 0.02266479, 0.0226707, 0.02267649, 0.02268215, 
    0.02268768, 0.02269309, 0.02269835, 0.02270347, 0.02270844, 0.02271326, 
    0.02271792, 0.02272242, 0.02272674, 0.02273089, 0.02273486, 0.02273864, 
    0.02274222, 0.02274561, 0.02274879, 0.02275176, 0.02275451, 0.02275703, 
    0.02275959, 0.02277218, 0.02278762, 0.0227995, 0.02280808, 0.0228136, 
    0.0228163, 0.0228164, 0.02281411, 0.02280962, 0.02280872, 0.02281175, 
    0.02281369, 0.02281446, 0.02281393, 0.02281201, 0.02280856, 0.02280346, 
    0.02279659, 0.02278709, 0.02277531, 0.02276325, 0.02275095, 0.02273844, 
    0.0227257, 0.02271276, 0.0226996, 0.02268625, 0.02267271, 0.02265898, 
    0.02264507, 0.02263098, 0.02261672, 0.0226023, 0.02258772, 0.02257299, 
    0.02255811, 0.02254308, 0.02252792, 0.02251263, 0.0224972, 0.02248166, 
    0.02246599, 0.02245021, 0.02243431, 0.02241832, 0.02217826, 0.02216419, 
    0.02215012, 0.02213606, 0.02212201, 0.02210798, 0.02209395, 0.02207994, 
    0.02206594, 0.02205196, 0.02203799, 0.02202404, 0.02201011, 0.02199619, 
    0.0219823, 0.02196843, 0.02195458, 0.02194075, 0.02192696, 0.02191318, 
    0.02189944, 0.02188572, 0.02187204, 0.02185839, 0.02184477, 0.02183119, 
    0.0218177, 0.02180661, 0.02179683, 0.02178679, 0.02177651, 0.02176602, 
    0.02175534, 0.02174448, 0.02173346, 0.02172229, 0.02170967, 0.02169588, 
    0.02168329, 0.02167202, 0.02166221, 0.02165399, 0.02164753, 0.02164298, 
    0.02164052, 0.02163799, 0.02163299, 0.02162805, 0.02162323, 0.02161855, 
    0.02161399, 0.02160955, 0.02160523, 0.02160102, 0.02159693, 0.02159293, 
    0.02158904, 0.02158525, 0.02158156, 0.02157796, 0.02157444, 0.02157102, 
    0.02156767, 0.02156441, 0.02156122, 0.0215581, 0.02155506, 0.02155208, 
    0.02154917, 0.02154632, 0.02154353, 0.02154079, 0.02159664, 0.02159347, 
    0.02159035, 0.02158728, 0.02158427, 0.02158133, 0.02157844, 0.02157563, 
    0.02157288, 0.02157021, 0.02156761, 0.02156509, 0.02156266, 0.02156032, 
    0.02155806, 0.0215559, 0.02155384, 0.02155188, 0.02155003, 0.02154828, 
    0.02154665, 0.02154514, 0.02154375, 0.02154248, 0.02154135, 0.02154035, 
    0.0215393, 0.02153153, 0.02152222, 0.02151566, 0.02151168, 0.02151009, 
    0.02151073, 0.02151344, 0.02151806, 0.02152445, 0.02152488, 0.02151961, 
    0.0215163, 0.02151515, 0.02151636, 0.02152017, 0.0215268, 0.02153649, 
    0.02154949, 0.02156491, 0.02158006, 0.02159536, 0.02161084, 0.02162649, 
    0.02164232, 0.02165831, 0.02167445, 0.02169074, 0.02170718, 0.02172376, 
    0.02174048, 0.02175732, 0.02177429, 0.02179139, 0.02180859, 0.02182591, 
    0.02184333, 0.02186086, 0.02187848, 0.0218962, 0.021914, 0.02193189, 
    0.02194986, 0.0219679, 0.02198602, 0.02200421, 0.02198792, 0.02200098, 
    0.02201402, 0.02202705, 0.02204005, 0.02205303, 0.022066, 0.02207893,
  0.02197557, 0.02198026, 0.02198494, 0.02198963, 0.02199431, 0.021999, 
    0.02200369, 0.02200837, 0.02201306, 0.02201774, 0.02202243, 0.02202711, 
    0.0220318, 0.02203649, 0.02204117, 0.02204586, 0.02205054, 0.02205523, 
    0.02205991, 0.0220646, 0.02206929, 0.02207397, 0.02207866, 0.02208334, 
    0.02208803, 0.02209271, 0.0220974, 0.02210209, 0.02210677, 0.02211146, 
    0.02211614, 0.02212083, 0.02212551, 0.0221302, 0.02213489, 0.02213957, 
    0.02214426, 0.02214894, 0.02215363, 0.02215832, 0.022163, 0.02216769, 
    0.02217237, 0.02217706, 0.02218174, 0.02218643, 0.02219112, 0.0221958, 
    0.02220049, 0.02220517, 0.02220986, 0.02221454, 0.02221923, 0.02222392, 
    0.0222286, 0.02223329, 0.02223797, 0.02224266, 0.02224734, 0.02225203, 
    0.02225672, 0.0222614, 0.02226609, 0.02227077, 0.02216773, 0.0221652, 
    0.02216267, 0.02216015, 0.02215762, 0.02215509, 0.02215256, 0.02215003, 
    0.02214751, 0.02214498, 0.02214245, 0.02213992, 0.02213739, 0.02213487, 
    0.02213234, 0.02212981, 0.02212728, 0.02212475, 0.02212223, 0.0221197, 
    0.02211717, 0.02211464, 0.02211211, 0.02210958, 0.02210706, 0.02210453, 
    0.022102, 0.02209947, 0.02209694, 0.02209442, 0.02209189, 0.02208936, 
    0.02208683, 0.02208431, 0.02208178, 0.02207925, 0.02207672, 0.02207419, 
    0.02207167, 0.02206914, 0.02206661, 0.02206408, 0.02206155, 0.02205902, 
    0.0220565, 0.02205397, 0.02205144, 0.02204891, 0.02204638, 0.02204386, 
    0.02204133, 0.0220388, 0.02203627, 0.02203374, 0.02203122, 0.02202869, 
    0.02202616, 0.02202363, 0.0220211, 0.02201858, 0.02201605, 0.02201352, 
    0.02201099, 0.02200846, 0.02200593, 0.02200341, 0.02200088, 0.02199835, 
    0.02199582, 0.02199329, 0.02199077, 0.02198824, 0.02205664, 0.02205153, 
    0.02204642, 0.02204131, 0.0220362, 0.0220311, 0.02202599, 0.02202088, 
    0.02201577, 0.02201067, 0.02200556, 0.02200045, 0.02199534, 0.02199024, 
    0.02198513, 0.02198002, 0.02197491, 0.02196981, 0.0219647, 0.02195959, 
    0.02195448, 0.02194938, 0.02194427, 0.02193916, 0.02193405, 0.02192895, 
    0.02192384, 0.02191873, 0.02191362, 0.02190851, 0.02190341, 0.0218983, 
    0.02189319, 0.02188808, 0.02188298, 0.02187787, 0.02187276, 0.02186765, 
    0.02186255, 0.02185744, 0.02185233, 0.02184722, 0.02184211, 0.02183701, 
    0.0218319, 0.02182679, 0.02182169, 0.02181658, 0.02181147, 0.02180636, 
    0.02180126, 0.02179615, 0.02179104, 0.02178593, 0.02178082, 0.02177572, 
    0.02177061, 0.0217655, 0.02176039, 0.02175529, 0.02175018, 0.02174507, 
    0.02173996, 0.02173486, 0.02172975, 0.02172464, 0.02171953, 0.02171443, 
    0.02170932, 0.02170421, 0.0216991, 0.021694, 0.02171504, 0.02171799, 
    0.02172094, 0.02172389, 0.02172684, 0.02172979, 0.02173274, 0.02173569, 
    0.02173864, 0.02174159, 0.02174454, 0.02174749, 0.02175044, 0.02175339, 
    0.02175634, 0.02175929, 0.02176224, 0.02176519, 0.02176814, 0.02177108, 
    0.02177403, 0.02177699, 0.02177994, 0.02178288, 0.02178583, 0.02178879, 
    0.02179174, 0.02179468, 0.02179763, 0.02180059, 0.02180353, 0.02180648, 
    0.02180943, 0.02181238, 0.02181533, 0.02181828, 0.02182123, 0.02182418, 
    0.02182713, 0.02183008, 0.02183303, 0.02183598, 0.02183893, 0.02184188, 
    0.02184483, 0.02184778, 0.02185073, 0.02185368, 0.02185663, 0.02185958, 
    0.02186253, 0.02186548, 0.02186843, 0.02187138, 0.02187433, 0.02187728, 
    0.02188023, 0.02188318, 0.02188613, 0.02188908, 0.02189203, 0.02189498, 
    0.02189793, 0.02190088, 0.02190383, 0.02190678, 0.02190973, 0.02191268, 
    0.02191563, 0.02191858, 0.02192153, 0.02192448, 0.02193809, 0.02194277, 
    0.02194746, 0.02195214, 0.02195683, 0.02196151, 0.0219662, 0.02197088 ;

 bnds = 1, 2 ;

 lat = -89.5, -88.5, -87.5, -86.5, -85.5, -84.5, -83.5, -82.5, -81.5, -80.5, 
    -79.5, -78.5, -77.5, -76.5, -75.5, -74.5, -73.5, -72.5, -71.5, -70.5, 
    -69.5, -68.5, -67.5, -66.5, -65.5, -64.5, -63.5, -62.5, -61.5, -60.5, 
    -59.5, -58.5, -57.5, -56.5, -55.5, -54.5, -53.5, -52.5, -51.5, -50.5, 
    -49.5, -48.5, -47.5, -46.5, -45.5, -44.5, -43.5, -42.5, -41.5, -40.5, 
    -39.5, -38.5, -37.5, -36.5, -35.5, -34.5, -33.5, -32.5, -31.5, -30.5, 
    -29.5, -28.5, -27.5, -26.5, -25.5, -24.5, -23.5, -22.5, -21.5, -20.5, 
    -19.5, -18.5, -17.5, -16.5, -15.5, -14.5, -13.5, -12.5, -11.5, -10.5, 
    -9.5, -8.5, -7.5, -6.5, -5.5, -4.5, -3.5, -2.5, -1.5, -0.5, 0.5, 1.5, 
    2.5, 3.5, 4.5, 5.5, 6.5, 7.5, 8.5, 9.5, 10.5, 11.5, 12.5, 13.5, 14.5, 
    15.5, 16.5, 17.5, 18.5, 19.5, 20.5, 21.5, 22.5, 23.5, 24.5, 25.5, 26.5, 
    27.5, 28.5, 29.5, 30.5, 31.5, 32.5, 33.5, 34.5, 35.5, 36.5, 37.5, 38.5, 
    39.5, 40.5, 41.5, 42.5, 43.5, 44.5, 45.5, 46.5, 47.5, 48.5, 49.5, 50.5, 
    51.5, 52.5, 53.5, 54.5, 55.5, 56.5, 57.5, 58.5, 59.5, 60.5, 61.5, 62.5, 
    63.5, 64.5, 65.5, 66.5, 67.5, 68.5, 69.5, 70.5, 71.5, 72.5, 73.5, 74.5, 
    75.5, 76.5, 77.5, 78.5, 79.5, 80.5, 81.5, 82.5, 83.5, 84.5, 85.5, 86.5, 
    87.5, 88.5, 89.5 ;

 lat_bnds =
  -90, -89,
  -89, -88,
  -88, -87,
  -87, -86,
  -86, -85,
  -85, -84,
  -84, -83,
  -83, -82,
  -82, -81,
  -81, -80,
  -80, -79,
  -79, -78,
  -78, -77,
  -77, -76,
  -76, -75,
  -75, -74,
  -74, -73,
  -73, -72,
  -72, -71,
  -71, -70,
  -70, -69,
  -69, -68,
  -68, -67,
  -67, -66,
  -66, -65,
  -65, -64,
  -64, -63,
  -63, -62,
  -62, -61,
  -61, -60,
  -60, -59,
  -59, -58,
  -58, -57,
  -57, -56,
  -56, -55,
  -55, -54,
  -54, -53,
  -53, -52,
  -52, -51,
  -51, -50,
  -50, -49,
  -49, -48,
  -48, -47,
  -47, -46,
  -46, -45,
  -45, -44,
  -44, -43,
  -43, -42,
  -42, -41,
  -41, -40,
  -40, -39,
  -39, -38,
  -38, -37,
  -37, -36,
  -36, -35,
  -35, -34,
  -34, -33,
  -33, -32,
  -32, -31,
  -31, -30,
  -30, -29,
  -29, -28,
  -28, -27,
  -27, -26,
  -26, -25,
  -25, -24,
  -24, -23,
  -23, -22,
  -22, -21,
  -21, -20,
  -20, -19,
  -19, -18,
  -18, -17,
  -17, -16,
  -16, -15,
  -15, -14,
  -14, -13,
  -13, -12,
  -12, -11,
  -11, -10,
  -10, -9,
  -9, -8,
  -8, -7,
  -7, -6,
  -6, -5,
  -5, -4,
  -4, -3,
  -3, -2,
  -2, -1,
  -1, 0,
  0, 1,
  1, 2,
  2, 3,
  3, 4,
  4, 5,
  5, 6,
  6, 7,
  7, 8,
  8, 9,
  9, 10,
  10, 11,
  11, 12,
  12, 13,
  13, 14,
  14, 15,
  15, 16,
  16, 17,
  17, 18,
  18, 19,
  19, 20,
  20, 21,
  21, 22,
  22, 23,
  23, 24,
  24, 25,
  25, 26,
  26, 27,
  27, 28,
  28, 29,
  29, 30,
  30, 31,
  31, 32,
  32, 33,
  33, 34,
  34, 35,
  35, 36,
  36, 37,
  37, 38,
  38, 39,
  39, 40,
  40, 41,
  41, 42,
  42, 43,
  43, 44,
  44, 45,
  45, 46,
  46, 47,
  47, 48,
  48, 49,
  49, 50,
  50, 51,
  51, 52,
  52, 53,
  53, 54,
  54, 55,
  55, 56,
  56, 57,
  57, 58,
  58, 59,
  59, 60,
  60, 61,
  61, 62,
  62, 63,
  63, 64,
  64, 65,
  65, 66,
  66, 67,
  67, 68,
  68, 69,
  69, 70,
  70, 71,
  71, 72,
  72, 73,
  73, 74,
  74, 75,
  75, 76,
  76, 77,
  77, 78,
  78, 79,
  79, 80,
  80, 81,
  81, 82,
  82, 83,
  83, 84,
  84, 85,
  85, 86,
  86, 87,
  87, 88,
  88, 89,
  89, 90 ;

 lon = 0.625, 1.875, 3.125, 4.375, 5.625, 6.875, 8.125, 9.375, 10.625, 
    11.875, 13.125, 14.375, 15.625, 16.875, 18.125, 19.375, 20.625, 21.875, 
    23.125, 24.375, 25.625, 26.875, 28.125, 29.375, 30.625, 31.875, 33.125, 
    34.375, 35.625, 36.875, 38.125, 39.375, 40.625, 41.875, 43.125, 44.375, 
    45.625, 46.875, 48.125, 49.375, 50.625, 51.875, 53.125, 54.375, 55.625, 
    56.875, 58.125, 59.375, 60.625, 61.875, 63.125, 64.375, 65.625, 66.875, 
    68.125, 69.375, 70.625, 71.875, 73.125, 74.375, 75.625, 76.875, 78.125, 
    79.375, 80.625, 81.875, 83.125, 84.375, 85.625, 86.875, 88.125, 89.375, 
    90.625, 91.875, 93.125, 94.375, 95.625, 96.875, 98.125, 99.375, 100.625, 
    101.875, 103.125, 104.375, 105.625, 106.875, 108.125, 109.375, 110.625, 
    111.875, 113.125, 114.375, 115.625, 116.875, 118.125, 119.375, 120.625, 
    121.875, 123.125, 124.375, 125.625, 126.875, 128.125, 129.375, 130.625, 
    131.875, 133.125, 134.375, 135.625, 136.875, 138.125, 139.375, 140.625, 
    141.875, 143.125, 144.375, 145.625, 146.875, 148.125, 149.375, 150.625, 
    151.875, 153.125, 154.375, 155.625, 156.875, 158.125, 159.375, 160.625, 
    161.875, 163.125, 164.375, 165.625, 166.875, 168.125, 169.375, 170.625, 
    171.875, 173.125, 174.375, 175.625, 176.875, 178.125, 179.375, 180.625, 
    181.875, 183.125, 184.375, 185.625, 186.875, 188.125, 189.375, 190.625, 
    191.875, 193.125, 194.375, 195.625, 196.875, 198.125, 199.375, 200.625, 
    201.875, 203.125, 204.375, 205.625, 206.875, 208.125, 209.375, 210.625, 
    211.875, 213.125, 214.375, 215.625, 216.875, 218.125, 219.375, 220.625, 
    221.875, 223.125, 224.375, 225.625, 226.875, 228.125, 229.375, 230.625, 
    231.875, 233.125, 234.375, 235.625, 236.875, 238.125, 239.375, 240.625, 
    241.875, 243.125, 244.375, 245.625, 246.875, 248.125, 249.375, 250.625, 
    251.875, 253.125, 254.375, 255.625, 256.875, 258.125, 259.375, 260.625, 
    261.875, 263.125, 264.375, 265.625, 266.875, 268.125, 269.375, 270.625, 
    271.875, 273.125, 274.375, 275.625, 276.875, 278.125, 279.375, 280.625, 
    281.875, 283.125, 284.375, 285.625, 286.875, 288.125, 289.375, 290.625, 
    291.875, 293.125, 294.375, 295.625, 296.875, 298.125, 299.375, 300.625, 
    301.875, 303.125, 304.375, 305.625, 306.875, 308.125, 309.375, 310.625, 
    311.875, 313.125, 314.375, 315.625, 316.875, 318.125, 319.375, 320.625, 
    321.875, 323.125, 324.375, 325.625, 326.875, 328.125, 329.375, 330.625, 
    331.875, 333.125, 334.375, 335.625, 336.875, 338.125, 339.375, 340.625, 
    341.875, 343.125, 344.375, 345.625, 346.875, 348.125, 349.375, 350.625, 
    351.875, 353.125, 354.375, 355.625, 356.875, 358.125, 359.375 ;

 lon_bnds =
  0, 1.25,
  1.25, 2.5,
  2.5, 3.75,
  3.75, 5,
  5, 6.25,
  6.25, 7.5,
  7.5, 8.75,
  8.75, 10,
  10, 11.25,
  11.25, 12.5,
  12.5, 13.75,
  13.75, 15,
  15, 16.25,
  16.25, 17.5,
  17.5, 18.75,
  18.75, 20,
  20, 21.25,
  21.25, 22.5,
  22.5, 23.75,
  23.75, 25,
  25, 26.25,
  26.25, 27.5,
  27.5, 28.75,
  28.75, 30,
  30, 31.25,
  31.25, 32.5,
  32.5, 33.75,
  33.75, 35,
  35, 36.25,
  36.25, 37.5,
  37.5, 38.75,
  38.75, 40,
  40, 41.25,
  41.25, 42.5,
  42.5, 43.75,
  43.75, 45,
  45, 46.25,
  46.25, 47.5,
  47.5, 48.75,
  48.75, 50,
  50, 51.25,
  51.25, 52.5,
  52.5, 53.75,
  53.75, 55,
  55, 56.25,
  56.25, 57.5,
  57.5, 58.75,
  58.75, 60,
  60, 61.25,
  61.25, 62.5,
  62.5, 63.75,
  63.75, 65,
  65, 66.25,
  66.25, 67.5,
  67.5, 68.75,
  68.75, 70,
  70, 71.25,
  71.25, 72.5,
  72.5, 73.75,
  73.75, 75,
  75, 76.25,
  76.25, 77.5,
  77.5, 78.75,
  78.75, 80,
  80, 81.25,
  81.25, 82.5,
  82.5, 83.75,
  83.75, 85,
  85, 86.25,
  86.25, 87.5,
  87.5, 88.75,
  88.75, 90,
  90, 91.25,
  91.25, 92.5,
  92.5, 93.75,
  93.75, 95,
  95, 96.25,
  96.25, 97.5,
  97.5, 98.75,
  98.75, 100,
  100, 101.25,
  101.25, 102.5,
  102.5, 103.75,
  103.75, 105,
  105, 106.25,
  106.25, 107.5,
  107.5, 108.75,
  108.75, 110,
  110, 111.25,
  111.25, 112.5,
  112.5, 113.75,
  113.75, 115,
  115, 116.25,
  116.25, 117.5,
  117.5, 118.75,
  118.75, 120,
  120, 121.25,
  121.25, 122.5,
  122.5, 123.75,
  123.75, 125,
  125, 126.25,
  126.25, 127.5,
  127.5, 128.75,
  128.75, 130,
  130, 131.25,
  131.25, 132.5,
  132.5, 133.75,
  133.75, 135,
  135, 136.25,
  136.25, 137.5,
  137.5, 138.75,
  138.75, 140,
  140, 141.25,
  141.25, 142.5,
  142.5, 143.75,
  143.75, 145,
  145, 146.25,
  146.25, 147.5,
  147.5, 148.75,
  148.75, 150,
  150, 151.25,
  151.25, 152.5,
  152.5, 153.75,
  153.75, 155,
  155, 156.25,
  156.25, 157.5,
  157.5, 158.75,
  158.75, 160,
  160, 161.25,
  161.25, 162.5,
  162.5, 163.75,
  163.75, 165,
  165, 166.25,
  166.25, 167.5,
  167.5, 168.75,
  168.75, 170,
  170, 171.25,
  171.25, 172.5,
  172.5, 173.75,
  173.75, 175,
  175, 176.25,
  176.25, 177.5,
  177.5, 178.75,
  178.75, 180,
  180, 181.25,
  181.25, 182.5,
  182.5, 183.75,
  183.75, 185,
  185, 186.25,
  186.25, 187.5,
  187.5, 188.75,
  188.75, 190,
  190, 191.25,
  191.25, 192.5,
  192.5, 193.75,
  193.75, 195,
  195, 196.25,
  196.25, 197.5,
  197.5, 198.75,
  198.75, 200,
  200, 201.25,
  201.25, 202.5,
  202.5, 203.75,
  203.75, 205,
  205, 206.25,
  206.25, 207.5,
  207.5, 208.75,
  208.75, 210,
  210, 211.25,
  211.25, 212.5,
  212.5, 213.75,
  213.75, 215,
  215, 216.25,
  216.25, 217.5,
  217.5, 218.75,
  218.75, 220,
  220, 221.25,
  221.25, 222.5,
  222.5, 223.75,
  223.75, 225,
  225, 226.25,
  226.25, 227.5,
  227.5, 228.75,
  228.75, 230,
  230, 231.25,
  231.25, 232.5,
  232.5, 233.75,
  233.75, 235,
  235, 236.25,
  236.25, 237.5,
  237.5, 238.75,
  238.75, 240,
  240, 241.25,
  241.25, 242.5,
  242.5, 243.75,
  243.75, 245,
  245, 246.25,
  246.25, 247.5,
  247.5, 248.75,
  248.75, 250,
  250, 251.25,
  251.25, 252.5,
  252.5, 253.75,
  253.75, 255,
  255, 256.25,
  256.25, 257.5,
  257.5, 258.75,
  258.75, 260,
  260, 261.25,
  261.25, 262.5,
  262.5, 263.75,
  263.75, 265,
  265, 266.25,
  266.25, 267.5,
  267.5, 268.75,
  268.75, 270,
  270, 271.25,
  271.25, 272.5,
  272.5, 273.75,
  273.75, 275,
  275, 276.25,
  276.25, 277.5,
  277.5, 278.75,
  278.75, 280,
  280, 281.25,
  281.25, 282.5,
  282.5, 283.75,
  283.75, 285,
  285, 286.25,
  286.25, 287.5,
  287.5, 288.75,
  288.75, 290,
  290, 291.25,
  291.25, 292.5,
  292.5, 293.75,
  293.75, 295,
  295, 296.25,
  296.25, 297.5,
  297.5, 298.75,
  298.75, 300,
  300, 301.25,
  301.25, 302.5,
  302.5, 303.75,
  303.75, 305,
  305, 306.25,
  306.25, 307.5,
  307.5, 308.75,
  308.75, 310,
  310, 311.25,
  311.25, 312.5,
  312.5, 313.75,
  313.75, 315,
  315, 316.25,
  316.25, 317.5,
  317.5, 318.75,
  318.75, 320,
  320, 321.25,
  321.25, 322.5,
  322.5, 323.75,
  323.75, 325,
  325, 326.25,
  326.25, 327.5,
  327.5, 328.75,
  328.75, 330,
  330, 331.25,
  331.25, 332.5,
  332.5, 333.75,
  333.75, 335,
  335, 336.25,
  336.25, 337.5,
  337.5, 338.75,
  338.75, 340,
  340, 341.25,
  341.25, 342.5,
  342.5, 343.75,
  343.75, 345,
  345, 346.25,
  346.25, 347.5,
  347.5, 348.75,
  348.75, 350,
  350, 351.25,
  351.25, 352.5,
  352.5, 353.75,
  353.75, 355,
  355, 356.25,
  356.25, 357.5,
  357.5, 358.75,
  358.75, 360 ;

 time = 913 ;

 time_bnds =
  0, 1826 ;

 average_T1 = 0 ;

 average_T2 = 1826 ;

 average_DT = 1826 ;
}
