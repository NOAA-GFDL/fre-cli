netcdf \00010101.atmos_daily.tile1.temp {
dimensions:
	time = UNLIMITED ; // (181 currently)
	phalf = 66 ;
	grid_xt = 15 ;
	grid_yt = 10 ;
	scalar_axis = 1 ;
	nv = 2 ;
	pfull = 1 ;
variables:
	double average_DT(time) ;
		average_DT:_FillValue = 1.e+20 ;
		average_DT:missing_value = 1.e+20 ;
		average_DT:units = "days" ;
		average_DT:long_name = "Length of average period" ;
	double average_T1(time) ;
		average_T1:_FillValue = 1.e+20 ;
		average_T1:missing_value = 1.e+20 ;
		average_T1:units = "days since 0001-01-01 00:00:00" ;
		average_T1:long_name = "Start time for average period" ;
	double average_T2(time) ;
		average_T2:_FillValue = 1.e+20 ;
		average_T2:missing_value = 1.e+20 ;
		average_T2:units = "days since 0001-01-01 00:00:00" ;
		average_T2:long_name = "End time for average period" ;
	float bk(phalf) ;
		bk:_FillValue = 1.e+20f ;
		bk:missing_value = 1.e+20f ;
		bk:long_name = "vertical coordinate sigma value" ;
		bk:cell_methods = "time: point" ;
	double grid_xt(grid_xt) ;
		grid_xt:units = "degrees_E" ;
		grid_xt:long_name = "T-cell longitude" ;
		grid_xt:axis = "X" ;
	double grid_yt(grid_yt) ;
		grid_yt:units = "degrees_N" ;
		grid_yt:long_name = "T-cell latitude" ;
		grid_yt:axis = "Y" ;
	float height10m(scalar_axis) ;
		height10m:_FillValue = 1.e+20f ;
		height10m:missing_value = 1.e+20f ;
		height10m:units = "m" ;
		height10m:long_name = "Height" ;
		height10m:cell_methods = "time: point" ;
		height10m:axis = "Z" ;
		height10m:positive = "up" ;
		height10m:standard_name = "height" ;
	float height2m(scalar_axis) ;
		height2m:_FillValue = 1.e+20f ;
		height2m:missing_value = 1.e+20f ;
		height2m:units = "m" ;
		height2m:long_name = "Height" ;
		height2m:cell_methods = "time: point" ;
		height2m:axis = "Z" ;
		height2m:positive = "up" ;
		height2m:standard_name = "height" ;
	float land_mask(grid_yt, grid_xt) ;
		land_mask:_FillValue = 1.e+20f ;
		land_mask:missing_value = 1.e+20f ;
		land_mask:valid_range = -0.01f, 1.01f ;
		land_mask:long_name = "fractional amount of land" ;
		land_mask:cell_methods = "time: point" ;
		land_mask:interp_method = "conserve_order1" ;
	double nv(nv) ;
		nv:long_name = "vertex number" ;
	double pfull(pfull) ;
		pfull:units = "mb" ;
		pfull:long_name = "ref full pressure level" ;
		pfull:axis = "Z" ;
		pfull:positive = "down" ;
	double phalf(phalf) ;
		phalf:units = "mb" ;
		phalf:long_name = "ref half pressure level" ;
		phalf:axis = "Z" ;
		phalf:positive = "down" ;
	float pk(phalf) ;
		pk:_FillValue = 1.e+20f ;
		pk:missing_value = 1.e+20f ;
		pk:units = "pascal" ;
		pk:long_name = "pressure part of the hybrid coordinate" ;
		pk:cell_methods = "time: point" ;
	double scalar_axis(scalar_axis) ;
		scalar_axis:long_name = "none" ;
	float sftlf(grid_yt, grid_xt) ;
		sftlf:_FillValue = 1.e+20f ;
		sftlf:missing_value = 1.e+20f ;
		sftlf:units = "1.0" ;
		sftlf:long_name = "Fraction of the Grid Cell Occupied by Land" ;
		sftlf:cell_methods = "time: point" ;
		sftlf:cell_measures = "area: area" ;
		sftlf:standard_name = "land_area_fraction" ;
		sftlf:interp_method = "conserve_order1" ;
	float temp(time, pfull, grid_yt, grid_xt) ;
		temp:_FillValue = -1.e+10f ;
		temp:missing_value = -1.e+10f ;
		temp:valid_range = 100.f, 350.f ;
		temp:units = "K" ;
		temp:long_name = "temperature" ;
		temp:cell_methods = "time: mean" ;
		temp:time_avg_info = "average_T1,average_T2,average_DT" ;
	double time(time) ;
		time:units = "days since 0001-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "NOLEAP" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bnds" ;
	double time_bnds(time, nv) ;
		time_bnds:long_name = "time axis boundaries" ;
	float zsurf(grid_yt, grid_xt) ;
		zsurf:_FillValue = 1.e+20f ;
		zsurf:missing_value = 1.e+20f ;
		zsurf:units = "m" ;
		zsurf:long_name = "surface height" ;
		zsurf:cell_methods = "time: point" ;
		zsurf:interp_method = "conserve_order1" ;

// global attributes:
		:title = "cm5_c96_am5f7c1r0_b06_piC_galb_noiceinit_alb" ;
		:associated_files = "area: 00010101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:history = "Mon Feb  2 22:06:42 2026: ncks -d time,0,180 old/00010101.atmos_daily.tile1.temp.nc 00010101.atmos_daily.tile1.temp.nc\nMon Feb  2 15:24:42 2026: ncks -d pfull,0,0 out.nc 00010101.atmos_daily.tile1.temp.nc\nFri Aug 29 13:34:10 2025: ncks -d grid_xt,0,14 -d grid_yt,0,9 -d time,0,181 /work/cew/scratch//00010101.atmos_daily.tile1.nc -O /work/cew/scratch/workflow-test/atmos_daily//ncks_out//00010101.atmos_daily.tile1.nc" ;
		:NCO = "netCDF Operators version 5.2.4 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 average_DT = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 average_T1 = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 
    18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 
    36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 
    54, 55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 
    72, 73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 
    90, 91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 
    106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 
    120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 
    134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 
    148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 
    162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 
    176, 177, 178, 179, 180 ;

 average_T2 = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 
    19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 
    37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 
    55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 
    73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 
    91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 106, 
    107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 
    121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 
    135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 
    149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 
    163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 
    177, 178, 179, 180, 181 ;

 bk = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.00193294, 0.00749994, 0.01640714, 0.02841953, 
    0.04334756, 0.06103661, 0.0813586, 0.1042054, 0.1294836, 0.1571101, 
    0.1870091, 0.2191095, 0.2533426, 0.2896406, 0.3279357, 0.3681587, 
    0.4102391, 0.454293, 0.5001689, 0.5468886, 0.5935643, 0.6397641, 
    0.6851825, 0.729505, 0.7723162, 0.8125153, 0.8492141, 0.8817441, 
    0.909788, 0.9332725, 0.9524949, 0.9678352, 0.9798011, 0.9889621, 0.99575, 1 ;

 grid_xt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15 ;

 grid_yt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10 ;

 height10m = 10 ;

 height2m = 2 ;

 land_mask =
  0.1986115, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.9611561, 0.1583273, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 0.7949425, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 0.7552791, 0.2484612, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 0.9872221, 0.4156101, 0.04560489, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 0.8345782, 0.2958934, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 0.7792858, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 0.9990003, 0.3505592, 0.06537855, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 0.8140894, 0.2409153, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 0.9453563, 0.02902743, 0, 0, 0, 0, 0, 0, 0, 0 ;

 nv = 1, 2 ;

 pfull = 0.0252729048206747 ;

 phalf = 0.01, 0.0513470268, 0.1404240036, 0.3072783852, 0.5379505539, 
    0.8245489502, 1.170559845, 1.5862843323, 2.0879000854, 2.700272522, 
    3.4550848389, 4.3841940308, 5.5185266113, 6.8925054932, 8.5440936279, 
    10.5147802734, 12.8495031738, 15.5965148926, 18.8071691895, 
    22.5356542969, 26.8386547852, 31.7749560547, 37.4049951172, 
    43.7903613281, 50.9932617188, 59.0759326172, 68.100078125, 78.1262353516, 
    89.2131933594, 101.4173632812, 114.7922466406, 129.3878501562, 
    145.2501478125, 162.4206823438, 180.9360560938, 200.8276451562, 
    222.1212074219, 244.8367185938, 268.9881007812, 294.5831945312, 
    321.6236510156, 350.1049399219, 380.0163883594, 411.3414303125, 
    444.0575547656, 478.1367280469, 513.5456339062, 550.403556875, 
    588.6019571094, 627.3470909766, 665.9273852344, 704.0097012891, 
    741.2475327734, 777.2856108203, 811.7659041211, 843.9830114648, 
    873.3803854492, 899.5263707422, 922.2501762402, 941.5376650684, 
    957.6070185254, 970.7426572876, 981.30107, 989.65107, 995.9000099865, 1000 ;

 pk = 1, 5.134703, 14.0424, 30.72784, 53.79506, 82.4549, 117.056, 158.6284, 
    208.79, 270.0273, 345.5085, 438.4194, 551.8527, 689.2505, 854.4094, 
    1051.478, 1284.95, 1559.651, 1880.717, 2253.565, 2683.865, 3177.496, 
    3740.5, 4379.036, 5099.326, 5907.593, 6810.008, 7812.624, 8921.319, 
    10141.74, 11285.93, 12188.79, 12884.3, 13400.12, 13758.85, 13979.1, 
    14076.26, 14063.13, 13950.46, 13747.31, 13461.45, 13099.54, 12667.38, 
    12170.08, 11612.19, 10997.8, 10330.65, 9611.055, 8843.304, 8045.85, 
    7236.312, 6424.557, 5606.509, 4778.059, 3944.972, 3146.775, 2416.634, 
    1778.226, 1246.215, 826.5195, 511.2139, 290.7407, 150, 68.893, 14.999, 0 ;

 scalar_axis = 0 ;

 sftlf =
  0.1986115, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.9611561, 0.1583273, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 0.7949425, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 0.7552791, 0.2484612, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 0.9872221, 0.4156101, 0.04560489, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 0.8345782, 0.2958934, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 0.7792858, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 0.9990003, 0.3505592, 0.06537855, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 0.8140894, 0.2409153, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 0.9453563, 0.02902743, 0, 0, 0, 0, 0, 0, 0, 0 ;

 temp =
  208.4635, 208.4194, 208.3678, 208.3111, 208.28, 208.2588, 208.264, 
    208.2572, 208.2392, 208.1897, 208.1172, 208.0198, 207.9185, 207.8336, 
    207.7737,
  208.699, 208.6725, 208.6208, 208.5544, 208.5045, 208.4645, 208.4583, 
    208.4631, 208.4673, 208.4495, 208.407, 208.3336, 208.2427, 208.1455, 
    208.0561,
  208.6891, 208.701, 208.6814, 208.6083, 208.551, 208.5075, 208.501, 
    208.5308, 208.5639, 208.5924, 208.5999, 208.5672, 208.4985, 208.3997, 
    208.2924,
  208.8424, 208.8699, 208.8607, 208.821, 208.751, 208.6781, 208.6407, 
    208.6486, 208.6992, 208.7618, 208.8182, 208.8369, 208.8115, 208.7351, 
    208.627,
  208.8215, 208.8781, 208.8903, 208.8715, 208.8365, 208.7707, 208.7203, 
    208.703, 208.7376, 208.8129, 208.9003, 208.9746, 209.0067, 208.9809, 
    208.9066,
  208.8997, 208.9688, 209.0045, 208.993, 208.9657, 208.9237, 208.8728, 
    208.8393, 208.8501, 208.9094, 209.0145, 209.1328, 209.2153, 209.2505, 
    209.2187,
  208.8504, 208.9283, 208.9876, 209.0336, 209.0429, 208.9932, 208.9529, 
    208.9049, 208.9107, 208.9427, 209.0481, 209.1828, 209.3256, 209.426, 
    209.4653,
  208.8611, 208.9474, 209.0175, 209.0806, 209.1368, 209.1075, 209.0728, 
    209.0204, 208.9922, 209.0213, 209.0934, 209.244, 209.4078, 209.5706, 
    209.6783,
  208.772, 208.8943, 209.0072, 209.0595, 209.152, 209.1864, 209.1552, 
    209.0986, 209.0592, 209.0484, 209.1186, 209.235, 209.4199, 209.612, 
    209.787,
  208.7096, 208.8593, 208.994, 209.1085, 209.2084, 209.2517, 209.2431, 
    209.2048, 209.1703, 209.1381, 209.1587, 209.2627, 209.4147, 209.6303, 
    209.8408,
  210.3387, 210.2716, 210.2551, 210.219, 210.1703, 210.0922, 210.0163, 
    209.9483, 209.8922, 209.8327, 209.7596, 209.6541, 209.5165, 209.3435, 
    209.1556,
  210.6138, 210.5299, 210.4781, 210.4366, 210.3918, 210.3309, 210.2633, 
    210.1938, 210.1306, 210.0651, 209.9879, 209.8764, 209.7409, 209.566, 
    209.3711,
  210.6581, 210.5719, 210.5103, 210.4483, 210.3933, 210.3411, 210.2886, 
    210.2342, 210.1889, 210.1375, 210.0773, 209.9827, 209.8632, 209.7054, 
    209.5192,
  210.8645, 210.77, 210.6887, 210.6206, 210.5595, 210.4913, 210.4356, 
    210.3771, 210.3315, 210.2885, 210.2409, 210.1656, 210.0571, 209.9122, 
    209.7341,
  210.9275, 210.8231, 210.7315, 210.6516, 210.5894, 210.5201, 210.4562, 
    210.3979, 210.3505, 210.3177, 210.2848, 210.237, 210.1614, 210.0415, 
    209.8806,
  211.065, 210.963, 210.8639, 210.7596, 210.6866, 210.6187, 210.5585, 
    210.496, 210.4385, 210.3956, 210.3629, 210.3344, 210.2889, 210.2017, 
    210.0704,
  211.0497, 210.9716, 210.8811, 210.8, 210.7147, 210.6364, 210.5731, 
    210.5197, 210.4626, 210.4099, 210.3727, 210.3443, 210.3263, 210.2766, 
    210.1928,
  211.0808, 211.0289, 210.9578, 210.8885, 210.8079, 210.7257, 210.6614, 
    210.5963, 210.5385, 210.4776, 210.4256, 210.3834, 210.3673, 210.345, 
    210.2994,
  211.0717, 211.0325, 210.9725, 210.8933, 210.8375, 210.7834, 210.7131, 
    210.6452, 210.5784, 210.5035, 210.4426, 210.3788, 210.3499, 210.3386, 
    210.325,
  211.1274, 211.0866, 211.0245, 210.9595, 210.8959, 210.8228, 210.7683, 
    210.7124, 210.6519, 210.5654, 210.4829, 210.3979, 210.3417, 210.3151, 
    210.3175,
  209.2334, 209.2643, 209.3478, 209.3565, 209.3357, 209.2693, 209.1786, 
    209.0705, 208.9595, 208.8492, 208.7626, 208.6944, 208.6524, 208.6291, 
    208.6359,
  209.3273, 209.3876, 209.4408, 209.4659, 209.4819, 209.4682, 209.4281, 
    209.3452, 209.2409, 209.1227, 209.0121, 208.9186, 208.8516, 208.8139, 
    208.8042,
  209.2857, 209.3968, 209.463, 209.4993, 209.5262, 209.5401, 209.5333, 
    209.4948, 209.4251, 209.3203, 209.2, 209.087, 209.0032, 208.9431, 208.9192,
  209.3386, 209.454, 209.5648, 209.6345, 209.6807, 209.692, 209.7078, 
    209.6983, 209.6713, 209.5995, 209.5002, 209.3827, 209.2731, 209.1807, 
    209.1249,
  209.2589, 209.3417, 209.4648, 209.5771, 209.6677, 209.7094, 209.7349, 
    209.7425, 209.7455, 209.7277, 209.6803, 209.5963, 209.4924, 209.3923, 
    209.3116,
  209.4225, 209.4425, 209.4912, 209.5631, 209.6527, 209.7298, 209.7929, 
    209.837, 209.868, 209.8787, 209.8687, 209.8299, 209.7529, 209.6608, 
    209.5737,
  209.4768, 209.4988, 209.5137, 209.5437, 209.5977, 209.6484, 209.7319, 
    209.8238, 209.9054, 209.9554, 209.9729, 209.9666, 209.9233, 209.8484, 
    209.7658,
  209.4787, 209.556, 209.602, 209.6234, 209.6472, 209.6743, 209.7351, 
    209.836, 209.965, 210.0627, 210.1226, 210.1378, 210.1189, 210.0613, 
    209.9823,
  209.4438, 209.5791, 209.6246, 209.635, 209.6669, 209.7046, 209.7327, 
    209.8046, 209.9352, 210.0782, 210.1939, 210.2431, 210.2462, 210.2133, 
    210.1485,
  209.4542, 209.593, 209.6911, 209.7229, 209.7486, 209.7693, 209.7792, 
    209.8319, 209.9558, 210.0935, 210.2385, 210.3335, 210.3679, 210.3575, 
    210.3074,
  210.9213, 210.859, 210.8355, 210.7602, 210.6738, 210.5651, 210.4466, 
    210.3198, 210.2033, 210.095, 209.9914, 209.8901, 209.796, 209.7071, 
    209.6258,
  211.1872, 211.1087, 211.0563, 210.9938, 210.9222, 210.8233, 210.7106, 
    210.5818, 210.4538, 210.3284, 210.2117, 210.1045, 210.0048, 209.9146, 
    209.8248,
  211.2531, 211.1672, 211.1154, 211.0448, 210.9691, 210.8692, 210.765, 
    210.6485, 210.5298, 210.4172, 210.3083, 210.2096, 210.1116, 210.0217, 
    209.9365,
  211.4785, 211.3703, 211.2996, 211.2195, 211.1433, 211.0555, 210.9549, 
    210.8456, 210.7253, 210.6138, 210.5078, 210.4121, 210.3209, 210.2314, 
    210.1466,
  211.5859, 211.4545, 211.3586, 211.2612, 211.1849, 211.1098, 211.0163, 
    210.9076, 210.7939, 210.6818, 210.5815, 210.4933, 210.4193, 210.3438, 
    210.2716,
  211.7933, 211.6594, 211.5499, 211.4258, 211.3338, 211.2618, 211.1806, 
    211.0706, 210.9532, 210.8373, 210.7344, 210.6481, 210.5754, 210.5078, 
    210.4388,
  211.9003, 211.7482, 211.6252, 211.5279, 211.4478, 211.3476, 211.258, 
    211.1374, 211.0101, 210.8903, 210.7808, 210.6897, 210.6175, 210.5623, 
    210.5154,
  212.0213, 211.872, 211.7442, 211.6545, 211.5851, 211.4981, 211.3987, 
    211.2687, 211.1344, 211.0025, 210.8754, 210.765, 210.6779, 210.6222, 
    210.6016,
  212.0626, 211.9273, 211.8, 211.6734, 211.6053, 211.5648, 211.4707, 
    211.3589, 211.226, 211.0789, 210.9466, 210.8249, 210.7282, 210.6622, 
    210.6319,
  212.1459, 212.0105, 211.8991, 211.7841, 211.6953, 211.6282, 211.53, 
    211.4314, 211.328, 211.1697, 211.0422, 210.9156, 210.8035, 210.7172, 
    210.6653,
  212.3093, 212.1735, 212.0835, 211.9536, 211.8651, 211.7985, 211.772, 
    211.771, 211.7763, 211.7628, 211.7355, 211.7013, 211.6405, 211.5729, 
    211.5036,
  212.6312, 212.5063, 212.4404, 212.3194, 212.2255, 212.1386, 212.0923, 
    212.0453, 212.0303, 212.0125, 211.9938, 211.9688, 211.9259, 211.8746, 
    211.8127,
  212.7264, 212.6378, 212.6028, 212.4939, 212.4091, 212.3202, 212.2645, 
    212.2069, 212.1763, 212.1527, 212.1351, 212.1183, 212.0945, 212.0696, 
    212.0309,
  212.946, 212.8671, 212.8459, 212.7616, 212.679, 212.5936, 212.5247, 
    212.4554, 212.4058, 212.3719, 212.3538, 212.3326, 212.3082, 212.2842, 
    212.2562,
  212.996, 212.9677, 212.9784, 212.9289, 212.8763, 212.806, 212.7372, 
    212.6603, 212.5931, 212.5407, 212.5107, 212.4836, 212.4593, 212.4379, 
    212.4168,
  213.1053, 213.107, 213.1488, 213.1203, 213.1067, 213.0634, 213.018, 
    212.945, 212.8719, 212.7939, 212.7369, 212.695, 212.6588, 212.6277, 
    212.6028,
  213.0659, 213.0885, 213.1577, 213.1864, 213.2246, 213.2177, 213.2, 
    213.1573, 213.0993, 213.0239, 212.9447, 212.8823, 212.8343, 212.795, 
    212.7636,
  213.0429, 213.0922, 213.1737, 213.2389, 213.323, 213.35, 213.3692, 
    213.3588, 213.3377, 213.2833, 213.1909, 213.1025, 213.034, 212.9758, 
    212.9354,
  212.9544, 213.0284, 213.1182, 213.1857, 213.3115, 213.4024, 213.4544, 
    213.4755, 213.4911, 213.471, 213.4136, 213.3258, 213.2452, 213.1703, 
    213.1088,
  212.9197, 213.0011, 213.1106, 213.2001, 213.3172, 213.4247, 213.5065, 
    213.5581, 213.6088, 213.6059, 213.5865, 213.5304, 213.4654, 213.3895, 
    213.3246,
  212.0979, 212.0076, 211.8932, 211.7525, 211.582, 211.3712, 211.1428, 
    210.9015, 210.6733, 210.4684, 210.3009, 210.1761, 210.0865, 210.0145, 
    209.9425,
  212.18, 212.1273, 212.0339, 211.945, 211.8348, 211.6757, 211.4699, 
    211.2278, 210.9928, 210.7699, 210.5659, 210.3885, 210.2483, 210.1432, 
    210.0638,
  212.0371, 212.0433, 212.0021, 211.9489, 211.8593, 211.7478, 211.5898, 
    211.3971, 211.1844, 210.9593, 210.7393, 210.5308, 210.3502, 210.2069, 
    210.1016,
  212.1275, 212.103, 212.0572, 211.9879, 211.9181, 211.8267, 211.7203, 
    211.5658, 211.3831, 211.1927, 210.9839, 210.7626, 210.5531, 210.3676, 
    210.2316,
  212.1016, 212.0301, 211.9662, 211.9058, 211.8497, 211.7901, 211.6958, 
    211.568, 211.4315, 211.2858, 211.1013, 210.8947, 210.6797, 210.492, 
    210.3459,
  212.0651, 212.0181, 211.9783, 211.9301, 211.86, 211.7959, 211.7199, 
    211.6369, 211.5406, 211.4057, 211.2455, 211.0619, 210.8507, 210.6597, 
    210.5007,
  211.9791, 211.921, 211.8839, 211.8601, 211.8243, 211.7607, 211.683, 
    211.5999, 211.5172, 211.4132, 211.2928, 211.1362, 210.952, 210.7656, 
    210.6066,
  211.9299, 211.8723, 211.8261, 211.8084, 211.784, 211.7322, 211.6434, 
    211.5562, 211.4933, 211.4316, 211.3445, 211.2171, 211.0603, 210.8914, 
    210.731,
  211.8299, 211.8163, 211.7788, 211.7262, 211.7016, 211.6544, 211.5751, 
    211.509, 211.45, 211.3896, 211.3201, 211.219, 211.0928, 210.947, 210.8014,
  211.7502, 211.754, 211.7132, 211.6682, 211.6211, 211.5747, 211.5095, 
    211.4513, 211.4171, 211.3451, 211.2875, 211.2001, 211.0985, 210.977, 
    210.8532,
  210.9064, 210.9189, 210.9865, 211.0451, 211.1293, 211.2006, 211.2691, 
    211.3049, 211.3097, 211.2754, 211.2103, 211.1193, 211.0196, 210.9343, 
    210.8715,
  211.1564, 211.1147, 211.152, 211.181, 211.243, 211.3024, 211.3712, 
    211.4226, 211.4556, 211.4471, 211.405, 211.3315, 211.2438, 211.1616, 
    211.0983,
  211.2504, 211.2071, 211.2161, 211.205, 211.2217, 211.2521, 211.306, 
    211.3616, 211.4235, 211.4643, 211.4801, 211.4584, 211.4014, 211.3254, 
    211.2511,
  211.4201, 211.3714, 211.352, 211.301, 211.2799, 211.2705, 211.2887, 
    211.3243, 211.3962, 211.4625, 211.5295, 211.5562, 211.5387, 211.4796, 
    211.3988,
  211.4861, 211.4136, 211.3879, 211.335, 211.3062, 211.2814, 211.2865, 
    211.3084, 211.3739, 211.4437, 211.5251, 211.5913, 211.6206, 211.6009, 
    211.54,
  211.5885, 211.5203, 211.4949, 211.4366, 211.4101, 211.3888, 211.3854, 
    211.3895, 211.4207, 211.4809, 211.5629, 211.6587, 211.716, 211.7233, 
    211.6814,
  211.6665, 211.612, 211.5857, 211.5653, 211.5576, 211.5163, 211.4859, 
    211.4585, 211.462, 211.5047, 211.5682, 211.6534, 211.7361, 211.7773, 
    211.7709,
  211.7643, 211.7247, 211.718, 211.7279, 211.74, 211.6979, 211.655, 211.6043, 
    211.5759, 211.5743, 211.6133, 211.678, 211.7601, 211.8271, 211.8483,
  211.8103, 211.8257, 211.8475, 211.8524, 211.8662, 211.8345, 211.7939, 
    211.7527, 211.7057, 211.6509, 211.6532, 211.692, 211.7681, 211.8432, 
    211.8986,
  211.894, 211.9066, 211.9562, 211.995, 212.0072, 211.9712, 211.9448, 
    211.9188, 211.892, 211.792, 211.7489, 211.7622, 211.8209, 211.9078, 
    211.9746,
  210.3648, 210.2375, 210.1955, 210.1771, 210.2043, 210.2341, 210.2789, 
    210.2906, 210.2775, 210.227, 210.15, 210.0561, 209.953, 209.8483, 209.7467,
  210.5881, 210.45, 210.367, 210.3386, 210.3506, 210.3834, 210.4323, 
    210.4705, 210.4843, 210.4666, 210.413, 210.3324, 210.2295, 210.1203, 
    210.0107,
  210.6279, 210.5223, 210.4194, 210.3519, 210.3522, 210.3804, 210.4326, 
    210.4929, 210.5338, 210.5503, 210.5338, 210.4833, 210.4098, 210.3114, 
    210.2099,
  210.7943, 210.6942, 210.5748, 210.4816, 210.444, 210.4586, 210.5012, 
    210.5646, 210.6246, 210.6661, 210.678, 210.6552, 210.597, 210.5124, 
    210.4117,
  210.8717, 210.7707, 210.6466, 210.5426, 210.4693, 210.4484, 210.4799, 
    210.5378, 210.6097, 210.6717, 210.7079, 210.7133, 210.6896, 210.6341, 
    210.5586,
  210.9695, 210.8698, 210.7453, 210.6293, 210.5415, 210.4929, 210.5112, 
    210.5566, 210.6359, 210.7077, 210.7688, 210.8013, 210.8031, 210.7742, 
    210.7121,
  211.0158, 210.9209, 210.8089, 210.7003, 210.6105, 210.5283, 210.5065, 
    210.5348, 210.6044, 210.6845, 210.7539, 210.8078, 210.8332, 210.8375, 
    210.8116,
  211.0358, 210.9627, 210.8731, 210.7771, 210.6907, 210.6117, 210.5702, 
    210.5665, 210.6205, 210.6867, 210.7677, 210.8358, 210.8882, 210.9214, 
    210.9221,
  211.0132, 210.9673, 210.8791, 210.7808, 210.7001, 210.6241, 210.575, 
    210.5603, 210.595, 210.645, 210.723, 210.8023, 210.861, 210.9062, 210.9178,
  210.9867, 210.945, 210.8996, 210.849, 210.7651, 210.6736, 210.6053, 
    210.5856, 210.6041, 210.6284, 210.6846, 210.7585, 210.8221, 210.8773, 
    210.9095,
  212.2787, 212.1641, 212.0433, 211.8848, 211.7186, 211.5289, 211.3448, 
    211.1592, 210.9974, 210.8677, 210.779, 210.7397, 210.7507, 210.8119, 
    210.9074,
  212.5175, 212.4081, 212.2878, 212.1297, 211.9636, 211.7859, 211.6049, 
    211.4204, 211.2455, 211.0892, 210.966, 210.8799, 210.8439, 210.8643, 
    210.9417,
  212.5354, 212.4817, 212.4113, 212.2702, 212.0951, 211.9077, 211.7244, 
    211.5315, 211.3541, 211.1909, 211.0618, 210.9529, 210.8898, 210.8714, 
    210.9146,
  212.6841, 212.6321, 212.5859, 212.4764, 212.3373, 212.155, 211.9742, 
    211.7646, 211.5644, 211.3726, 211.2101, 211.0774, 210.9796, 210.9353, 
    210.9453,
  212.7662, 212.713, 212.6626, 212.5625, 212.458, 212.3191, 212.1624, 
    211.9626, 211.7517, 211.5294, 211.3341, 211.1674, 211.0392, 210.9597, 
    210.9365,
  212.8549, 212.8336, 212.7834, 212.6904, 212.5945, 212.4756, 212.3436, 
    212.1619, 211.9615, 211.7336, 211.5209, 211.326, 211.1642, 211.0468, 
    210.9881,
  212.832, 212.8363, 212.8215, 212.763, 212.6848, 212.5729, 212.4613, 
    212.3029, 212.1216, 211.9032, 211.6795, 211.4677, 211.283, 211.1364, 
    211.0402,
  212.8364, 212.8626, 212.8911, 212.8576, 212.8052, 212.7174, 212.6144, 
    212.4696, 212.3111, 212.1137, 211.8976, 211.6741, 211.4616, 211.2843, 
    211.1539,
  212.8724, 212.9108, 212.9538, 212.9448, 212.9161, 212.847, 212.7272, 
    212.5994, 212.4516, 212.2867, 212.1055, 211.8876, 211.6768, 211.467, 
    211.3026,
  212.8948, 212.932, 213.0075, 213.0436, 213.0417, 212.9815, 212.8658, 
    212.7442, 212.6101, 212.4393, 212.282, 212.0935, 211.8944, 211.6906, 
    211.5042,
  209.0141, 209.0995, 209.2378, 209.4044, 209.5845, 209.7048, 209.803, 
    209.8261, 209.803, 209.7216, 209.6154, 209.4906, 209.3577, 209.2288, 
    209.1027,
  209.2437, 209.2075, 209.2933, 209.4286, 209.6014, 209.7706, 209.908, 
    209.978, 209.9921, 209.9364, 209.8388, 209.7134, 209.5873, 209.4627, 
    209.3383,
  209.3034, 209.2239, 209.2591, 209.3552, 209.51, 209.702, 209.8667, 
    209.9979, 210.0569, 210.0542, 209.9807, 209.8694, 209.7337, 209.615, 
    209.5047,
  209.5059, 209.3874, 209.3386, 209.365, 209.482, 209.6566, 209.8706, 
    210.0397, 210.179, 210.2285, 210.2114, 210.1279, 210.0056, 209.8733, 
    209.7505,
  209.7137, 209.534, 209.4324, 209.3736, 209.4285, 209.5647, 209.7673, 
    209.9762, 210.1474, 210.2593, 210.3041, 210.283, 210.2018, 210.0899, 
    209.968,
  209.9225, 209.7499, 209.6178, 209.4986, 209.4696, 209.5388, 209.6919, 
    209.903, 210.0938, 210.2584, 210.3468, 210.3941, 210.3787, 210.3176, 
    210.2187,
  210.0782, 209.9247, 209.766, 209.6348, 209.5519, 209.5326, 209.6106, 
    209.7754, 209.9923, 210.1688, 210.311, 210.376, 210.4111, 210.3993, 
    210.3555,
  210.2336, 210.0925, 209.9499, 209.8249, 209.7191, 209.6365, 209.6454, 
    209.7429, 209.9573, 210.1744, 210.3354, 210.4314, 210.4588, 210.4627, 
    210.4429,
  210.2659, 210.1789, 210.0707, 209.9451, 209.8458, 209.7681, 209.7139, 
    209.7488, 209.8991, 210.1217, 210.3322, 210.4798, 210.5409, 210.5519, 
    210.5379,
  210.2929, 210.2345, 210.1729, 210.0864, 210.0106, 209.932, 209.8258, 
    209.7878, 209.8542, 209.9853, 210.1891, 210.3921, 210.5374, 210.6155, 
    210.6426,
  212.1442, 211.9078, 211.6787, 211.4323, 211.2095, 211.0075, 210.8417, 
    210.7123, 210.6206, 210.569, 210.5463, 210.5343, 210.532, 210.5192, 
    210.4967,
  212.4529, 212.2545, 212.0075, 211.7686, 211.5372, 211.3297, 211.1337, 
    210.9674, 210.8389, 210.7399, 210.6915, 210.6685, 210.6743, 210.6828, 
    210.6826,
  212.4369, 212.3133, 212.101, 211.8771, 211.6533, 211.4514, 211.2606, 
    211.0798, 210.9232, 210.7989, 210.7185, 210.685, 210.6899, 210.7118, 
    210.7362,
  212.5861, 212.4827, 212.2953, 212.0916, 211.8923, 211.7016, 211.5225, 
    211.3372, 211.1574, 210.987, 210.8615, 210.7916, 210.7749, 210.7898, 
    210.8191,
  212.5764, 212.4864, 212.325, 212.1406, 211.9757, 211.8146, 211.6644, 
    211.4878, 211.3072, 211.1251, 210.9639, 210.8533, 210.8064, 210.8035, 
    210.8266,
  212.64, 212.5728, 212.442, 212.2609, 212.1063, 211.9724, 211.8478, 
    211.7006, 211.5307, 211.3334, 211.1476, 211.0044, 210.9134, 210.8741, 
    210.8663,
  212.6111, 212.5648, 212.4664, 212.3067, 212.1616, 212.0296, 211.937, 
    211.8249, 211.6847, 211.5074, 211.31, 211.138, 211.0083, 210.9267, 
    210.8896,
  212.6423, 212.633, 212.5665, 212.4208, 212.2717, 212.1323, 212.0471, 
    211.9612, 211.8516, 211.7055, 211.5133, 211.3247, 211.1639, 211.0452, 
    210.9642,
  212.6217, 212.6427, 212.6242, 212.5006, 212.3649, 212.224, 212.1266, 
    212.0623, 211.9785, 211.8579, 211.6926, 211.4983, 211.3258, 211.1699, 
    211.0701,
  212.6081, 212.6634, 212.6912, 212.6157, 212.4984, 212.3416, 212.2318, 
    212.1634, 212.1253, 212.0206, 211.8926, 211.7041, 211.5139, 211.3455, 
    211.216,
  211.8876, 211.8495, 211.8293, 211.7646, 211.7164, 211.6585, 211.6168, 
    211.585, 211.5679, 211.5587, 211.5594, 211.5806, 211.6295, 211.6891, 
    211.7541,
  212.079, 212.054, 212.0363, 211.9821, 211.9401, 211.8806, 211.8407, 
    211.8098, 211.7976, 211.7965, 211.8136, 211.8362, 211.8792, 211.9278, 
    211.9825,
  212.15, 212.1481, 212.1419, 212.1025, 212.0594, 212.007, 211.9666, 211.934, 
    211.9283, 211.9292, 211.9504, 211.9655, 211.9905, 212.0278, 212.0764,
  212.2787, 212.2854, 212.3057, 212.2797, 212.254, 212.201, 212.1676, 
    212.1248, 212.1096, 212.1016, 212.1126, 212.1193, 212.1286, 212.149, 
    212.1879,
  212.3417, 212.3433, 212.3792, 212.3659, 212.3589, 212.321, 212.297, 
    212.2609, 212.2344, 212.2174, 212.2135, 212.2124, 212.2138, 212.2286, 
    212.2563,
  212.4595, 212.4555, 212.5001, 212.4921, 212.5008, 212.4806, 212.4741, 
    212.447, 212.4264, 212.3984, 212.3855, 212.3737, 212.3616, 212.3629, 
    212.3848,
  212.5447, 212.509, 212.5468, 212.5555, 212.5742, 212.5706, 212.5802, 
    212.5811, 212.5784, 212.5599, 212.5391, 212.521, 212.4994, 212.4853, 
    212.4886,
  212.676, 212.6347, 212.6566, 212.6504, 212.6629, 212.6701, 212.7023, 
    212.7107, 212.7355, 212.7433, 212.7381, 212.7206, 212.6964, 212.674, 
    212.6551,
  212.7912, 212.7507, 212.7416, 212.7271, 212.7402, 212.7401, 212.7586, 
    212.7905, 212.8277, 212.8617, 212.8877, 212.8869, 212.8744, 212.856, 
    212.8366,
  212.9465, 212.8887, 212.8841, 212.8779, 212.8609, 212.8297, 212.8426, 
    212.8666, 212.9158, 212.9572, 213.0154, 213.0414, 213.0454, 213.0385, 
    213.0308,
  211.74, 211.7443, 211.7417, 211.7043, 211.6287, 211.5091, 211.3593, 
    211.1769, 210.9856, 210.7739, 210.5597, 210.3472, 210.1409, 209.944, 
    209.7726,
  211.8221, 211.8316, 211.8304, 211.8364, 211.7961, 211.715, 211.5945, 
    211.4341, 211.26, 211.0625, 210.8512, 210.6343, 210.4105, 210.1945, 
    209.9895,
  211.7834, 211.7485, 211.7378, 211.7628, 211.7612, 211.7283, 211.6493, 
    211.5316, 211.3893, 211.221, 211.0293, 210.8266, 210.6155, 210.3988, 
    210.1908,
  211.8999, 211.8298, 211.7849, 211.7781, 211.7952, 211.7988, 211.753, 
    211.6675, 211.5408, 211.3982, 211.2325, 211.0463, 210.8461, 210.6432, 
    210.431,
  211.9549, 211.8643, 211.7971, 211.767, 211.7542, 211.7753, 211.7593, 
    211.7037, 211.5964, 211.4665, 211.3304, 211.1813, 211.0112, 210.8354, 
    210.6414,
  212.0636, 211.9744, 211.8802, 211.8157, 211.7787, 211.7988, 211.8001, 
    211.7685, 211.6815, 211.5598, 211.4265, 211.2965, 211.1568, 211.0098, 
    210.8361,
  212.0989, 212.0216, 211.9218, 211.8489, 211.7883, 211.7841, 211.7935, 
    211.78, 211.7177, 211.6052, 211.4732, 211.3527, 211.2358, 211.1208, 
    210.989,
  212.1464, 212.0982, 212.0114, 211.9105, 211.8269, 211.8139, 211.8183, 
    211.8086, 211.7673, 211.6796, 211.5451, 211.4205, 211.3136, 211.2195, 
    211.1217,
  212.1452, 212.1281, 212.0403, 211.9454, 211.8685, 211.8253, 211.8076, 
    211.8119, 211.7871, 211.7136, 211.6036, 211.4681, 211.3613, 211.2838, 
    211.2169,
  212.1404, 212.1427, 212.0782, 212.0291, 211.9285, 211.853, 211.8285, 
    211.8343, 211.8185, 211.7633, 211.6586, 211.5326, 211.4145, 211.3428, 
    211.2933,
  211.846, 211.7386, 211.6261, 211.4713, 211.3214, 211.1516, 211.0133, 
    210.9146, 210.8672, 210.8606, 210.886, 210.9319, 210.9782, 211.0226, 
    211.0579,
  212.0621, 211.9493, 211.8472, 211.6931, 211.5458, 211.3692, 211.2069, 
    211.0699, 210.9949, 210.9655, 210.979, 211.0221, 211.0833, 211.1404, 
    211.1874,
  212.1283, 212.043, 211.9643, 211.8237, 211.6844, 211.5242, 211.3506, 
    211.1899, 211.0722, 211.0121, 211.0052, 211.0333, 211.0905, 211.1576, 
    211.2201,
  212.2686, 212.202, 212.1515, 212.0245, 211.8914, 211.7401, 211.5748, 
    211.4035, 211.2559, 211.1551, 211.1173, 211.1279, 211.1696, 211.2353, 
    211.2977,
  212.2854, 212.2617, 212.2361, 212.1381, 212.023, 211.8811, 211.7309, 
    211.5639, 211.399, 211.2689, 211.203, 211.1863, 211.2148, 211.2702, 211.34,
  212.3309, 212.3518, 212.3407, 212.2789, 212.192, 212.0665, 211.9332, 
    211.7693, 211.6018, 211.4413, 211.3361, 211.2956, 211.3058, 211.3563, 
    211.4229,
  212.2974, 212.3433, 212.3634, 212.3376, 212.2981, 212.1911, 212.0767, 
    211.9353, 211.7727, 211.5993, 211.4568, 211.3804, 211.3715, 211.4114, 
    211.4757,
  212.2576, 212.3472, 212.3957, 212.4003, 212.3933, 212.3376, 212.2579, 
    212.1349, 211.982, 211.8099, 211.6412, 211.5164, 211.466, 211.4882, 
    211.5432,
  212.1748, 212.3047, 212.3718, 212.4052, 212.4411, 212.4246, 212.3806, 
    212.3033, 212.1753, 211.9959, 211.8206, 211.6606, 211.566, 211.5495, 
    211.5934,
  212.1281, 212.2427, 212.3493, 212.4125, 212.4671, 212.4763, 212.4912, 
    212.4686, 212.3767, 212.2159, 212.0352, 211.8516, 211.7165, 211.657, 
    211.6669,
  210.2915, 210.1856, 210.1198, 210.0507, 209.9913, 209.9399, 209.8902, 
    209.8412, 209.7935, 209.76, 209.764, 209.7957, 209.8119, 209.784, 209.6946,
  210.4222, 210.3044, 210.2027, 210.1329, 210.0848, 210.0502, 210.0105, 
    209.9653, 209.9118, 209.864, 209.8329, 209.8269, 209.8429, 209.8464, 
    209.8207,
  210.4424, 210.3055, 210.199, 210.1146, 210.074, 210.0643, 210.0535, 
    210.0238, 209.9846, 209.9375, 209.8915, 209.8595, 209.862, 209.8784, 
    209.8905,
  210.5769, 210.4396, 210.2998, 210.1837, 210.1378, 210.1268, 210.1345, 
    210.139, 210.1167, 210.0829, 210.0409, 210.0064, 209.9869, 209.9987, 
    210.0135,
  210.6183, 210.4786, 210.3311, 210.2089, 210.1424, 210.127, 210.1485, 
    210.1814, 210.187, 210.1692, 210.1371, 210.0988, 210.0783, 210.0689, 
    210.0803,
  210.7023, 210.5622, 210.3947, 210.2566, 210.1542, 210.1322, 210.1588, 
    210.217, 210.2585, 210.2737, 210.263, 210.2268, 210.1907, 210.1698, 
    210.1599,
  210.7284, 210.5857, 210.4133, 210.2763, 210.1496, 210.0867, 210.1002, 
    210.1581, 210.2299, 210.2809, 210.3044, 210.301, 210.2708, 210.2474, 
    210.2281,
  210.8069, 210.6585, 210.4979, 210.3449, 210.1947, 210.0958, 210.0804, 
    210.1162, 210.1953, 210.285, 210.3318, 210.3625, 210.3537, 210.3306, 
    210.3115,
  210.8574, 210.7134, 210.5596, 210.4009, 210.2631, 210.1391, 210.0629, 
    210.0831, 210.1319, 210.2362, 210.3169, 210.3643, 210.3955, 210.3856, 
    210.377,
  210.9216, 210.7779, 210.6454, 210.5231, 210.3661, 210.21, 210.109, 
    210.0907, 210.1238, 210.2063, 210.3139, 210.3894, 210.446, 210.4672, 
    210.4675,
  211.0997, 210.929, 210.776, 210.6533, 210.5741, 210.5468, 210.5382, 
    210.5459, 210.5626, 210.5604, 210.5632, 210.5859, 210.6086, 210.6638, 
    210.7219,
  211.4407, 211.2266, 211.0619, 210.9064, 210.791, 210.7226, 210.6972, 
    210.6944, 210.7057, 210.7092, 210.7138, 210.7177, 210.7197, 210.7519, 
    210.791,
  211.6281, 211.4204, 211.2733, 211.0899, 210.9456, 210.8509, 210.8043, 
    210.7981, 210.8089, 210.8208, 210.8367, 210.8389, 210.8468, 210.858, 
    210.8876,
  211.816, 211.6701, 211.5576, 211.387, 211.2305, 211.0929, 211.0113, 
    210.962, 210.9604, 210.9795, 211.0108, 211.0314, 211.0467, 211.0552, 
    211.0708,
  211.9559, 211.85, 211.7588, 211.6011, 211.425, 211.2488, 211.1338, 
    211.0507, 211.0208, 211.0311, 211.0663, 211.0969, 211.1148, 211.1302, 
    211.1272,
  212.1308, 212.0424, 211.9723, 211.8289, 211.6801, 211.5082, 211.3751, 
    211.2694, 211.1896, 211.1646, 211.1779, 211.2155, 211.2348, 211.2592, 
    211.2473,
  212.2439, 212.1678, 212.1336, 212.0289, 211.9056, 211.7311, 211.58, 
    211.4455, 211.3526, 211.2892, 211.2769, 211.2951, 211.3219, 211.3415, 
    211.3462,
  212.3585, 212.3158, 212.2985, 212.2184, 212.1215, 211.9853, 211.8277, 
    211.6902, 211.5788, 211.5144, 211.4669, 211.4628, 211.4673, 211.479, 
    211.4779,
  212.417, 212.3734, 212.3788, 212.3262, 212.2834, 212.1779, 212.0359, 
    211.8827, 211.7655, 211.6763, 211.6308, 211.6005, 211.5905, 211.5875, 
    211.5723,
  212.505, 212.4687, 212.4955, 212.4743, 212.4478, 212.3465, 212.2321, 
    212.09, 211.9518, 211.8372, 211.7779, 211.7391, 211.7213, 211.7091, 
    211.6871,
  208.429, 208.3677, 208.3725, 208.3926, 208.436, 208.4671, 208.5057, 
    208.5251, 208.535, 208.5196, 208.4848, 208.4364, 208.3847, 208.3355, 
    208.3036,
  208.3809, 208.3574, 208.353, 208.3662, 208.3863, 208.4047, 208.4388, 
    208.4932, 208.5509, 208.5855, 208.5877, 208.5579, 208.513, 208.4704, 
    208.431,
  208.4592, 208.3923, 208.3123, 208.2968, 208.3365, 208.4024, 208.4749, 
    208.5525, 208.6263, 208.6781, 208.6995, 208.6803, 208.6395, 208.5922, 
    208.551,
  208.5214, 208.4387, 208.3735, 208.3895, 208.4326, 208.4878, 208.5327, 
    208.59, 208.6552, 208.7248, 208.7716, 208.78, 208.7543, 208.7104, 208.6626,
  208.545, 208.4826, 208.4141, 208.3451, 208.2932, 208.2862, 208.3168, 
    208.3874, 208.4747, 208.5782, 208.6687, 208.7312, 208.7504, 208.7493, 
    208.7269,
  208.6217, 208.5489, 208.4476, 208.3465, 208.3042, 208.3044, 208.3568, 
    208.4254, 208.5134, 208.6048, 208.6973, 208.7656, 208.7962, 208.7926, 
    208.7719,
  208.6696, 208.5862, 208.4882, 208.408, 208.3385, 208.2864, 208.2776, 
    208.3176, 208.3996, 208.5002, 208.6045, 208.6974, 208.7714, 208.8106, 
    208.82,
  208.6795, 208.621, 208.5221, 208.4205, 208.3054, 208.2245, 208.1915, 
    208.197, 208.2831, 208.3858, 208.5051, 208.6222, 208.7374, 208.8216, 
    208.8611,
  208.6622, 208.6323, 208.5589, 208.4678, 208.3833, 208.2909, 208.2084, 
    208.1746, 208.2019, 208.2936, 208.4221, 208.5526, 208.688, 208.7968, 
    208.8686,
  208.7001, 208.7003, 208.6566, 208.5781, 208.462, 208.3397, 208.231, 
    208.1836, 208.1793, 208.2368, 208.3487, 208.4871, 208.6395, 208.7819, 
    208.889,
  211.4837, 211.3156, 211.1459, 210.9528, 210.7607, 210.5791, 210.4233, 
    210.2979, 210.2067, 210.1498, 210.1171, 210.0887, 210.0604, 210.0316, 
    210.0044,
  211.7743, 211.6491, 211.5013, 211.3154, 211.1096, 210.8899, 210.6859, 
    210.5149, 210.3893, 210.305, 210.2542, 210.2241, 210.1995, 210.1778, 
    210.1468,
  211.8242, 211.746, 211.655, 211.4817, 211.2948, 211.0857, 210.8938, 
    210.7185, 210.5736, 210.4527, 210.3754, 210.3365, 210.319, 210.304, 
    210.2755,
  211.9551, 211.9126, 211.8622, 211.7371, 211.5853, 211.3812, 211.1676, 
    210.9601, 210.7816, 210.6379, 210.548, 210.5019, 210.4717, 210.4572, 
    210.4274,
  212.1386, 212.1151, 212.0681, 211.9762, 211.8444, 211.6504, 211.4361, 
    211.2171, 211.0229, 210.8626, 210.7226, 210.6267, 210.5628, 210.5248, 
    210.4882,
  212.1767, 212.1468, 212.1337, 212.1014, 212.0199, 211.9034, 211.7386, 
    211.53, 211.3027, 211.0821, 210.9093, 210.7916, 210.7262, 210.6892, 
    210.6501,
  212.2176, 212.2401, 212.2705, 212.2842, 212.2446, 212.1265, 211.9692, 
    211.753, 211.5252, 211.2953, 211.0973, 210.9566, 210.8588, 210.8046, 
    210.7582,
  212.2741, 212.3197, 212.3495, 212.3754, 212.3955, 212.3439, 212.2263, 
    212.0596, 211.8531, 211.613, 211.3717, 211.1629, 211.0275, 210.9305, 
    210.8741,
  212.2177, 212.2672, 212.3193, 212.3706, 212.4448, 212.4887, 212.4322, 
    212.3051, 212.1072, 211.8595, 211.6024, 211.368, 211.1918, 211.0731, 
    210.9988,
  212.2046, 212.2831, 212.3521, 212.4292, 212.5172, 212.5889, 212.5951, 
    212.517, 212.3671, 212.1387, 211.8839, 211.6229, 211.4037, 211.2511, 
    211.1481,
  208.9654, 208.9964, 209.0713, 209.1311, 209.16, 209.1423, 209.0744, 
    208.9524, 208.8246, 208.703, 208.6158, 208.5728, 208.5771, 208.6218, 
    208.6791,
  208.9949, 209.0256, 209.0963, 209.1798, 209.257, 209.2869, 209.2715, 
    209.1898, 209.0952, 208.9865, 208.8868, 208.8089, 208.7613, 208.751, 
    208.7699,
  209.0021, 208.9979, 209.0466, 209.1131, 209.1957, 209.2715, 209.2956, 
    209.2548, 209.1807, 209.0871, 208.9917, 208.9086, 208.8505, 208.8358, 
    208.8586,
  209.0606, 209.0413, 209.0527, 209.0898, 209.1675, 209.2601, 209.3375, 
    209.3443, 209.3088, 209.2234, 209.1397, 209.0436, 209.004, 208.989, 
    209.0084,
  209.0542, 209.0292, 209.0407, 209.0712, 209.1345, 209.2328, 209.3384, 
    209.3917, 209.3828, 209.3114, 209.2171, 209.1165, 209.0376, 209.0099, 
    209.0023,
  209.1122, 209.0881, 209.0775, 209.0681, 209.0898, 209.1668, 209.3003, 
    209.4014, 209.4617, 209.4438, 209.3653, 209.2639, 209.1657, 209.0875, 
    209.0603,
  209.1612, 209.1259, 209.114, 209.1055, 209.0995, 209.1103, 209.1979, 
    209.3151, 209.4231, 209.478, 209.4656, 209.3885, 209.2929, 209.1966, 
    209.1245,
  209.1419, 209.0917, 209.0711, 209.0692, 209.0719, 209.0739, 209.12, 
    209.221, 209.3461, 209.4609, 209.5164, 209.5038, 209.4367, 209.3482, 
    209.2744,
  209.1352, 209.0582, 209.0024, 208.9612, 208.9799, 209.0106, 209.0456, 
    209.1092, 209.2259, 209.3452, 209.4583, 209.5062, 209.5025, 209.4395, 
    209.3772,
  209.2332, 209.1292, 209.0635, 209.0157, 209.0204, 209.0312, 209.0485, 
    209.0894, 209.1651, 209.2571, 209.3712, 209.4722, 209.5266, 209.536, 
    209.4885,
  212.2849, 212.1564, 212.0006, 211.8063, 211.6161, 211.4541, 211.3306, 
    211.2286, 211.144, 211.0651, 210.9901, 210.9096, 210.8283, 210.7403, 
    210.6436,
  212.5236, 212.4025, 212.2796, 212.1022, 211.9248, 211.745, 211.6083, 
    211.4866, 211.3847, 211.2841, 211.1917, 211.1035, 211.012, 210.923, 
    210.8212,
  212.5621, 212.4807, 212.403, 212.2599, 212.1016, 211.9217, 211.7685, 
    211.6338, 211.5206, 211.4106, 211.3069, 211.2094, 211.1062, 211.0104, 
    210.906,
  212.6894, 212.6304, 212.576, 212.4719, 212.3456, 212.1777, 212.0175, 
    211.8672, 211.7391, 211.6306, 211.5192, 211.4068, 211.2861, 211.1752, 
    211.0579,
  212.6958, 212.6578, 212.6207, 212.5444, 212.4593, 212.3218, 212.1648, 
    212.0088, 211.8622, 211.7401, 211.6245, 211.5117, 211.3941, 211.2842, 
    211.1709,
  212.7768, 212.7533, 212.7257, 212.6575, 212.5831, 212.4836, 212.3519, 
    212.1925, 212.0332, 211.9052, 211.7916, 211.684, 211.5775, 211.4681, 
    211.3548,
  212.8128, 212.7745, 212.7438, 212.6922, 212.6327, 212.5435, 212.4353, 
    212.2954, 212.1465, 212.0005, 211.8698, 211.7728, 211.6748, 211.5851, 
    211.482,
  212.8608, 212.8327, 212.8022, 212.7554, 212.7023, 212.6319, 212.538, 
    212.4188, 212.2841, 212.1382, 212.0009, 211.8828, 211.7947, 211.7075, 
    211.6056,
  212.8444, 212.8406, 212.8297, 212.7768, 212.7328, 212.6877, 212.5873, 
    212.4763, 212.3583, 212.2183, 212.0934, 211.965, 211.8763, 211.7869, 
    211.703,
  212.8419, 212.8485, 212.855, 212.8384, 212.8074, 212.7522, 212.6459, 
    212.5381, 212.4414, 212.2934, 212.1658, 212.0403, 211.9375, 211.8613, 
    211.7945,
  210.5735, 210.5497, 210.4642, 210.2974, 210.0896, 209.8531, 209.6299, 
    209.4251, 209.2717, 209.1641, 209.1156, 209.112, 209.1445, 209.1981, 
    209.2672,
  210.6629, 210.6915, 210.6925, 210.5977, 210.4432, 210.2088, 209.9662, 
    209.7308, 209.5506, 209.4153, 209.3436, 209.3166, 209.3299, 209.3681, 
    209.4275,
  210.5797, 210.63, 210.6909, 210.668, 210.5911, 210.4207, 210.2093, 209.983, 
    209.7866, 209.6343, 209.5408, 209.4918, 209.4874, 209.5104, 209.558,
  210.6095, 210.6691, 210.7512, 210.787, 210.7884, 210.6756, 210.5097, 
    210.2913, 210.0878, 209.9124, 209.7982, 209.7262, 209.6998, 209.7052, 
    209.7369,
  210.5361, 210.5932, 210.6835, 210.7563, 210.8257, 210.7909, 210.6906, 
    210.5036, 210.3079, 210.1219, 209.9886, 209.9056, 209.8736, 209.8751, 
    209.9021,
  210.5366, 210.5778, 210.6691, 210.7484, 210.8515, 210.8883, 210.8624, 
    210.7373, 210.5603, 210.3751, 210.2174, 210.1167, 210.0715, 210.071, 
    210.1024,
  210.4662, 210.4974, 210.5841, 210.6814, 210.7978, 210.8784, 210.9184, 
    210.8649, 210.7426, 210.5711, 210.4142, 210.2961, 210.2444, 210.2369, 
    210.2753,
  210.4082, 210.4539, 210.5479, 210.6356, 210.7515, 210.8567, 210.9492, 
    210.9625, 210.8998, 210.7716, 210.6193, 210.4959, 210.4298, 210.4218, 
    210.4624,
  210.3388, 210.401, 210.4717, 210.548, 210.6696, 210.7717, 210.8945, 
    210.9802, 210.9778, 210.8988, 210.7792, 210.6613, 210.5911, 210.5699, 
    210.6101,
  210.2928, 210.3758, 210.455, 210.5448, 210.6337, 210.69, 210.8018, 
    210.9572, 211.0118, 210.9915, 210.9245, 210.8222, 210.7584, 210.7276, 
    210.755,
  211.2321, 210.9914, 210.6926, 210.3775, 210.0827, 209.8247, 209.6315, 
    209.4809, 209.3736, 209.2863, 209.2131, 209.1415, 209.0656, 208.976, 
    208.869,
  211.531, 211.3357, 211.0526, 210.7457, 210.4178, 210.1152, 209.8609, 
    209.672, 209.5353, 209.4388, 209.3613, 209.2921, 209.2213, 209.1369, 
    209.04,
  211.5459, 211.4027, 211.1878, 210.9171, 210.5968, 210.2787, 209.9938, 
    209.7774, 209.6172, 209.5118, 209.4358, 209.3753, 209.3167, 209.2496, 
    209.1694,
  211.6657, 211.5593, 211.3914, 211.1547, 210.856, 210.5319, 210.2198, 
    209.9684, 209.7873, 209.6658, 209.5876, 209.5302, 209.4796, 209.4178, 
    209.345,
  211.6551, 211.585, 211.4676, 211.277, 211.0202, 210.7103, 210.3953, 
    210.1088, 209.8885, 209.7441, 209.6566, 209.6034, 209.5618, 209.5147, 
    209.4558,
  211.6756, 211.634, 211.5577, 211.4119, 211.205, 210.9368, 210.6305, 
    210.3276, 210.0684, 209.8827, 209.7681, 209.7041, 209.665, 209.6235, 
    209.5724,
  211.631, 211.5904, 211.5447, 211.4542, 211.3021, 211.0867, 210.8178, 
    210.5312, 210.2579, 210.0374, 209.8881, 209.8002, 209.7551, 209.7182, 
    209.6737,
  211.6505, 211.6024, 211.5603, 211.4939, 211.3728, 211.2199, 210.9991, 
    210.7321, 210.4705, 210.233, 210.0558, 209.9443, 209.8734, 209.8406, 
    209.7915,
  211.6614, 211.6007, 211.5389, 211.4828, 211.4067, 211.285, 211.11, 
    210.8928, 210.6464, 210.4111, 210.2119, 210.0716, 209.9888, 209.9412, 
    209.896,
  211.7415, 211.6519, 211.5758, 211.5461, 211.4574, 211.3374, 211.1926, 
    211.0293, 210.814, 210.5889, 210.3802, 210.2179, 210.1125, 210.0421, 
    209.998,
  210.4593, 210.5325, 210.6073, 210.588, 210.5421, 210.4423, 210.3434, 
    210.2271, 210.1222, 210.0162, 209.9234, 209.8177, 209.7227, 209.6499, 
    209.6126,
  210.6388, 210.6869, 210.7912, 210.8047, 210.8061, 210.7205, 210.6287, 
    210.4885, 210.3666, 210.2415, 210.1198, 209.9988, 209.8781, 209.7797, 
    209.7215,
  210.633, 210.6922, 210.801, 210.8281, 210.8657, 210.8262, 210.7556, 
    210.6464, 210.5321, 210.4118, 210.295, 210.18, 210.0595, 209.9589, 209.888,
  210.7098, 210.8205, 210.9494, 210.9888, 211.0176, 210.9667, 210.8942, 
    210.7898, 210.6763, 210.5674, 210.4632, 210.3591, 210.2543, 210.1557, 
    210.0732,
  210.6701, 210.8323, 211.0045, 211.0701, 211.0906, 211.0584, 210.9986, 
    210.8926, 210.7833, 210.6607, 210.5565, 210.4455, 210.3406, 210.239, 
    210.1537,
  210.7339, 210.8786, 211.0647, 211.1509, 211.1867, 211.1586, 211.1123, 
    211.0234, 210.9302, 210.8102, 210.7042, 210.5941, 210.4914, 210.3853, 
    210.2937,
  210.7062, 210.8304, 211.0387, 211.1779, 211.2501, 211.2282, 211.1969, 
    211.1205, 211.0366, 210.9202, 210.8109, 210.7021, 210.5919, 210.4836, 
    210.3856,
  210.654, 210.8015, 211.0287, 211.1868, 211.301, 211.34, 211.3288, 211.2502, 
    211.1742, 211.0692, 210.9587, 210.8442, 210.731, 210.6205, 210.5181,
  210.5943, 210.7508, 210.9495, 211.1265, 211.3135, 211.4, 211.3955, 
    211.3468, 211.2571, 211.1743, 211.0752, 210.971, 210.8673, 210.7529, 
    210.6519,
  210.565, 210.7146, 210.9159, 211.15, 211.3438, 211.4495, 211.4936, 
    211.4514, 211.3752, 211.2694, 211.1834, 211.0827, 210.9808, 210.8681, 
    210.7669,
  210.979, 210.8012, 210.6509, 210.4894, 210.3787, 210.287, 210.234, 
    210.1663, 210.1127, 210.0761, 210.0535, 210.0409, 210.037, 210.0136, 
    209.9575,
  211.0493, 210.8744, 210.7504, 210.6164, 210.5128, 210.4091, 210.326, 
    210.2457, 210.1806, 210.1083, 210.0517, 210.0222, 210.0237, 210.0324, 
    210.0208,
  211.0348, 210.901, 210.8111, 210.6996, 210.6185, 210.5228, 210.4447, 
    210.3646, 210.2942, 210.2126, 210.1426, 210.0941, 210.0788, 210.0853, 
    210.0858,
  211.1734, 211.0775, 211.0059, 210.9232, 210.847, 210.7197, 210.6124, 
    210.5162, 210.4497, 210.387, 210.3203, 210.2578, 210.2079, 210.1846, 
    210.1651,
  211.2423, 211.1775, 211.1358, 211.0225, 210.8995, 210.7337, 210.6119, 
    210.5115, 210.4488, 210.3882, 210.3363, 210.3136, 210.2897, 210.2646, 
    210.2338,
  211.3175, 211.1902, 211.1091, 210.963, 210.8599, 210.7576, 210.6703, 
    210.5781, 210.4806, 210.3996, 210.3362, 210.3053, 210.279, 210.2363, 
    210.195,
  211.3331, 211.1376, 211.0358, 210.9415, 210.895, 210.7987, 210.6873, 
    210.5819, 210.5069, 210.454, 210.3864, 210.3153, 210.2645, 210.2137, 
    210.1996,
  211.5083, 211.2884, 211.1535, 210.9998, 210.9133, 210.8217, 210.7317, 
    210.6675, 210.6497, 210.6162, 210.5259, 210.4047, 210.3199, 210.261, 
    210.2463,
  211.6694, 211.4327, 211.2689, 211.0731, 210.9893, 210.9405, 210.8615, 
    210.8074, 210.7752, 210.729, 210.6568, 210.5234, 210.4015, 210.3257, 
    210.2888,
  211.7776, 211.5406, 211.4017, 211.2323, 211.124, 211.0232, 210.911, 
    210.8186, 210.783, 210.6922, 210.6467, 210.5531, 210.4764, 210.4081, 
    210.3685,
  210.9548, 210.9052, 210.8532, 210.7576, 210.6924, 210.6151, 210.5585, 
    210.5078, 210.4778, 210.4624, 210.464, 210.4817, 210.5263, 210.5828, 
    210.627,
  211.1624, 211.1082, 211.0688, 210.9803, 210.8987, 210.7985, 210.725, 
    210.662, 210.6238, 210.5923, 210.5762, 210.5843, 210.6384, 210.7131, 
    210.778,
  211.1784, 211.1263, 211.1043, 211.0487, 210.9773, 210.8833, 210.8181, 
    210.7677, 210.7507, 210.7494, 210.7571, 210.8023, 210.873, 210.934, 
    210.9465,
  211.2974, 211.2446, 211.2134, 211.1692, 211.1087, 211.0303, 210.9751, 
    210.9457, 210.9504, 210.9677, 210.9896, 211.0406, 211.0982, 211.1409, 
    211.1257,
  211.3312, 211.2727, 211.2422, 211.194, 211.1412, 211.0671, 210.9923, 
    210.9567, 210.9604, 210.9545, 210.9391, 210.9464, 210.9913, 211.0878, 
    211.1374,
  211.4403, 211.3996, 211.378, 211.3088, 211.2454, 211.1646, 211.0833, 
    211.0074, 211.0112, 211.0123, 211.0221, 211.001, 210.9978, 211.0798, 
    211.1416,
  211.5153, 211.4932, 211.4732, 211.4232, 211.3778, 211.2639, 211.1563, 
    211.0465, 211.03, 211.0746, 211.1477, 211.1595, 211.1453, 211.1684, 
    211.1805,
  211.6029, 211.6164, 211.6242, 211.5999, 211.5629, 211.4539, 211.3273, 
    211.1721, 211.0786, 211.0688, 211.1203, 211.1689, 211.211, 211.2303, 
    211.2401,
  211.6083, 211.6772, 211.7166, 211.6855, 211.6649, 211.6232, 211.5001, 
    211.3324, 211.1808, 211.1041, 211.1249, 211.203, 211.2726, 211.2925, 
    211.2876,
  211.5917, 211.6843, 211.7622, 211.7717, 211.7664, 211.7131, 211.5941, 
    211.451, 211.3179, 211.1808, 211.1393, 211.1919, 211.2567, 211.299, 
    211.2983,
  209.5054, 209.4042, 209.3046, 209.163, 209.0253, 208.8633, 208.7186, 
    208.5634, 208.4193, 208.2618, 208.0971, 207.9394, 207.8119, 207.7513, 
    207.7323,
  209.7464, 209.6412, 209.5472, 209.4032, 209.2577, 209.081, 208.9247, 
    208.7683, 208.6271, 208.4801, 208.3291, 208.1893, 208.0685, 208.0211, 
    207.9753,
  209.7936, 209.7275, 209.6515, 209.5313, 209.3847, 209.2077, 209.0461, 
    208.8873, 208.7473, 208.6083, 208.4665, 208.3317, 208.2087, 208.1136, 
    208.0247,
  209.9298, 209.8866, 209.8345, 209.7268, 209.6009, 209.4213, 209.2497, 
    209.0831, 208.9361, 208.7966, 208.6567, 208.5019, 208.3517, 208.2116, 
    208.0887,
  209.983, 209.9395, 209.9081, 209.8331, 209.7303, 209.5737, 209.3965, 
    209.2224, 209.0649, 208.919, 208.7708, 208.6095, 208.4487, 208.3123, 
    208.2278,
  210.0807, 210.0334, 210.015, 209.9545, 209.876, 209.7501, 209.5866, 
    209.3997, 209.2281, 209.0659, 208.9147, 208.7533, 208.6004, 208.4667, 
    208.375,
  210.123, 210.0422, 210.0312, 210.0271, 209.9978, 209.8828, 209.7365, 
    209.5443, 209.3624, 209.1845, 209.0314, 208.8768, 208.7261, 208.5719, 
    208.4656,
  210.1635, 210.0741, 210.0597, 210.0979, 210.1116, 210.0491, 209.9194, 
    209.7231, 209.525, 209.3327, 209.1602, 209.0066, 208.8558, 208.7094, 
    208.5974,
  210.1952, 210.0921, 210.0681, 210.1158, 210.1914, 210.2163, 210.1148, 
    209.9356, 209.7161, 209.4973, 209.3117, 209.1344, 208.9847, 208.8478, 
    208.7327,
  210.2662, 210.1345, 210.1064, 210.1884, 210.2833, 210.3453, 210.3063, 
    210.1721, 209.9727, 209.7207, 209.5098, 209.3193, 209.1514, 209.0042, 
    208.8775,
  210.198, 210.129, 210.1107, 210.0715, 210.058, 210.0484, 210.0552, 
    210.0759, 210.104, 210.1191, 210.1106, 210.0765, 210.0066, 209.9064, 
    209.783,
  210.4635, 210.3876, 210.3583, 210.316, 210.2948, 210.2779, 210.2792, 
    210.2946, 210.3227, 210.3467, 210.3542, 210.3403, 210.294, 210.2162, 
    210.1114,
  210.5419, 210.5248, 210.505, 210.4753, 210.438, 210.4111, 210.4, 210.4152, 
    210.4441, 210.4872, 210.5222, 210.5433, 210.5301, 210.4798, 210.3992,
  210.7078, 210.7147, 210.704, 210.6845, 210.6495, 210.6066, 210.5729, 
    210.5691, 210.5898, 210.6259, 210.6694, 210.7113, 210.7268, 210.7174, 
    210.6697,
  210.7621, 210.7943, 210.7993, 210.7955, 210.768, 210.7288, 210.6768, 
    210.6517, 210.6632, 210.6961, 210.7477, 210.7985, 210.8395, 210.852, 
    210.8334,
  210.8632, 210.9048, 210.9296, 210.9314, 210.901, 210.859, 210.8048, 
    210.7557, 210.7468, 210.7717, 210.8279, 210.887, 210.943, 210.9775, 
    210.9821,
  210.9118, 210.9415, 210.991, 211.0218, 211.0168, 210.9569, 210.8961, 
    210.8308, 210.7956, 210.8014, 210.8441, 210.9171, 210.9902, 211.0468, 
    211.0688,
  211.0049, 211.0263, 211.0815, 211.1187, 211.1396, 211.1039, 211.054, 
    210.9759, 210.9099, 210.8752, 210.8939, 210.9441, 211.0304, 211.0989, 
    211.156,
  211.0692, 211.073, 211.1242, 211.1605, 211.2237, 211.2437, 211.214, 
    211.159, 211.0607, 210.9727, 210.9516, 210.9757, 211.0387, 211.1267, 
    211.1949,
  211.1939, 211.1368, 211.1863, 211.2452, 211.3158, 211.3563, 211.3784, 
    211.3475, 211.2673, 211.1395, 211.0502, 211.0372, 211.0664, 211.1483, 
    211.2323,
  209.5154, 209.5949, 209.7128, 209.765, 209.7632, 209.6609, 209.5037, 
    209.2618, 208.9965, 208.7166, 208.4608, 208.2436, 208.0807, 207.9696, 
    207.9132,
  209.5348, 209.605, 209.7422, 209.8374, 209.8988, 209.8709, 209.7643, 
    209.5739, 209.3267, 209.0432, 208.7758, 208.536, 208.3469, 208.2075, 
    208.1262,
  209.5165, 209.5915, 209.7143, 209.8469, 209.9407, 209.9742, 209.9282, 
    209.7812, 209.5699, 209.2928, 209.0163, 208.7646, 208.5589, 208.4067, 
    208.3096,
  209.5582, 209.6031, 209.6985, 209.8377, 209.9882, 210.0738, 210.0881, 
    210.0079, 209.8236, 209.5846, 209.2998, 209.0478, 208.8199, 208.6585, 
    208.5451,
  209.625, 209.601, 209.6536, 209.7742, 209.9426, 210.0812, 210.163, 
    210.1554, 210.0445, 209.8287, 209.5683, 209.2844, 209.0639, 208.8703, 
    208.755,
  209.7483, 209.6623, 209.6528, 209.7164, 209.8657, 210.0546, 210.2124, 
    210.2807, 210.2472, 210.0896, 209.8549, 209.5692, 209.3106, 209.0988, 
    208.9457,
  209.8548, 209.726, 209.6484, 209.6682, 209.7769, 209.9498, 210.1544, 
    210.3191, 210.3905, 210.316, 210.1228, 209.8436, 209.5418, 209.2892, 
    209.0997,
  209.9857, 209.8426, 209.7306, 209.6744, 209.7162, 209.8547, 210.096, 
    210.31, 210.4674, 210.4742, 210.3404, 210.1006, 209.7857, 209.4907, 
    209.268,
  210.0961, 209.9715, 209.8222, 209.6803, 209.681, 209.7991, 209.9852, 
    210.2334, 210.4224, 210.5288, 210.493, 210.3026, 210.008, 209.6994, 
    209.4513,
  210.2012, 210.0974, 209.9769, 209.8442, 209.7818, 209.7744, 209.9004, 
    210.1342, 210.3791, 210.5337, 210.5857, 210.4709, 210.2496, 209.9732, 
    209.7041,
  210.9946, 211.0579, 211.1549, 211.2555, 211.3644, 211.4682, 211.583, 
    211.6924, 211.799, 211.8888, 211.956, 211.9888, 211.9808, 211.9293, 
    211.8333,
  211.0812, 211.101, 211.1629, 211.2489, 211.3558, 211.471, 211.5949, 
    211.721, 211.8452, 211.9639, 212.0571, 212.1199, 212.1477, 212.1277, 
    212.0572,
  211.0545, 211.0507, 211.0785, 211.1444, 211.2282, 211.3433, 211.4662, 
    211.5945, 211.7306, 211.869, 212.005, 212.1113, 212.1889, 212.2142, 
    212.1777,
  211.1136, 211.0872, 211.0876, 211.1419, 211.2258, 211.3258, 211.4462, 
    211.5545, 211.6774, 211.8066, 211.9562, 212.0973, 212.2089, 212.2725, 
    212.2744,
  211.1253, 211.0646, 211.0362, 211.0544, 211.1317, 211.2197, 211.3352, 
    211.4419, 211.5469, 211.6735, 211.8245, 211.998, 212.1534, 212.2616, 
    212.3073,
  211.2669, 211.1406, 211.0786, 211.0407, 211.0757, 211.172, 211.2771, 
    211.3897, 211.4803, 211.5856, 211.7249, 211.9007, 212.082, 212.224, 
    212.3127,
  211.4078, 211.201, 211.0905, 211.015, 211.0196, 211.0656, 211.1601, 
    211.2692, 211.3795, 211.4829, 211.609, 211.7739, 211.9553, 212.1263, 
    212.2483,
  211.5973, 211.3884, 211.1993, 211.0731, 211.0075, 211.0233, 211.0954, 
    211.178, 211.2862, 211.4002, 211.514, 211.6668, 211.8355, 212.0126, 
    212.1658,
  211.7228, 211.5668, 211.3585, 211.1461, 211.0285, 210.9884, 211.0162, 
    211.0906, 211.1768, 211.2935, 211.4189, 211.5609, 211.7161, 211.879, 
    212.0471,
  211.8307, 211.7305, 211.5767, 211.3606, 211.1739, 211.0274, 210.972, 
    211.0087, 211.1169, 211.2044, 211.3504, 211.4863, 211.6264, 211.7656, 
    211.9206,
  210.0089, 210.1717, 210.3584, 210.5117, 210.6323, 210.6794, 210.6804, 
    210.6215, 210.5238, 210.3772, 210.2077, 210.025, 209.8552, 209.7081, 
    209.6034,
  210.0738, 210.2042, 210.369, 210.5361, 210.6946, 210.7957, 210.8532, 
    210.8286, 210.7605, 210.6333, 210.4932, 210.3369, 210.1844, 210.0372, 
    209.9106,
  210.1064, 210.2083, 210.3627, 210.5159, 210.6782, 210.8101, 210.9114, 
    210.9493, 210.9362, 210.8498, 210.7229, 210.5679, 210.4104, 210.2597, 
    210.127,
  210.1637, 210.2443, 210.3869, 210.5316, 210.7003, 210.8608, 211.0067, 
    211.0954, 211.1234, 211.066, 210.9382, 210.7809, 210.6172, 210.4721, 
    210.3505,
  210.2258, 210.261, 210.3814, 210.5226, 210.691, 210.8637, 211.0284, 
    211.149, 211.2077, 211.1888, 211.106, 210.9734, 210.8331, 210.7004, 
    210.5786,
  210.3414, 210.345, 210.4316, 210.5214, 210.6578, 210.841, 211.013, 
    211.1463, 211.2404, 211.2681, 211.2368, 211.1565, 211.0471, 210.9307, 
    210.8156,
  210.4414, 210.4035, 210.441, 210.5085, 210.6559, 210.7984, 210.9618, 
    211.1027, 211.2164, 211.2842, 211.3027, 211.2656, 211.1931, 211.0971, 
    210.9961,
  210.5354, 210.4789, 210.4844, 210.5372, 210.653, 210.77, 210.914, 211.0497, 
    211.1845, 211.2932, 211.3536, 211.3619, 211.3223, 211.2509, 211.1625,
  210.5916, 210.5403, 210.5395, 210.5379, 210.621, 210.7653, 210.8942, 
    211.013, 211.1459, 211.2547, 211.3564, 211.3983, 211.3939, 211.3413, 
    211.2719,
  210.6342, 210.5869, 210.5933, 210.615, 210.6789, 210.7998, 210.8773, 
    210.9813, 211.1219, 211.2203, 211.3262, 211.4008, 211.4224, 211.3966, 
    211.3476,
  211.3759, 211.1983, 211.0316, 210.8867, 210.7729, 210.695, 210.6482, 
    210.6261, 210.6317, 210.645, 210.674, 210.6984, 210.7227, 210.7268, 
    210.7094,
  211.5823, 211.4055, 211.2207, 211.0634, 210.9369, 210.8416, 210.7883, 
    210.7534, 210.7461, 210.754, 210.7766, 210.8071, 210.8356, 210.8532, 
    210.8499,
  211.6181, 211.4767, 211.3054, 211.1425, 211.0044, 210.8998, 210.8421, 
    210.8007, 210.7898, 210.7865, 210.8058, 210.8375, 210.8775, 210.9095, 
    210.9296,
  211.7412, 211.6201, 211.4688, 211.2973, 211.1487, 211.025, 210.948, 
    210.8976, 210.8774, 210.8745, 210.8877, 210.9243, 210.965, 211.0065, 
    211.0329,
  211.7745, 211.6806, 211.5536, 211.392, 211.2496, 211.1051, 211.0051, 
    210.9421, 210.9166, 210.9091, 210.9197, 210.9488, 210.9997, 211.0453, 
    211.0829,
  211.8362, 211.7747, 211.6889, 211.5317, 211.3842, 211.2334, 211.107, 
    211.0153, 210.9682, 210.9557, 210.9593, 210.9836, 211.0291, 211.079, 
    211.1213,
  211.8243, 211.779, 211.728, 211.6356, 211.5232, 211.3438, 211.2019, 
    211.0649, 211.0002, 210.966, 210.9715, 210.9853, 211.027, 211.0713, 
    211.1167,
  211.8227, 211.7923, 211.773, 211.7379, 211.663, 211.4933, 211.3245, 
    211.1592, 211.0575, 210.9939, 210.9911, 211.0042, 211.0328, 211.0699, 
    211.11,
  211.7654, 211.7543, 211.7725, 211.7564, 211.7294, 211.6385, 211.4648, 
    211.2835, 211.1366, 211.0341, 211.004, 211.0094, 211.0293, 211.054, 
    211.0857,
  211.7387, 211.7156, 211.768, 211.8237, 211.838, 211.7757, 211.6066, 
    211.4267, 211.2827, 211.12, 211.0501, 211.0306, 211.0363, 211.0449, 
    211.0583,
  210.2235, 210.0802, 209.9276, 209.7639, 209.6133, 209.4789, 209.3636, 
    209.251, 209.1454, 209.0437, 208.9528, 208.8877, 208.8557, 208.8542, 
    208.8788,
  210.4155, 210.3182, 210.1614, 210.0067, 209.8395, 209.6906, 209.5707, 
    209.4601, 209.3647, 209.2657, 209.1684, 209.0823, 209.0152, 208.9798, 
    208.9866,
  210.4353, 210.3872, 210.2594, 210.1247, 209.9688, 209.8228, 209.6915, 
    209.5848, 209.4932, 209.406, 209.3186, 209.2281, 209.1467, 209.0864, 
    209.0587,
  210.487, 210.4635, 210.3635, 210.2417, 210.1076, 209.9698, 209.8483, 
    209.7386, 209.6577, 209.5857, 209.5082, 209.4222, 209.3294, 209.2492, 
    209.1942,
  210.4827, 210.4764, 210.423, 210.3139, 210.1954, 210.0699, 209.9612, 
    209.8526, 209.773, 209.71, 209.6512, 209.5742, 209.4856, 209.394, 209.3192,
  210.4896, 210.5096, 210.4869, 210.3963, 210.2807, 210.171, 210.0759, 
    209.9932, 209.9239, 209.8623, 209.8082, 209.74, 209.6616, 209.5644, 
    209.4756,
  210.4472, 210.4545, 210.4565, 210.4227, 210.3542, 210.2413, 210.1555, 
    210.0929, 210.0492, 209.9992, 209.9474, 209.8845, 209.812, 209.7212, 
    209.6206,
  210.433, 210.4332, 210.4444, 210.444, 210.4083, 210.332, 210.2616, 
    210.1977, 210.1615, 210.1352, 210.0889, 210.0459, 209.978, 209.8982, 
    209.7984,
  210.4389, 210.4273, 210.4205, 210.4107, 210.4222, 210.4053, 210.3436, 
    210.2943, 210.2512, 210.222, 210.2004, 210.1705, 210.1317, 210.0625, 
    209.974,
  210.5024, 210.4581, 210.4495, 210.4611, 210.4561, 210.4348, 210.3957, 
    210.3714, 210.3421, 210.2992, 210.2857, 210.2814, 210.2687, 210.2278, 
    210.1653,
  210.7937, 210.7904, 210.7838, 210.7623, 210.7331, 210.681, 210.6382, 
    210.5832, 210.5358, 210.4911, 210.4437, 210.3861, 210.3182, 210.2432, 
    210.1718,
  210.9023, 210.901, 210.9078, 210.9203, 210.9124, 210.8798, 210.8464, 
    210.7949, 210.7531, 210.6925, 210.6337, 210.5612, 210.4887, 210.4106, 
    210.3321,
  210.9752, 210.9516, 210.9678, 210.9719, 211.0008, 211.0112, 211.0061, 
    210.9689, 210.9401, 210.8718, 210.7983, 210.712, 210.6381, 210.5544, 
    210.4721,
  211.0959, 211.0526, 211.0481, 211.0456, 211.0633, 211.0818, 211.1228, 
    211.1337, 211.1324, 211.094, 211.0331, 210.9366, 210.8426, 210.7354, 
    210.6382,
  211.1673, 211.1086, 211.1167, 211.1022, 211.0962, 211.1026, 211.1429, 
    211.1775, 211.2191, 211.2193, 211.206, 211.1256, 211.0351, 210.9157, 
    210.7979,
  211.2934, 211.2391, 211.2263, 211.1969, 211.1514, 211.1437, 211.1699, 
    211.2076, 211.2718, 211.2933, 211.3171, 211.2856, 211.2229, 211.1229, 
    211.001,
  211.4115, 211.3315, 211.2951, 211.266, 211.2374, 211.1759, 211.1773, 
    211.208, 211.292, 211.358, 211.4087, 211.419, 211.3932, 211.3193, 211.2173,
  211.5634, 211.4702, 211.4184, 211.3751, 211.3414, 211.2717, 211.2234, 
    211.2254, 211.2976, 211.3983, 211.4807, 211.5263, 211.5384, 211.5061, 
    211.4277,
  211.7131, 211.6061, 211.5383, 211.4641, 211.4358, 211.3985, 211.3043, 
    211.2502, 211.2876, 211.3838, 211.514, 211.6, 211.6513, 211.66, 211.6035,
  211.8281, 211.7026, 211.6432, 211.6145, 211.5869, 211.5249, 211.434, 
    211.3436, 211.3237, 211.3626, 211.4915, 211.6188, 211.7167, 211.77, 
    211.7642,
  209.7754, 209.7545, 209.7491, 209.7337, 209.7122, 209.6618, 209.5919, 
    209.5095, 209.4382, 209.3972, 209.3845, 209.4068, 209.4551, 209.5326, 
    209.6355,
  209.8477, 209.8571, 209.849, 209.8371, 209.8095, 209.7661, 209.7138, 
    209.6428, 209.5841, 209.5374, 209.5244, 209.5272, 209.5668, 209.6174, 
    209.6931,
  209.835, 209.8534, 209.8738, 209.8996, 209.9126, 209.8952, 209.8674, 
    209.8102, 209.7484, 209.6731, 209.6158, 209.5938, 209.6066, 209.6584, 
    209.7319,
  209.8875, 209.864, 209.884, 209.9187, 209.9497, 209.9447, 209.9057, 
    209.835, 209.7524, 209.668, 209.6039, 209.5714, 209.5901, 209.6563, 
    209.7556,
  209.9649, 209.8954, 209.9014, 209.912, 209.9428, 209.9533, 209.9395, 
    209.9036, 209.8532, 209.7968, 209.7346, 209.6752, 209.6598, 209.7042, 
    209.7931,
  210.0566, 209.9811, 209.9569, 209.9354, 209.9598, 210.001, 210.0336, 
    210.0333, 209.987, 209.9038, 209.8028, 209.6949, 209.6351, 209.6425, 
    209.7168,
  210.1114, 210.0145, 209.956, 209.9303, 209.9307, 209.9444, 209.9849, 
    209.9986, 209.9975, 209.962, 209.9162, 209.8482, 209.782, 209.7377, 
    209.7442,
  210.114, 210.0388, 209.9754, 209.9514, 209.9267, 209.9427, 209.9962, 
    210.0277, 210.0528, 210.045, 210.0068, 209.9551, 209.8938, 209.8529, 
    209.8313,
  210.1753, 210.1199, 210.0396, 209.9625, 209.9395, 209.9539, 209.9879, 
    210.0169, 210.0349, 210.0173, 209.9782, 209.9082, 209.8465, 209.7988, 
    209.8015,
  210.2379, 210.1606, 210.0898, 210.0205, 209.9618, 209.9567, 209.9439, 
    209.979, 210.0232, 210.0262, 210.0086, 209.9431, 209.8753, 209.8271, 
    209.8158,
  211.1334, 211.0743, 211.0037, 210.9321, 210.8835, 210.8761, 210.9004, 
    210.9444, 211, 211.072, 211.1361, 211.1871, 211.2008, 211.1747, 211.1085,
  211.283, 211.2524, 211.1923, 211.1261, 211.0716, 211.0356, 211.0268, 
    211.0488, 211.0966, 211.1525, 211.2164, 211.273, 211.3205, 211.3334, 
    211.3162,
  211.3538, 211.3255, 211.2669, 211.1968, 211.1184, 211.0678, 211.0336, 
    211.033, 211.0616, 211.1048, 211.1639, 211.2323, 211.3042, 211.3468, 
    211.3432,
  211.3885, 211.3597, 211.2999, 211.2288, 211.157, 211.0882, 211.0293, 
    211.0051, 211.0067, 211.0349, 211.0812, 211.1468, 211.2316, 211.3065, 
    211.3387,
  211.4418, 211.4233, 211.401, 211.3396, 211.2774, 211.2108, 211.1531, 
    211.1163, 211.0876, 211.0822, 211.089, 211.1219, 211.1835, 211.2621, 
    211.3211,
  211.5475, 211.5321, 211.5318, 211.4741, 211.4198, 211.3781, 211.3398, 
    211.3015, 211.2538, 211.218, 211.1911, 211.1849, 211.1954, 211.2262, 
    211.2582,
  211.6141, 211.5615, 211.5419, 211.512, 211.4862, 211.4355, 211.4008, 
    211.369, 211.3308, 211.2931, 211.2485, 211.2169, 211.2014, 211.2178, 
    211.2515,
  211.6658, 211.6, 211.5672, 211.548, 211.5534, 211.5408, 211.5345, 211.5219, 
    211.4991, 211.4663, 211.4118, 211.3676, 211.3291, 211.3065, 211.3062,
  211.7055, 211.67, 211.6345, 211.6183, 211.6355, 211.6629, 211.6487, 
    211.6282, 211.5922, 211.5537, 211.5217, 211.4755, 211.4158, 211.3441, 
    211.3003,
  211.7825, 211.7251, 211.6939, 211.7124, 211.7242, 211.7389, 211.6924, 
    211.6696, 211.6654, 211.6197, 211.5938, 211.571, 211.5219, 211.4507, 
    211.3731,
  210.0608, 210.0841, 210.1019, 210.1115, 210.1114, 210.1099, 210.1114, 
    210.1132, 210.1217, 210.1376, 210.1621, 210.1993, 210.2407, 210.295, 
    210.3622,
  210.1124, 210.1108, 210.1222, 210.1425, 210.164, 210.1918, 210.2255, 
    210.2491, 210.2789, 210.3041, 210.3429, 210.3763, 210.4248, 210.4714, 
    210.5336,
  210.1503, 210.1346, 210.1424, 210.151, 210.1843, 210.2291, 210.2886, 
    210.3388, 210.3827, 210.4154, 210.4521, 210.4888, 210.5302, 210.5806, 
    210.6396,
  210.2261, 210.1887, 210.1831, 210.1927, 210.2421, 210.296, 210.3638, 
    210.4217, 210.4672, 210.4959, 210.5237, 210.5591, 210.5999, 210.652, 
    210.7163,
  210.3043, 210.237, 210.2246, 210.2339, 210.2853, 210.3359, 210.4014, 
    210.4476, 210.4941, 210.5229, 210.5495, 210.5864, 210.6405, 210.7072, 
    210.7876,
  210.457, 210.3739, 210.3515, 210.3135, 210.338, 210.3901, 210.4422, 
    210.4819, 210.5196, 210.5522, 210.5853, 210.6306, 210.7001, 210.7883, 
    210.8876,
  210.6117, 210.5107, 210.4523, 210.4156, 210.4342, 210.444, 210.4854, 
    210.5058, 210.5424, 210.5771, 210.6287, 210.6881, 210.7737, 210.8712, 
    210.9778,
  210.7368, 210.6698, 210.6105, 210.5644, 210.5444, 210.5078, 210.5302, 
    210.5595, 210.6005, 210.647, 210.6972, 210.7604, 210.8384, 210.9407, 
    211.0453,
  210.8177, 210.7954, 210.744, 210.6582, 210.6036, 210.5871, 210.5825, 
    210.6208, 210.6802, 210.7177, 210.7637, 210.8209, 210.8952, 210.984, 
    211.0807,
  210.8618, 210.855, 210.8186, 210.7531, 210.696, 210.6468, 210.6104, 
    210.6418, 210.7245, 210.7683, 210.8212, 210.8737, 210.9379, 211.0096, 
    211.0863,
  210.6008, 210.4997, 210.3842, 210.281, 210.1833, 210.0994, 210.0269, 
    209.9755, 209.9282, 209.8943, 209.868, 209.8595, 209.8625, 209.869, 
    209.8765,
  210.6837, 210.5751, 210.4481, 210.3344, 210.2327, 210.1445, 210.0694, 
    210.0023, 209.9511, 209.9098, 209.8904, 209.8817, 209.8865, 209.8908, 
    209.8984,
  210.6938, 210.5851, 210.4722, 210.3553, 210.2388, 210.1372, 210.0594, 
    209.9892, 209.9417, 209.9058, 209.8901, 209.8813, 209.8772, 209.8668, 
    209.8555,
  210.7373, 210.6368, 210.5419, 210.4231, 210.3047, 210.194, 210.1053, 
    210.0304, 209.9774, 209.9447, 209.9292, 209.9187, 209.9028, 209.8786, 
    209.8471,
  210.7639, 210.655, 210.5675, 210.4532, 210.348, 210.237, 210.1376, 
    210.0621, 209.9987, 209.9557, 209.9324, 209.9161, 209.8921, 209.8567, 
    209.8144,
  210.8189, 210.7229, 210.6469, 210.5212, 210.4033, 210.2978, 210.2032, 
    210.1199, 210.0544, 209.9975, 209.9513, 209.923, 209.8994, 209.8711, 
    209.829,
  210.8348, 210.7439, 210.674, 210.5724, 210.4689, 210.3356, 210.2358, 
    210.1444, 210.0792, 210.0104, 209.9484, 209.9045, 209.8745, 209.859, 
    209.8359,
  210.858, 210.7797, 210.7219, 210.652, 210.5553, 210.4154, 210.2916, 
    210.1881, 210.1112, 210.0503, 209.982, 209.9265, 209.8805, 209.8569, 
    209.8431,
  210.8607, 210.8163, 210.7598, 210.672, 210.5884, 210.5, 210.3715, 210.2468, 
    210.1518, 210.0723, 210.0215, 209.9554, 209.9072, 209.8696, 209.8588,
  210.8706, 210.8348, 210.8195, 210.7663, 210.6884, 210.5803, 210.4481, 
    210.3299, 210.2519, 210.1458, 210.0744, 210.0082, 209.9415, 209.9055, 
    209.878,
  209.0869, 209.1237, 209.1592, 209.1554, 209.1498, 209.1163, 209.0668, 
    208.9918, 208.9215, 208.8432, 208.7741, 208.7101, 208.6599, 208.6189, 
    208.6092,
  209.0834, 209.1241, 209.1602, 209.1677, 209.1727, 209.1498, 209.1224, 
    209.0699, 209.0254, 208.9641, 208.9073, 208.8308, 208.7686, 208.7143, 
    208.6819,
  209.1047, 209.1646, 209.2142, 209.2379, 209.2422, 209.215, 209.1796, 
    209.1329, 209.0914, 209.0476, 208.9909, 208.9252, 208.8464, 208.7782, 
    208.7314,
  209.1303, 209.2098, 209.2854, 209.3389, 209.3626, 209.339, 209.3027, 
    209.2443, 209.2092, 209.1631, 209.1144, 209.0364, 208.958, 208.8767, 
    208.8173,
  209.1457, 209.2183, 209.3251, 209.3997, 209.4463, 209.438, 209.4039, 
    209.3611, 209.3205, 209.2752, 209.2187, 209.1435, 209.063, 208.9798, 
    208.9062,
  209.1748, 209.2522, 209.3586, 209.4275, 209.4716, 209.4957, 209.4998, 
    209.48, 209.4519, 209.3992, 209.3248, 209.2383, 209.1592, 209.0893, 
    209.0299,
  209.2085, 209.2536, 209.3287, 209.4101, 209.4935, 209.53, 209.5665, 
    209.5788, 209.5718, 209.4979, 209.4092, 209.3167, 209.2493, 209.2031, 
    209.1548,
  209.2452, 209.2708, 209.3358, 209.4305, 209.5164, 209.5735, 209.6318, 
    209.6497, 209.6441, 209.5825, 209.4935, 209.4173, 209.3551, 209.3068, 
    209.2607,
  209.2611, 209.2816, 209.3446, 209.4056, 209.5116, 209.6315, 209.6882, 
    209.6912, 209.6645, 209.621, 209.5749, 209.5231, 209.4655, 209.4088, 
    209.3594,
  209.2941, 209.2747, 209.343, 209.4474, 209.5615, 209.6735, 209.7011, 
    209.6934, 209.7056, 209.6719, 209.6906, 209.6682, 209.601, 209.5258, 
    209.4564,
  210.5184, 210.3878, 210.2761, 210.1735, 210.0897, 210.0072, 209.927, 
    209.8311, 209.7413, 209.6636, 209.6154, 209.585, 209.5701, 209.5511, 
    209.5394,
  210.6889, 210.5635, 210.4533, 210.3465, 210.2529, 210.1584, 210.0732, 
    209.9751, 209.8906, 209.8145, 209.7709, 209.7391, 209.7209, 209.7002, 
    209.6681,
  210.7519, 210.6473, 210.5456, 210.4386, 210.3441, 210.2461, 210.154, 
    210.0565, 209.9721, 209.9028, 209.8687, 209.846, 209.829, 209.8005, 
    209.7545,
  210.8772, 210.7798, 210.676, 210.5753, 210.4822, 210.3699, 210.268, 
    210.1615, 210.0797, 210.0087, 209.9747, 209.9513, 209.9364, 209.9042, 
    209.8532,
  210.955, 210.8512, 210.7713, 210.6756, 210.5873, 210.4685, 210.3537, 
    210.2348, 210.1603, 210.0984, 210.0565, 210.0257, 209.9959, 209.9662, 
    209.92,
  211.0584, 210.9682, 210.9085, 210.8005, 210.7039, 210.5989, 210.4891, 
    210.3629, 210.2793, 210.2158, 210.1642, 210.1101, 210.0726, 210.0312, 
    209.9935,
  211.0853, 210.9993, 210.9344, 210.8704, 210.8219, 210.7043, 210.6073, 
    210.4982, 210.409, 210.3406, 210.2661, 210.199, 210.1391, 210.1056, 
    210.0885,
  211.1088, 211.035, 210.9847, 210.9366, 210.9046, 210.807, 210.7316, 
    210.6453, 210.5614, 210.4897, 210.4067, 210.3327, 210.2704, 210.2339, 
    210.2193,
  211.0981, 211.0393, 211.0129, 210.9368, 210.9064, 210.8871, 210.8133, 
    210.7385, 210.6675, 210.5971, 210.5605, 210.5157, 210.4745, 210.4294, 
    210.396,
  211.0887, 211.0396, 211.0354, 211.0064, 210.9824, 210.949, 210.8585, 
    210.7811, 210.7518, 210.6827, 210.6665, 210.6543, 210.616, 210.5677, 
    210.5201,
  210.0333, 210.0199, 210.0155, 209.9925, 209.9605, 209.8988, 209.8339, 
    209.7557, 209.6826, 209.6143, 209.555, 209.488, 209.4121, 209.3262, 
    209.245,
  210.1364, 210.0978, 210.0876, 210.0688, 210.0452, 209.9988, 209.9471, 
    209.876, 209.8106, 209.7474, 209.6953, 209.6322, 209.5547, 209.4637, 
    209.3755,
  210.1785, 210.1406, 210.1325, 210.1031, 210.0819, 210.0439, 210.0003, 
    209.9429, 209.8829, 209.8282, 209.7759, 209.7208, 209.6508, 209.5706, 
    209.4957,
  210.2843, 210.2449, 210.2202, 210.1826, 210.1644, 210.1259, 210.0845, 
    210.0271, 209.9699, 209.9099, 209.86, 209.8069, 209.7558, 209.6976, 
    209.6514,
  210.3683, 210.3169, 210.2986, 210.266, 210.2401, 210.1978, 210.1536, 
    210.0846, 210.024, 209.9632, 209.917, 209.8751, 209.8416, 209.8113, 
    209.7867,
  210.4801, 210.4381, 210.4095, 210.3509, 210.3204, 210.2883, 210.2386, 
    210.164, 210.0939, 210.0312, 209.9868, 209.9545, 209.9356, 209.9206, 
    209.9132,
  210.585, 210.5203, 210.4748, 210.4324, 210.4158, 210.3735, 210.3128, 
    210.2308, 210.157, 210.0934, 210.0521, 210.0237, 210.0138, 210.0064, 
    210.0065,
  210.6313, 210.5807, 210.5527, 210.5207, 210.4979, 210.4348, 210.382, 
    210.2963, 210.2229, 210.1571, 210.1208, 210.0996, 210.0895, 210.0864, 
    210.0917,
  210.6574, 210.629, 210.6154, 210.5526, 210.5346, 210.5237, 210.4587, 
    210.3725, 210.2941, 210.2171, 210.1831, 210.1631, 210.1571, 210.1521, 
    210.1614,
  210.6498, 210.6188, 210.6315, 210.6233, 210.6228, 210.6038, 210.509, 
    210.429, 210.3829, 210.2829, 210.2447, 210.2155, 210.203, 210.2006, 
    210.2158,
  210.0448, 210.0048, 209.9683, 209.9151, 209.8609, 209.7825, 209.7066, 
    209.6194, 209.531, 209.4558, 209.3923, 209.3379, 209.2912, 209.2459, 
    209.2067,
  210.1775, 210.1205, 210.0753, 210.028, 209.983, 209.918, 209.8515, 209.765, 
    209.6736, 209.585, 209.5109, 209.4521, 209.4082, 209.3716, 209.3374,
  210.2234, 210.1606, 210.1232, 210.0813, 210.0393, 209.9877, 209.933, 
    209.8589, 209.7788, 209.6932, 209.6218, 209.5575, 209.5157, 209.4825, 
    209.4502,
  210.3148, 210.2579, 210.2105, 210.1563, 210.1194, 210.0902, 210.0609, 
    210.0157, 209.9544, 209.8763, 209.7959, 209.7258, 209.6651, 209.6105, 
    209.5706,
  210.3891, 210.3301, 210.2722, 210.2127, 210.1833, 210.1634, 210.1545, 
    210.1326, 210.1034, 210.0454, 209.9703, 209.8831, 209.8036, 209.7208, 
    209.6486,
  210.4769, 210.4215, 210.3777, 210.3205, 210.2857, 210.2817, 210.2851, 
    210.2707, 210.2622, 210.2203, 210.151, 210.0513, 209.9447, 209.8318, 
    209.7251,
  210.521, 210.4666, 210.4215, 210.3883, 210.3799, 210.3754, 210.378, 
    210.3708, 210.3581, 210.3257, 210.2609, 210.1641, 210.0456, 209.9196, 
    209.7983,
  210.5478, 210.5119, 210.4741, 210.4556, 210.4565, 210.4527, 210.4501, 
    210.4304, 210.4133, 210.374, 210.3157, 210.2308, 210.1192, 210.0032, 
    209.8936,
  210.5568, 210.5337, 210.5112, 210.469, 210.4675, 210.4836, 210.4597, 
    210.4417, 210.4142, 210.3702, 210.3241, 210.2664, 210.1882, 210.1054, 
    210.0314,
  210.5477, 210.5175, 210.517, 210.5181, 210.5147, 210.4891, 210.4267, 
    210.3907, 210.3981, 210.3558, 210.3468, 210.3256, 210.2968, 210.2542, 
    210.2222,
  208.4109, 208.3725, 208.3445, 208.3167, 208.3026, 208.2756, 208.2484, 
    208.1944, 208.1369, 208.0719, 208.0225, 207.9827, 207.9601, 207.9524, 
    207.9719,
  208.5381, 208.4956, 208.4422, 208.4085, 208.3862, 208.3517, 208.3401, 
    208.302, 208.2665, 208.2166, 208.1735, 208.1362, 208.1088, 208.0956, 
    208.1019,
  208.6303, 208.5814, 208.541, 208.496, 208.4534, 208.4144, 208.3971, 
    208.3717, 208.3528, 208.321, 208.2946, 208.267, 208.2518, 208.241, 
    208.2456,
  208.7312, 208.7036, 208.6586, 208.6014, 208.547, 208.5047, 208.4831, 
    208.4697, 208.4717, 208.4574, 208.4461, 208.4234, 208.4045, 208.387, 
    208.3824,
  208.8532, 208.8203, 208.7705, 208.7086, 208.6524, 208.6061, 208.5722, 
    208.5549, 208.569, 208.5706, 208.569, 208.5545, 208.5384, 208.5239, 
    208.5158,
  208.961, 208.9341, 208.8993, 208.8345, 208.7734, 208.7208, 208.6909, 
    208.6717, 208.6821, 208.6938, 208.7039, 208.6883, 208.6689, 208.6482, 
    208.6438,
  209.0189, 209.0157, 209.0042, 208.9618, 208.9232, 208.8641, 208.8155, 
    208.7861, 208.7903, 208.798, 208.8047, 208.7894, 208.7749, 208.7662, 
    208.772,
  209.0837, 209.1017, 209.1133, 209.1048, 209.0905, 209.0441, 208.9889, 
    208.9283, 208.8925, 208.8868, 208.8725, 208.8654, 208.853, 208.8686, 
    208.8944,
  209.1673, 209.1779, 209.2023, 209.2002, 209.2129, 209.1988, 209.1506, 
    209.0975, 209.0385, 208.9918, 208.9615, 208.9435, 208.934, 208.9571, 
    209.0201,
  209.2495, 209.2432, 209.2894, 209.3356, 209.3619, 209.3466, 209.2961, 
    209.2451, 209.2078, 209.1308, 209.0806, 209.0448, 209.0392, 209.0766, 
    209.1518,
  209.7347, 209.7312, 209.7389, 209.7567, 209.7536, 209.7284, 209.6894, 
    209.6329, 209.5671, 209.482, 209.3939, 209.3058, 209.2161, 209.1206, 
    209.0396,
  209.9127, 209.899, 209.8847, 209.9025, 209.9119, 209.8975, 209.8668, 
    209.8189, 209.759, 209.6788, 209.5829, 209.4786, 209.3723, 209.2605, 
    209.1648,
  209.9962, 209.9892, 209.9837, 209.9849, 209.9857, 209.9773, 209.965, 
    209.9388, 209.9048, 209.8464, 209.7657, 209.6562, 209.5295, 209.3884, 
    209.2622,
  210.158, 210.1496, 210.1495, 210.1322, 210.1311, 210.1211, 210.1137, 
    210.0972, 210.0824, 210.0394, 209.9619, 209.8428, 209.6988, 209.537, 
    209.3818,
  210.28, 210.2771, 210.2841, 210.2643, 210.2455, 210.2281, 210.2172, 
    210.2157, 210.2118, 210.1934, 210.1269, 210.0064, 209.8484, 209.6743, 
    209.5022,
  210.3896, 210.3933, 210.4166, 210.4057, 210.3825, 210.3741, 210.3622, 
    210.3478, 210.3574, 210.3557, 210.3058, 210.1877, 210.0211, 209.8373, 
    209.6616,
  210.4599, 210.4626, 210.488, 210.5041, 210.5118, 210.4944, 210.4759, 
    210.4703, 210.4742, 210.4836, 210.4494, 210.3515, 210.1864, 210.0081, 
    209.8356,
  210.5462, 210.5319, 210.5755, 210.605, 210.634, 210.6301, 210.6144, 
    210.5971, 210.5952, 210.5963, 210.5723, 210.4992, 210.3608, 210.1906, 
    210.0376,
  210.6223, 210.5843, 210.6155, 210.64, 210.6975, 210.7301, 210.7125, 
    210.7067, 210.7149, 210.713, 210.6891, 210.6244, 210.502, 210.3515, 
    210.2159,
  210.7067, 210.6615, 210.6748, 210.7329, 210.7962, 210.8199, 210.8088, 
    210.8057, 210.8384, 210.8333, 210.8113, 210.7619, 210.6638, 210.5445, 
    210.4264,
  208.5279, 208.4546, 208.3867, 208.3074, 208.2478, 208.1978, 208.1748, 
    208.1815, 208.2229, 208.2757, 208.3309, 208.409, 208.4782, 208.5416, 
    208.6128,
  208.6114, 208.5409, 208.4663, 208.4019, 208.3409, 208.2847, 208.2434, 
    208.2228, 208.2384, 208.2723, 208.3188, 208.3846, 208.4516, 208.5243, 
    208.6025,
  208.6551, 208.5987, 208.5494, 208.5031, 208.4464, 208.3922, 208.3442, 
    208.3061, 208.2901, 208.3037, 208.3327, 208.3832, 208.4424, 208.5216, 
    208.5941,
  208.7237, 208.6806, 208.6378, 208.6004, 208.5609, 208.5199, 208.4731, 
    208.4262, 208.3942, 208.3744, 208.3805, 208.4066, 208.4547, 208.5148, 
    208.5899,
  208.7948, 208.7455, 208.7115, 208.6871, 208.6623, 208.626, 208.5855, 
    208.5401, 208.4941, 208.4602, 208.4422, 208.4422, 208.465, 208.5104, 
    208.5708,
  208.8597, 208.8075, 208.7797, 208.7503, 208.7233, 208.7078, 208.6654, 
    208.621, 208.5771, 208.5449, 208.5124, 208.4981, 208.4946, 208.5182, 
    208.5657,
  208.9101, 208.8477, 208.8135, 208.7953, 208.7906, 208.7628, 208.7181, 
    208.6669, 208.628, 208.6019, 208.5756, 208.5567, 208.5388, 208.5476, 
    208.5769,
  208.9302, 208.8776, 208.8608, 208.8479, 208.8367, 208.803, 208.7603, 
    208.712, 208.6794, 208.6691, 208.6553, 208.6478, 208.6354, 208.6405, 
    208.6561,
  208.9484, 208.9116, 208.8826, 208.8508, 208.8495, 208.8328, 208.7772, 
    208.7494, 208.728, 208.7389, 208.7538, 208.7559, 208.75, 208.7513, 
    208.7657,
  208.9554, 208.9208, 208.9091, 208.9193, 208.9037, 208.8465, 208.7867, 
    208.7643, 208.7918, 208.8098, 208.847, 208.8589, 208.8596, 208.8661, 
    208.8911,
  209.6455, 209.7554, 209.8301, 209.8818, 209.8977, 209.8772, 209.8365, 
    209.7778, 209.7236, 209.673, 209.6316, 209.5931, 209.5567, 209.5171, 
    209.4817,
  209.5779, 209.6938, 209.7974, 209.8975, 209.9455, 209.9451, 209.9164, 
    209.8614, 209.8016, 209.7439, 209.6913, 209.65, 209.6164, 209.5777, 
    209.5392,
  209.4799, 209.5874, 209.723, 209.8448, 209.933, 209.9614, 209.9463, 
    209.902, 209.8315, 209.7711, 209.7108, 209.6619, 209.6216, 209.5834, 
    209.5496,
  209.4482, 209.5283, 209.6599, 209.7933, 209.915, 209.9876, 209.9929, 
    209.9583, 209.8943, 209.8174, 209.7492, 209.6873, 209.6432, 209.5991, 
    209.5616,
  209.4599, 209.4795, 209.5902, 209.7218, 209.8597, 209.952, 209.9921, 
    209.972, 209.9259, 209.847, 209.7697, 209.6965, 209.6405, 209.5968, 
    209.5559,
  209.5197, 209.5022, 209.574, 209.6653, 209.784, 209.8979, 209.9673, 
    209.9821, 209.9582, 209.9008, 209.8223, 209.7424, 209.6764, 209.6212, 
    209.571,
  209.6194, 209.5639, 209.5695, 209.6376, 209.7487, 209.832, 209.9019, 
    209.9382, 209.9545, 209.928, 209.8756, 209.8009, 209.7256, 209.664, 
    209.5997,
  209.7585, 209.6874, 209.6634, 209.6798, 209.7467, 209.8087, 209.8614, 
    209.9031, 209.9353, 209.9536, 209.9295, 209.8834, 209.8166, 209.7571, 
    209.6918,
  209.8696, 209.8373, 209.7941, 209.7415, 209.7603, 209.8173, 209.8401, 
    209.8781, 209.9234, 209.9559, 209.9677, 209.9347, 209.8831, 209.8272, 
    209.7662,
  209.9785, 209.9583, 209.9386, 209.9132, 209.8786, 209.8431, 209.8358, 
    209.8752, 209.9468, 209.9799, 210.0008, 209.9841, 209.927, 209.8703, 
    209.8101,
  208.843, 208.805, 208.7932, 208.7811, 208.7717, 208.7698, 208.7594, 
    208.7247, 208.6816, 208.6183, 208.556, 208.4947, 208.4494, 208.419, 
    208.4084,
  208.8706, 208.8346, 208.7991, 208.7801, 208.7737, 208.7788, 208.7767, 
    208.7629, 208.7325, 208.6801, 208.6229, 208.5618, 208.5113, 208.4798, 
    208.4703,
  208.8656, 208.8253, 208.7927, 208.7685, 208.7589, 208.7628, 208.7638, 
    208.7579, 208.7404, 208.6995, 208.649, 208.5916, 208.5395, 208.4991, 
    208.4866,
  208.9132, 208.8778, 208.8301, 208.7929, 208.7735, 208.7667, 208.7707, 
    208.7686, 208.767, 208.7388, 208.7003, 208.6461, 208.5843, 208.5355, 
    208.5059,
  208.9495, 208.915, 208.8681, 208.8248, 208.7927, 208.7671, 208.7583, 
    208.7553, 208.7569, 208.7472, 208.7203, 208.6854, 208.6324, 208.5816, 
    208.5447,
  208.9875, 208.9606, 208.921, 208.862, 208.8066, 208.7864, 208.7673, 
    208.7523, 208.7474, 208.7466, 208.7375, 208.7198, 208.6935, 208.654, 
    208.6165,
  209.0188, 208.9716, 208.9254, 208.9002, 208.8621, 208.8114, 208.7682, 
    208.745, 208.7427, 208.7447, 208.751, 208.7515, 208.7438, 208.7326, 
    208.7079,
  209.0657, 209.0053, 208.9677, 208.9504, 208.9172, 208.8648, 208.8109, 
    208.7578, 208.7428, 208.749, 208.764, 208.7856, 208.7967, 208.8055, 
    208.7934,
  209.1073, 209.0569, 209.0155, 208.9654, 208.9544, 208.9554, 208.8685, 
    208.8009, 208.7549, 208.7486, 208.7866, 208.821, 208.8472, 208.8559, 
    208.8488,
  209.1862, 209.1155, 209.0779, 209.0782, 209.08, 209.0064, 208.9173, 
    208.8554, 208.8191, 208.7842, 208.8121, 208.8569, 208.8914, 208.9081, 
    208.9069,
  208.7432, 208.6768, 208.6702, 208.7334, 208.8345, 208.9441, 209.047, 
    209.1105, 209.134, 209.0924, 209.0129, 208.9051, 208.7781, 208.6506, 
    208.5366,
  208.9053, 208.7998, 208.7458, 208.7776, 208.8605, 208.9751, 209.09, 
    209.1717, 209.2087, 209.1853, 209.112, 209.0131, 208.8972, 208.7763, 
    208.6588,
  209.0354, 208.8948, 208.8253, 208.8152, 208.8629, 208.969, 209.0851, 
    209.1793, 209.2287, 209.2239, 209.1686, 209.0721, 208.9618, 208.8458, 
    208.7332,
  209.1725, 209.0431, 208.9428, 208.8878, 208.8976, 208.9626, 209.0665, 
    209.1597, 209.238, 209.2556, 209.2326, 209.1492, 209.0568, 208.9398, 
    208.8285,
  209.2836, 209.1749, 209.072, 208.9862, 208.9555, 208.9695, 209.0306, 
    209.1211, 209.2146, 209.2702, 209.2816, 209.2286, 209.1519, 209.0424, 
    208.9299,
  209.3772, 209.3026, 209.2088, 209.11, 209.0358, 209.0192, 209.0498, 
    209.1086, 209.2139, 209.3033, 209.3557, 209.3495, 209.2805, 209.1816, 
    209.0642,
  209.4328, 209.384, 209.3082, 209.2231, 209.1626, 209.0853, 209.0895, 
    209.1352, 209.2365, 209.3522, 209.4418, 209.4665, 209.4203, 209.3221, 
    209.1996,
  209.4729, 209.4581, 209.4282, 209.369, 209.3021, 209.2015, 209.1682, 
    209.1874, 209.2902, 209.4144, 209.5387, 209.5887, 209.5585, 209.464, 
    209.3192,
  209.4659, 209.5047, 209.5186, 209.4745, 209.4257, 209.3417, 209.2488, 
    209.249, 209.3258, 209.4465, 209.5941, 209.6738, 209.6723, 209.5909, 
    209.4468,
  209.478, 209.5356, 209.5932, 209.6189, 209.5849, 209.4495, 209.3262, 
    209.289, 209.3575, 209.4551, 209.5966, 209.7021, 209.7214, 209.6738, 
    209.5542,
  208.7999, 208.8511, 208.9218, 208.9946, 209.0516, 209.0731, 209.0618, 
    209.0186, 208.9785, 208.9372, 208.8993, 208.8474, 208.774, 208.6881, 
    208.5939,
  208.8393, 208.8733, 208.9312, 209.0135, 209.0833, 209.1349, 209.1543, 
    209.1377, 209.1098, 209.0755, 209.041, 208.989, 208.9197, 208.8371, 
    208.7526,
  208.8699, 208.8777, 208.9209, 208.991, 209.0603, 209.1191, 209.157, 
    209.1839, 209.1985, 209.2051, 209.1903, 209.1448, 209.0687, 208.9828, 
    208.9036,
  208.93, 208.9104, 208.9324, 208.9846, 209.0517, 209.1198, 209.1665, 
    209.2227, 209.2761, 209.3286, 209.3419, 209.3048, 209.2288, 209.1389, 
    209.0611,
  209.0108, 208.9531, 208.9512, 208.9861, 209.0449, 209.1076, 209.1595, 
    209.2293, 209.3065, 209.3913, 209.4296, 209.4144, 209.3462, 209.2669, 
    209.188,
  209.1147, 209.0337, 209.0084, 209.0104, 209.0458, 209.1164, 209.1744, 
    209.2447, 209.3339, 209.4369, 209.4973, 209.4993, 209.4479, 209.3783, 
    209.3052,
  209.2101, 209.1051, 209.0517, 209.0362, 209.0716, 209.1111, 209.1778, 
    209.2478, 209.3444, 209.4436, 209.525, 209.548, 209.5299, 209.4787, 
    209.4167,
  209.318, 209.2127, 209.1439, 209.1131, 209.1228, 209.1444, 209.1912, 
    209.2575, 209.3406, 209.442, 209.5347, 209.5863, 209.601, 209.5764, 
    209.5314,
  209.4275, 209.3437, 209.2588, 209.1798, 209.1657, 209.2014, 209.2149, 
    209.2668, 209.3247, 209.4106, 209.5172, 209.595, 209.6523, 209.6577, 
    209.6416,
  209.5304, 209.4617, 209.4056, 209.3454, 209.3061, 209.2573, 209.235, 
    209.2617, 209.3269, 209.379, 209.4896, 209.5925, 209.682, 209.7195, 
    209.7302,
  209.9283, 209.7984, 209.6933, 209.5796, 209.5145, 209.4524, 209.4242, 
    209.4016, 209.3959, 209.4011, 209.4241, 209.4318, 209.4274, 209.4057, 
    209.3589,
  210.1331, 209.9477, 209.8164, 209.6812, 209.5921, 209.5085, 209.4743, 
    209.46, 209.4669, 209.4878, 209.5131, 209.5404, 209.5445, 209.5328, 
    209.4897,
  210.2639, 210.0826, 209.94, 209.7839, 209.6626, 209.5568, 209.5018, 
    209.4835, 209.4916, 209.5183, 209.5444, 209.5767, 209.6004, 209.6004, 
    209.5858,
  210.4388, 210.2651, 210.1153, 209.928, 209.78, 209.6495, 209.568, 209.5264, 
    209.5218, 209.5325, 209.5547, 209.5849, 209.6178, 209.6425, 209.6476,
  210.5963, 210.4317, 210.2863, 210.086, 209.9165, 209.7464, 209.6331, 
    209.5506, 209.5326, 209.5288, 209.5463, 209.574, 209.619, 209.6553, 
    209.6897,
  210.7207, 210.5999, 210.4737, 210.274, 210.0859, 209.8923, 209.7476, 
    209.6268, 209.5659, 209.5442, 209.5452, 209.5746, 209.6297, 209.6939, 
    209.7432,
  210.8059, 210.7231, 210.6132, 210.452, 210.2934, 210.0789, 209.9048, 
    209.7478, 209.6416, 209.5866, 209.5701, 209.5939, 209.6406, 209.7128, 
    209.771,
  210.8652, 210.8215, 210.7579, 210.6315, 210.4967, 210.2972, 210.104, 
    209.915, 209.7791, 209.6747, 209.6317, 209.6284, 209.653, 209.7231, 
    209.8032,
  210.9022, 210.8726, 210.8548, 210.7417, 210.6489, 210.5066, 210.318, 
    210.1087, 209.9383, 209.8028, 209.7215, 209.6861, 209.6969, 209.7334, 
    209.7986,
  210.9427, 210.9129, 210.9238, 210.8995, 210.8196, 210.6829, 210.5012, 
    210.3174, 210.1309, 209.9716, 209.8568, 209.7938, 209.7586, 209.7645, 
    209.8188,
  208.5519, 208.4683, 208.3588, 208.2676, 208.1826, 208.0803, 207.9818, 
    207.8838, 207.803, 207.7426, 207.7054, 207.6864, 207.6882, 207.6952, 
    207.7122,
  208.6183, 208.5375, 208.4319, 208.3576, 208.2804, 208.1814, 208.0784, 
    207.9621, 207.8648, 207.7834, 207.7352, 207.7086, 207.7023, 207.7103, 
    207.7316,
  208.631, 208.5414, 208.4674, 208.4057, 208.3307, 208.2457, 208.1444, 
    208.026, 207.922, 207.8336, 207.779, 207.7492, 207.741, 207.747, 207.7635,
  208.6812, 208.592, 208.5206, 208.446, 208.3802, 208.3043, 208.2077, 
    208.0976, 208.0034, 207.9209, 207.8673, 207.8304, 207.8149, 207.8049, 
    207.8077,
  208.7365, 208.6313, 208.5522, 208.4838, 208.43, 208.3579, 208.2665, 
    208.1668, 208.0788, 208.0077, 207.9506, 207.9085, 207.8802, 207.8602, 
    207.8503,
  208.7959, 208.6871, 208.602, 208.5218, 208.4473, 208.4047, 208.3258, 
    208.2404, 208.1583, 208.0922, 208.0323, 207.9776, 207.9367, 207.9112, 
    207.8885,
  208.8523, 208.7345, 208.6185, 208.5405, 208.4908, 208.4433, 208.3765, 
    208.3079, 208.2247, 208.1546, 208.0794, 208.0165, 207.9607, 207.9295, 
    207.9015,
  208.9065, 208.7928, 208.6765, 208.5973, 208.5452, 208.484, 208.436, 
    208.3682, 208.2901, 208.2138, 208.1334, 208.0636, 208.0052, 207.9658, 
    207.9362,
  208.9634, 208.8526, 208.734, 208.6295, 208.5726, 208.5441, 208.4866, 
    208.4221, 208.3515, 208.2722, 208.2024, 208.1277, 208.0568, 207.9912, 
    207.9386,
  209.0224, 208.8971, 208.7927, 208.7232, 208.6666, 208.5997, 208.5225, 
    208.4643, 208.4143, 208.3376, 208.2674, 208.1879, 208.0997, 208.0238, 
    207.9854,
  208.2579, 208.1358, 208.0346, 207.9325, 207.8561, 207.788, 207.7303, 
    207.667, 207.6012, 207.5335, 207.467, 207.4149, 207.3682, 207.3341, 
    207.3099,
  208.4834, 208.3485, 208.2185, 208.0957, 208.0161, 207.9455, 207.8994, 
    207.842, 207.7865, 207.7168, 207.6465, 207.5776, 207.5214, 207.4802, 
    207.451,
  208.6344, 208.5211, 208.4032, 208.2759, 208.171, 208.093, 208.052, 
    207.9986, 207.9522, 207.8886, 207.8226, 207.7521, 207.6856, 207.6329, 
    207.5902,
  208.7942, 208.7177, 208.6168, 208.4693, 208.3495, 208.2584, 208.2041, 
    208.1525, 208.1099, 208.054, 207.9912, 207.9169, 207.8465, 207.7888, 
    207.739,
  208.9443, 208.895, 208.8129, 208.6644, 208.5356, 208.4222, 208.3575, 
    208.3069, 208.2626, 208.2063, 208.1412, 208.0616, 207.9895, 207.9247, 
    207.8772,
  209.0437, 209.0392, 208.9952, 208.8542, 208.7064, 208.5928, 208.5191, 
    208.4639, 208.4261, 208.3676, 208.3008, 208.2089, 208.1296, 208.0607, 
    208.0143,
  209.0913, 209.124, 209.1087, 209.0043, 208.8887, 208.75, 208.6593, 
    208.6036, 208.574, 208.5272, 208.4597, 208.3701, 208.2794, 208.2057, 
    208.1513,
  209.1077, 209.1756, 209.2093, 209.1495, 209.0479, 208.9108, 208.8041, 
    208.7324, 208.7022, 208.6732, 208.6211, 208.5433, 208.4479, 208.3594, 
    208.2936,
  209.1222, 209.2065, 209.2776, 209.2308, 209.1657, 209.0651, 208.935, 
    208.8438, 208.8103, 208.7916, 208.778, 208.7178, 208.6344, 208.5383, 
    208.4518,
  209.167, 209.2143, 209.3096, 209.3528, 209.3306, 209.2001, 209.0595, 
    208.9521, 208.9026, 208.8797, 208.8829, 208.8634, 208.799, 208.7106, 
    208.6192,
  209.0182, 209.0437, 209.0575, 209.0617, 209.0318, 208.9846, 208.9409, 
    208.8918, 208.83, 208.7649, 208.6865, 208.613, 208.5353, 208.4621, 
    208.4033,
  209.0658, 209.1102, 209.133, 209.1545, 209.1396, 209.1119, 209.0675, 
    209.0061, 208.9422, 208.879, 208.8141, 208.748, 208.683, 208.6176, 
    208.5547,
  209.0473, 209.125, 209.1881, 209.233, 209.2208, 209.2111, 209.1772, 
    209.1278, 209.0749, 209.016, 208.9526, 208.887, 208.8237, 208.7605, 
    208.6976,
  209.0069, 209.1145, 209.2203, 209.2855, 209.3035, 209.3206, 209.296, 
    209.255, 209.2088, 209.1438, 209.0845, 209.0226, 208.9608, 208.8964, 
    208.8321,
  208.9726, 209.0797, 209.2067, 209.3039, 209.368, 209.4106, 209.4031, 
    209.3759, 209.3395, 209.2781, 209.2195, 209.1593, 209.0977, 209.0314, 
    208.9622,
  208.9433, 209.0414, 209.1725, 209.288, 209.3688, 209.4575, 209.4908, 
    209.4861, 209.4623, 209.4175, 209.3631, 209.304, 209.2452, 209.1781, 
    209.0994,
  208.9213, 208.9683, 209.0716, 209.2018, 209.3404, 209.4543, 209.5268, 
    209.5607, 209.5614, 209.5313, 209.4863, 209.433, 209.3825, 209.3207, 
    209.2462,
  208.9291, 208.9373, 208.996, 209.1306, 209.2715, 209.4103, 209.5255, 
    209.5837, 209.6123, 209.6085, 209.5841, 209.5501, 209.5122, 209.4683, 
    209.4051,
  208.9867, 208.9547, 208.9789, 209.0277, 209.1705, 209.3543, 209.4804, 
    209.558, 209.606, 209.6291, 209.638, 209.6256, 209.6084, 209.5846, 
    209.5469,
  209.0842, 209.0168, 208.995, 209.0461, 209.1873, 209.2917, 209.4149, 
    209.5222, 209.5909, 209.6221, 209.6449, 209.6614, 209.6523, 209.6657, 
    209.6582,
  209.9812, 209.9422, 209.9396, 209.9827, 210.017, 210.063, 210.081, 
    210.0696, 210.0367, 209.9905, 209.9341, 209.8759, 209.8159, 209.7736, 
    209.7412,
  210.1104, 210.0549, 210.0203, 210.0341, 210.0683, 210.1248, 210.164, 
    210.1673, 210.1432, 210.0956, 210.0362, 209.9704, 209.9066, 209.8657, 
    209.8374,
  210.22, 210.1763, 210.1408, 210.1031, 210.1199, 210.1656, 210.2031, 
    210.2257, 210.2227, 210.1817, 210.1173, 210.037, 209.9563, 209.8982, 
    209.8724,
  210.3337, 210.2798, 210.2588, 210.2055, 210.2025, 210.2369, 210.2653, 
    210.298, 210.304, 210.2798, 210.2352, 210.1545, 210.0473, 209.9621, 
    209.9083,
  210.4475, 210.3976, 210.3719, 210.3212, 210.2994, 210.3043, 210.3337, 
    210.3657, 210.3795, 210.3651, 210.3346, 210.2718, 210.1673, 210.0382, 
    209.947,
  210.5783, 210.5387, 210.4922, 210.4226, 210.391, 210.3791, 210.406, 
    210.4561, 210.4884, 210.4959, 210.4736, 210.4117, 210.3204, 210.18, 
    210.0314,
  210.6618, 210.6143, 210.5731, 210.5238, 210.4895, 210.4688, 210.4672, 
    210.5112, 210.5692, 210.5944, 210.5954, 210.567, 210.483, 210.3653, 
    210.2067,
  210.6982, 210.6888, 210.6705, 210.6261, 210.557, 210.5286, 210.5397, 
    210.5388, 210.611, 210.6678, 210.6873, 210.692, 210.6379, 210.5474, 
    210.4084,
  210.7156, 210.7333, 210.7261, 210.67, 210.639, 210.6195, 210.5866, 
    210.5833, 210.6077, 210.6761, 210.7333, 210.7635, 210.7605, 210.7067, 
    210.6138,
  210.7542, 210.7547, 210.755, 210.7674, 210.7542, 210.6773, 210.6525, 
    210.6303, 210.6352, 210.662, 210.7196, 210.7904, 210.8229, 210.8275, 
    210.7832,
  210.0197, 209.8503, 209.7449, 209.6828, 209.6677, 209.6679, 209.6747, 
    209.6722, 209.6352, 209.561, 209.4355, 209.2946, 209.1457, 208.9815, 
    208.8242,
  210.1838, 210.0223, 209.8708, 209.7673, 209.7057, 209.692, 209.705, 
    209.708, 209.7127, 209.6871, 209.6136, 209.5076, 209.3726, 209.2294, 
    209.059,
  210.3553, 210.217, 210.0503, 209.9065, 209.7937, 209.7374, 209.7198, 
    209.7253, 209.7428, 209.7497, 209.7222, 209.653, 209.5502, 209.4152, 
    209.2711,
  210.5157, 210.424, 210.2843, 210.1236, 209.9869, 209.8674, 209.7965, 
    209.7646, 209.769, 209.7832, 209.7816, 209.7494, 209.6856, 209.5931, 
    209.4767,
  210.6036, 210.5626, 210.48, 210.3481, 210.195, 210.0541, 209.948, 209.8726, 
    209.839, 209.8103, 209.813, 209.8026, 209.7717, 209.7055, 209.627,
  210.6509, 210.6499, 210.6315, 210.5294, 210.4047, 210.2558, 210.1296, 
    210.0276, 209.9791, 209.9388, 209.9095, 209.886, 209.8641, 209.8118, 
    209.7384,
  210.6828, 210.669, 210.6658, 210.6403, 210.5801, 210.4438, 210.2922, 
    210.1726, 210.1047, 210.0631, 210.0279, 209.9936, 209.9689, 209.9362, 
    209.879,
  210.7099, 210.7029, 210.7134, 210.6934, 210.6526, 210.5736, 210.4605, 
    210.3179, 210.2271, 210.1674, 210.1242, 210.0876, 210.0617, 210.0384, 
    210.0092,
  210.7259, 210.7321, 210.7381, 210.7054, 210.7117, 210.6985, 210.5821, 
    210.4652, 210.3429, 210.2805, 210.2254, 210.1897, 210.1522, 210.1368, 
    210.1254,
  210.7729, 210.752, 210.762, 210.7915, 210.8205, 210.7732, 210.703, 
    210.5955, 210.4707, 210.3408, 210.2919, 210.2408, 210.2074, 210.1818, 
    210.1912,
  208.6077, 208.5495, 208.4977, 208.4505, 208.4003, 208.3518, 208.3318, 
    208.3203, 208.3304, 208.3376, 208.3563, 208.3622, 208.3623, 208.3476, 
    208.317,
  208.7764, 208.6865, 208.6421, 208.5781, 208.5444, 208.4926, 208.4635, 
    208.4521, 208.456, 208.4658, 208.4898, 208.5088, 208.5259, 208.5294, 
    208.5169,
  208.8743, 208.7893, 208.7594, 208.7012, 208.6762, 208.6061, 208.5668, 
    208.5401, 208.5427, 208.5473, 208.5744, 208.6072, 208.6445, 208.6759, 
    208.6886,
  209.0233, 208.95, 208.9103, 208.8194, 208.7872, 208.7142, 208.6727, 
    208.649, 208.6427, 208.653, 208.6753, 208.7028, 208.7441, 208.7833, 
    208.8137,
  209.1591, 209.1082, 209.0614, 208.9776, 208.9374, 208.8588, 208.813, 
    208.7744, 208.7477, 208.7538, 208.768, 208.7855, 208.8167, 208.8645, 
    208.9107,
  209.2664, 209.2245, 209.1844, 209.1161, 209.0524, 208.9771, 208.9223, 
    208.8625, 208.8438, 208.8423, 208.8627, 208.8811, 208.9025, 208.9341, 
    208.9813,
  209.3989, 209.3217, 209.2796, 209.2473, 209.213, 209.1302, 209.0593, 
    208.9928, 208.9587, 208.9366, 208.9507, 208.9625, 208.9894, 209.0136, 
    209.0512,
  209.5227, 209.4355, 209.4081, 209.368, 209.3452, 209.2676, 209.2079, 
    209.1182, 209.0701, 209.0298, 209.0182, 209.0284, 209.0612, 209.0946, 
    209.1315,
  209.6431, 209.5747, 209.5268, 209.4467, 209.4621, 209.4333, 209.3455, 
    209.2699, 209.2023, 209.1363, 209.1011, 209.0891, 209.1262, 209.1647, 
    209.2126,
  209.7859, 209.6829, 209.6222, 209.6034, 209.6414, 209.5585, 209.4878, 
    209.4124, 209.3294, 209.2422, 209.1825, 209.1495, 209.1673, 209.2023, 
    209.2561,
  208.9999, 208.9482, 208.9081, 208.8743, 208.8386, 208.795, 208.7456, 
    208.6743, 208.5983, 208.5024, 208.417, 208.3257, 208.2454, 208.1681, 
    208.0924,
  209.1369, 209.0633, 209.0275, 208.9947, 208.9875, 208.959, 208.9183, 
    208.8492, 208.7821, 208.6915, 208.6136, 208.5235, 208.4364, 208.3473, 
    208.2604,
  209.1941, 209.1256, 209.115, 209.1022, 209.1011, 209.0796, 209.0534, 
    209.0095, 208.9629, 208.8892, 208.8236, 208.7429, 208.6585, 208.557, 
    208.4547,
  209.2455, 209.2144, 209.2072, 209.1909, 209.1987, 209.1926, 209.1909, 
    209.1658, 209.1263, 209.0676, 209.0087, 208.94, 208.8669, 208.7612, 
    208.6565,
  209.2668, 209.2583, 209.2537, 209.2551, 209.2788, 209.2711, 209.2789, 
    209.2614, 209.2299, 209.1932, 209.1509, 209.1012, 209.044, 208.9691, 
    208.8863,
  209.2518, 209.2677, 209.2719, 209.2812, 209.3011, 209.3091, 209.3356, 
    209.3257, 209.3013, 209.2675, 209.2298, 209.1886, 209.1493, 209.1079, 
    209.0589,
  209.2215, 209.2398, 209.2458, 209.2718, 209.3256, 209.3487, 209.382, 
    209.3756, 209.3502, 209.3079, 209.2544, 209.214, 209.1814, 209.1563, 
    209.128,
  209.1827, 209.1997, 209.2331, 209.2622, 209.3205, 209.3749, 209.4305, 
    209.425, 209.3982, 209.3564, 209.2962, 209.2497, 209.2092, 209.179, 
    209.1492,
  209.1685, 209.1907, 209.2289, 209.2213, 209.2978, 209.3799, 209.4285, 
    209.4592, 209.4509, 209.4096, 209.3643, 209.3105, 209.2581, 209.2085, 
    209.185,
  209.1916, 209.1851, 209.2045, 209.2487, 209.331, 209.3557, 209.4164, 
    209.4616, 209.4732, 209.4452, 209.4117, 209.3764, 209.3078, 209.2561, 
    209.2231,
  210.6251, 210.6004, 210.5711, 210.5354, 210.5187, 210.5367, 210.581, 
    210.6229, 210.6665, 210.6976, 210.707, 210.6982, 210.6935, 210.6662, 
    210.6253,
  210.6934, 210.7038, 210.6623, 210.6218, 210.6091, 210.6084, 210.6362, 
    210.66, 210.7013, 210.7476, 210.7872, 210.8115, 210.8303, 210.8185, 
    210.7939,
  210.7078, 210.7371, 210.7378, 210.7328, 210.7019, 210.6685, 210.6812, 
    210.7027, 210.7582, 210.8163, 210.8611, 210.8879, 210.9072, 210.8991, 
    210.8966,
  210.7101, 210.7756, 210.8194, 210.8225, 210.8097, 210.7633, 210.7684, 
    210.7795, 210.8163, 210.8645, 210.9214, 210.968, 211.0002, 211.011, 
    211.0214,
  210.721, 210.7825, 210.8528, 210.8792, 210.9083, 210.8694, 210.8573, 
    210.8427, 210.8618, 210.8939, 210.9657, 211.0168, 211.0481, 211.0791, 
    211.1055,
  210.735, 210.7699, 210.8578, 210.9158, 210.964, 210.9652, 210.9623, 
    210.9376, 210.9466, 210.9619, 211.0115, 211.0501, 211.0682, 211.1125, 
    211.1615,
  210.7452, 210.7538, 210.8173, 210.8967, 210.9823, 211.0212, 211.029, 
    211.0189, 211.0434, 211.0497, 211.0697, 211.1021, 211.1188, 211.1748, 
    211.2125,
  210.7678, 210.7527, 210.7988, 210.8724, 210.9632, 211.0425, 211.0912, 
    211.1012, 211.1505, 211.1678, 211.1668, 211.1748, 211.1923, 211.2445, 
    211.2822,
  210.7971, 210.7934, 210.829, 210.8433, 210.9268, 211.037, 211.1061, 
    211.1651, 211.2419, 211.271, 211.2762, 211.2775, 211.2809, 211.3316, 
    211.3511,
  210.8897, 210.8601, 210.8654, 210.8973, 210.9664, 211.0226, 211.092, 
    211.1827, 211.3014, 211.3552, 211.3886, 211.4037, 211.3962, 211.4204, 
    211.4352,
  211.717, 211.6832, 211.5692, 211.4775, 211.3969, 211.3368, 211.2283, 
    211.1192, 210.9873, 210.8279, 210.7039, 210.5905, 210.5029, 210.4068, 
    210.3473,
  211.7803, 211.7183, 211.59, 211.5008, 211.4226, 211.3575, 211.2836, 
    211.2112, 211.0839, 210.9433, 210.8005, 210.6746, 210.5933, 210.4935, 
    210.4258,
  211.7668, 211.6885, 211.5751, 211.484, 211.3895, 211.3335, 211.2855, 
    211.2346, 211.1427, 211.0288, 210.9036, 210.7786, 210.7034, 210.5871, 
    210.4945,
  211.7623, 211.7063, 211.6036, 211.505, 211.4072, 211.3369, 211.2945, 
    211.2615, 211.1922, 211.0988, 210.9859, 210.8776, 210.7859, 210.6902, 
    210.6073,
  211.7948, 211.729, 211.6122, 211.5202, 211.4338, 211.3469, 211.3027, 
    211.2816, 211.2476, 211.1785, 211.0787, 210.9808, 210.8774, 210.7855, 
    210.7017,
  211.8228, 211.7531, 211.652, 211.5494, 211.4409, 211.3646, 211.3297, 
    211.3048, 211.3044, 211.2578, 211.1708, 211.0851, 210.984, 210.895, 
    210.7971,
  211.8741, 211.7932, 211.6773, 211.5567, 211.4835, 211.4011, 211.3618, 
    211.3338, 211.355, 211.3351, 211.2835, 211.2114, 211.1173, 211.0241, 
    210.9063,
  211.9466, 211.8398, 211.7257, 211.6116, 211.533, 211.4675, 211.4286, 
    211.3824, 211.387, 211.3924, 211.366, 211.316, 211.2344, 211.1617, 
    211.0438,
  212.0069, 211.9202, 211.8139, 211.6726, 211.5776, 211.5415, 211.5043, 
    211.4528, 211.4278, 211.4277, 211.4266, 211.3916, 211.3285, 211.249, 
    211.1615,
  212.0527, 211.9841, 211.8843, 211.7806, 211.7136, 211.6454, 211.5719, 
    211.5186, 211.4937, 211.4753, 211.4674, 211.4342, 211.3864, 211.314, 
    211.2537,
  209.2146, 209.1168, 209.0117, 208.9331, 208.831, 208.7444, 208.6145, 
    208.5054, 208.3862, 208.2732, 208.1709, 208.0495, 207.959, 207.8303, 
    207.6786,
  209.2946, 209.2218, 209.1313, 209.0349, 208.9269, 208.8396, 208.7191, 
    208.6039, 208.464, 208.3459, 208.2307, 208.1342, 208.0555, 207.9426, 
    207.8227,
  209.3649, 209.3144, 209.2546, 209.1451, 209.0356, 208.936, 208.8076, 
    208.6949, 208.5695, 208.4428, 208.3121, 208.1966, 208.099, 207.9976, 
    207.9074,
  209.4738, 209.4021, 209.3422, 209.241, 209.1421, 209.0284, 208.9106, 
    208.8049, 208.6719, 208.5351, 208.4022, 208.2725, 208.1622, 208.0603, 
    207.9745,
  209.5757, 209.4966, 209.4329, 209.3565, 209.2673, 209.1545, 209.0437, 
    208.9172, 208.7791, 208.6324, 208.501, 208.3669, 208.2449, 208.1397, 
    208.055,
  209.6753, 209.6021, 209.5566, 209.4655, 209.3502, 209.2611, 209.1559, 
    209.029, 208.9051, 208.7725, 208.6342, 208.4948, 208.3633, 208.2429, 
    208.1445,
  209.7758, 209.7016, 209.6417, 209.546, 209.46, 209.3571, 209.2468, 
    209.1415, 209.0207, 208.8992, 208.7637, 208.6292, 208.5078, 208.3737, 
    208.2633,
  209.8932, 209.7917, 209.732, 209.6558, 209.5701, 209.4431, 209.3464, 
    209.2304, 209.1263, 209.0222, 208.8974, 208.7722, 208.6451, 208.5203, 
    208.4002,
  209.9948, 209.9062, 209.847, 209.7261, 209.6325, 209.5538, 209.4544, 
    209.3233, 209.2139, 209.1039, 208.9995, 208.8876, 208.7744, 208.657, 
    208.5469,
  210.1277, 210.0314, 209.9432, 209.8476, 209.7883, 209.6804, 209.5454, 
    209.4252, 209.3067, 209.1807, 209.084, 208.9784, 208.8813, 208.7746, 
    208.6685,
  207.3066, 207.2828, 207.2595, 207.2278, 207.1738, 207.0962, 207.0243, 
    206.9523, 206.8692, 206.7773, 206.7023, 206.6421, 206.6019, 206.5583, 
    206.5227,
  207.3594, 207.3305, 207.3068, 207.295, 207.2748, 207.2333, 207.1829, 
    207.102, 207.0235, 206.937, 206.8788, 206.8295, 206.7912, 206.7421, 
    206.6888,
  207.4546, 207.379, 207.3721, 207.3573, 207.3399, 207.3291, 207.295, 
    207.2181, 207.1496, 207.0744, 207.035, 206.9899, 206.9564, 206.9025, 
    206.8473,
  207.5494, 207.4707, 207.4614, 207.416, 207.3852, 207.3759, 207.3575, 
    207.3169, 207.2577, 207.2009, 207.1612, 207.1297, 207.0949, 207.0455, 
    206.9931,
  207.6257, 207.5638, 207.5389, 207.4964, 207.4561, 207.4271, 207.4152, 
    207.3991, 207.3536, 207.3172, 207.2765, 207.2498, 207.2025, 207.1567, 
    207.1034,
  207.6864, 207.628, 207.6042, 207.5631, 207.4995, 207.4648, 207.464, 
    207.4706, 207.4474, 207.421, 207.3764, 207.3351, 207.2889, 207.235, 
    207.1998,
  207.76, 207.683, 207.6232, 207.5869, 207.5508, 207.4959, 207.4832, 
    207.4975, 207.5035, 207.5004, 207.468, 207.4253, 207.3775, 207.3288, 
    207.2933,
  207.8533, 207.7416, 207.6668, 207.6235, 207.592, 207.5309, 207.5198, 
    207.5154, 207.5331, 207.5473, 207.535, 207.4999, 207.4586, 207.4166, 
    207.3802,
  207.9328, 207.8457, 207.7697, 207.6646, 207.6102, 207.5879, 207.5618, 
    207.5398, 207.5419, 207.5602, 207.5756, 207.5683, 207.5431, 207.5037, 
    207.471,
  208.0367, 207.9352, 207.8624, 207.7715, 207.7248, 207.6644, 207.5967, 
    207.5824, 207.5757, 207.58, 207.5925, 207.6077, 207.6004, 207.58, 207.5448,
  208.3607, 208.3844, 208.3752, 208.3831, 208.3724, 208.4083, 208.4629, 
    208.5036, 208.5263, 208.5399, 208.5634, 208.5775, 208.6053, 208.6213, 
    208.6449,
  208.487, 208.5003, 208.4919, 208.5188, 208.5261, 208.5668, 208.6191, 
    208.6463, 208.6659, 208.6864, 208.7198, 208.7532, 208.8004, 208.8442, 
    208.8809,
  208.6416, 208.6184, 208.619, 208.6454, 208.6429, 208.6818, 208.7181, 
    208.7459, 208.7904, 208.841, 208.8937, 208.9425, 209.0072, 209.0648, 
    209.1019,
  208.7876, 208.77, 208.7572, 208.7482, 208.7383, 208.7501, 208.789, 
    208.8339, 208.8783, 208.9242, 208.9819, 209.04, 209.1018, 209.1573, 
    209.1929,
  208.9318, 208.9227, 208.8985, 208.9091, 208.8864, 208.871, 208.8915, 
    208.9298, 208.9824, 209.0284, 209.0904, 209.1552, 209.2245, 209.2867, 
    209.3453,
  209.0529, 209.0535, 209.0707, 209.0897, 209.0472, 209.0175, 208.9975, 
    209.031, 209.0813, 209.1321, 209.1864, 209.2424, 209.3136, 209.3949, 
    209.4812,
  209.1822, 209.1671, 209.1942, 209.2129, 209.2176, 209.1751, 209.1157, 
    209.1296, 209.1693, 209.224, 209.2867, 209.3463, 209.4322, 209.5208, 
    209.6305,
  209.3282, 209.2933, 209.3295, 209.3448, 209.359, 209.338, 209.2829, 209.25, 
    209.2494, 209.3129, 209.3752, 209.4396, 209.5134, 209.6113, 209.7318,
  209.4794, 209.443, 209.4825, 209.4464, 209.4509, 209.4977, 209.4404, 
    209.4062, 209.3707, 209.3896, 209.434, 209.4942, 209.5777, 209.6758, 
    209.8107,
  209.651, 209.5845, 209.5948, 209.5861, 209.6329, 209.6388, 209.5674, 
    209.5453, 209.4956, 209.4819, 209.4906, 209.5446, 209.6224, 209.7233, 
    209.8503,
  210.0802, 210.0431, 210.0598, 210.0838, 210.0956, 210.1198, 210.1412, 
    210.1387, 210.1188, 210.1076, 210.1096, 210.1049, 210.0873, 210.089, 
    210.054,
  210.2092, 210.1776, 210.1805, 210.2088, 210.2278, 210.2486, 210.27, 
    210.2814, 210.2781, 210.2783, 210.2732, 210.2451, 210.223, 210.2235, 
    210.2094,
  210.3516, 210.3057, 210.3051, 210.3033, 210.278, 210.2813, 210.323, 
    210.3798, 210.4131, 210.4568, 210.4747, 210.4634, 210.4736, 210.4839, 
    210.5177,
  210.5274, 210.4435, 210.4174, 210.4079, 210.3913, 210.3943, 210.411, 
    210.4846, 210.5383, 210.5937, 210.6112, 210.6131, 210.6208, 210.6014, 
    210.6535,
  210.7314, 210.594, 210.5452, 210.5402, 210.5331, 210.5051, 210.4734, 
    210.5403, 210.6054, 210.6824, 210.7271, 210.7717, 210.7679, 210.7211, 
    210.7564,
  210.9457, 210.8189, 210.7665, 210.7137, 210.6579, 210.6126, 210.5654, 
    210.6026, 210.6607, 210.7181, 210.7715, 210.8484, 210.8789, 210.8811, 
    210.8938,
  211.1735, 211.0448, 210.9326, 210.8327, 210.8412, 210.7721, 210.6956, 
    210.6814, 210.7, 210.7395, 210.7916, 210.864, 210.9403, 211.0193, 211.0679,
  211.3593, 211.2367, 211.092, 210.975, 210.9629, 210.8942, 210.8136, 
    210.741, 210.7254, 210.7637, 210.8219, 210.8762, 210.9632, 211.0746, 
    211.1512,
  211.4929, 211.3955, 211.2676, 211.1164, 211.0266, 211.0213, 210.9487, 
    210.8637, 210.7953, 210.7862, 210.8351, 210.8669, 210.922, 211.0164, 
    211.1101,
  211.5756, 211.4831, 211.3543, 211.2273, 211.1693, 211.1447, 211.035, 
    210.9204, 210.8599, 210.8066, 210.8116, 210.8528, 210.8895, 210.9743, 
    211.0689,
  209.4055, 209.3383, 209.302, 209.2791, 209.2622, 209.2225, 209.1814, 
    209.1238, 209.0675, 208.9993, 208.9293, 208.858, 208.7948, 208.7349, 
    208.7081,
  209.5166, 209.406, 209.3412, 209.2976, 209.2798, 209.2531, 209.2272, 
    209.1704, 209.1104, 209.0361, 208.979, 208.9139, 208.8194, 208.751, 
    208.6902,
  209.6384, 209.5112, 209.4165, 209.3583, 209.3148, 209.2863, 209.2628, 
    209.2278, 209.1781, 209.1082, 209.0435, 208.9744, 208.9001, 208.8433, 
    208.7511,
  209.7626, 209.6501, 209.5368, 209.4359, 209.3536, 209.3048, 209.2773, 
    209.2556, 209.2229, 209.1736, 209.1043, 209.0258, 208.9689, 208.8954, 
    208.8136,
  209.8397, 209.7348, 209.642, 209.5365, 209.4182, 209.3247, 209.2627, 
    209.237, 209.2237, 209.1932, 209.1321, 209.0629, 209.0082, 208.9455, 
    208.8866,
  209.8881, 209.799, 209.7347, 209.6429, 209.5173, 209.4061, 209.3235, 
    209.2644, 209.2556, 209.2205, 209.1878, 209.1116, 209.0441, 208.9658, 
    208.904,
  209.9003, 209.792, 209.6981, 209.6446, 209.588, 209.4742, 209.3694, 
    209.2901, 209.247, 209.2348, 209.2047, 209.1475, 209.0705, 208.9785, 
    208.9102,
  209.8526, 209.7219, 209.6264, 209.5754, 209.5414, 209.4774, 209.4118, 
    209.3144, 209.2509, 209.2254, 209.1912, 209.1433, 209.0844, 209.0238, 
    208.9805,
  209.7901, 209.6549, 209.5527, 209.452, 209.4365, 209.4241, 209.3777, 
    209.3246, 209.2855, 209.2502, 209.2147, 209.1618, 209.091, 209.0414, 
    209.0027,
  209.761, 209.6182, 209.4913, 209.4108, 209.383, 209.3142, 209.2858, 
    209.241, 209.2359, 209.2188, 209.2074, 209.1647, 209.1107, 209.065, 
    209.0292,
  207.976, 207.9076, 207.9012, 207.8976, 207.9096, 207.921, 207.9501, 
    207.9743, 208.0243, 208.0779, 208.1396, 208.1782, 208.2038, 208.2157, 
    208.2045,
  208.0352, 207.9656, 207.926, 207.9057, 207.9004, 207.9033, 207.9212, 
    207.9528, 208.0079, 208.0648, 208.1262, 208.178, 208.2254, 208.2579, 
    208.2877,
  208.1335, 208.0269, 207.9753, 207.9428, 207.9148, 207.908, 207.9135, 
    207.929, 207.9688, 208.0167, 208.0872, 208.1589, 208.2288, 208.3, 208.351,
  208.2688, 208.1261, 208.0437, 207.9852, 207.9453, 207.931, 207.9314, 
    207.9412, 207.9618, 207.9976, 208.0498, 208.1214, 208.2135, 208.3087, 
    208.3907,
  208.4613, 208.2732, 208.1484, 208.0646, 208.0083, 207.972, 207.9555, 
    207.9689, 207.9716, 207.9852, 208.0182, 208.0971, 208.1966, 208.3154, 
    208.4161,
  208.6456, 208.4628, 208.3293, 208.2105, 208.0851, 208.042, 208.0151, 
    208.0183, 208.01, 208.0149, 208.0282, 208.0725, 208.1635, 208.294, 
    208.4172,
  208.7886, 208.6585, 208.5005, 208.361, 208.2286, 208.148, 208.087, 
    208.0771, 208.0766, 208.0793, 208.0755, 208.0941, 208.1555, 208.264, 
    208.4008,
  208.8922, 208.7986, 208.6694, 208.549, 208.4079, 208.2862, 208.2161, 
    208.1545, 208.1519, 208.1653, 208.1602, 208.1544, 208.1777, 208.2557, 
    208.3672,
  208.9536, 208.8949, 208.8177, 208.7021, 208.5454, 208.4725, 208.3678, 
    208.2734, 208.2443, 208.2405, 208.2504, 208.2406, 208.2429, 208.2713, 
    208.3507,
  208.9968, 208.9471, 208.9207, 208.8841, 208.7853, 208.6743, 208.5307, 
    208.4122, 208.366, 208.3267, 208.3343, 208.3354, 208.3251, 208.33, 
    208.3723,
  208.5824, 208.6521, 208.6886, 208.7589, 208.79, 208.8427, 208.8927, 
    208.9335, 208.9435, 208.9238, 208.8824, 208.8196, 208.7521, 208.6772, 
    208.6201,
  208.5585, 208.6685, 208.6911, 208.766, 208.807, 208.8647, 208.9142, 
    208.9614, 208.9973, 209.0062, 208.9954, 208.9501, 208.888, 208.8071, 
    208.7439,
  208.5078, 208.6324, 208.691, 208.7802, 208.8234, 208.8792, 208.9315, 
    208.9706, 209.024, 209.0565, 209.0869, 209.0776, 209.0442, 208.962, 
    208.8776,
  208.4531, 208.5832, 208.6829, 208.7766, 208.8338, 208.8931, 208.9536, 
    209.0001, 209.0591, 209.0961, 209.136, 209.1533, 209.1515, 209.1082, 
    209.0436,
  208.4623, 208.5434, 208.6582, 208.7463, 208.8428, 208.9079, 208.972, 
    209.0324, 209.0986, 209.1333, 209.1734, 209.1991, 209.2188, 209.2217, 
    209.1992,
  208.5222, 208.5536, 208.6602, 208.7325, 208.8147, 208.9023, 208.9913, 
    209.0713, 209.1287, 209.176, 209.2148, 209.2426, 209.2638, 209.2843, 
    209.2755,
  208.6268, 208.6208, 208.6809, 208.7263, 208.8208, 208.9081, 208.9864, 
    209.0848, 209.169, 209.2317, 209.2733, 209.2941, 209.307, 209.3136, 
    209.3111,
  208.7802, 208.7431, 208.7511, 208.7791, 208.8605, 208.9164, 208.9976, 
    209.0809, 209.1788, 209.2707, 209.3399, 209.3614, 209.3608, 209.3485, 
    209.326,
  208.9594, 208.9044, 208.8914, 208.8736, 208.9046, 208.9641, 209.0219, 
    209.0849, 209.191, 209.2822, 209.3733, 209.4124, 209.4255, 209.4072, 
    209.3918,
  209.2402, 209.1401, 209.0813, 209.0437, 209.0546, 209.0792, 209.0764, 
    209.1141, 209.2059, 209.2851, 209.3774, 209.4357, 209.4727, 209.4751, 
    209.4611,
  208.3091, 208.3206, 208.2745, 208.2303, 208.1645, 208.1081, 208.0532, 
    207.9823, 207.8889, 207.781, 207.6801, 207.5891, 207.5348, 207.4971, 
    207.4369,
  208.2474, 208.275, 208.2469, 208.246, 208.2153, 208.1835, 208.1461, 
    208.081, 207.9957, 207.882, 207.7716, 207.6743, 207.6088, 207.5427, 
    207.4635,
  208.1644, 208.1986, 208.1899, 208.2202, 208.2128, 208.2132, 208.1874, 
    208.1423, 208.0719, 207.9659, 207.8509, 207.7496, 207.6783, 207.604, 
    207.5425,
  208.0672, 208.1228, 208.1372, 208.1718, 208.1886, 208.201, 208.1821, 
    208.1443, 208.09, 208.0059, 207.9124, 207.8158, 207.7275, 207.6485, 
    207.5845,
  208.0251, 208.0419, 208.078, 208.1433, 208.1643, 208.1762, 208.1579, 
    208.1271, 208.0871, 208.036, 207.9721, 207.908, 207.8475, 207.7805, 
    207.6928,
  207.9971, 208.0012, 208.0811, 208.1407, 208.1244, 208.1399, 208.1327, 
    208.1043, 208.081, 208.0784, 208.0531, 208.0283, 207.9935, 207.9404, 
    207.8371,
  208.0202, 208.025, 208.0622, 208.0904, 208.14, 208.1399, 208.1397, 
    208.1331, 208.105, 208.1039, 208.0899, 208.0668, 208.033, 207.9816, 
    207.8994,
  208.0653, 208.061, 208.0507, 208.0714, 208.1399, 208.1266, 208.1387, 
    208.1299, 208.1203, 208.1165, 208.0974, 208.0794, 208.0361, 207.9846, 
    207.9444,
  208.104, 208.1146, 208.1246, 208.1002, 208.071, 208.1024, 208.1366, 
    208.1197, 208.1193, 208.1076, 208.0901, 208.0774, 208.0448, 207.9953, 
    207.9549,
  208.232, 208.2113, 208.1865, 208.1656, 208.1475, 208.1609, 208.1216, 
    208.0439, 208.0979, 208.1162, 208.1356, 208.1241, 208.0778, 208.0029, 
    207.9434,
  207.4881, 207.3671, 207.2387, 207.0941, 206.9635, 206.8285, 206.7128, 
    206.6155, 206.5414, 206.4697, 206.388, 206.3132, 206.2431, 206.1855, 
    206.1372,
  207.608, 207.5122, 207.3702, 207.2232, 207.1026, 206.9661, 206.8449, 
    206.7303, 206.6373, 206.5393, 206.4452, 206.3668, 206.3025, 206.2375, 
    206.1796,
  207.685, 207.5977, 207.4869, 207.3839, 207.2651, 207.1411, 207.0205, 
    206.8906, 206.757, 206.6328, 206.5218, 206.4289, 206.3543, 206.2841, 
    206.2192,
  207.7438, 207.6566, 207.5848, 207.4893, 207.3912, 207.2898, 207.1835, 
    207.0534, 206.924, 206.7801, 206.6352, 206.5115, 206.4165, 206.3391, 
    206.2711,
  207.8234, 207.7316, 207.6459, 207.5414, 207.4501, 207.365, 207.2769, 
    207.1749, 207.0555, 206.9316, 206.7821, 206.627, 206.4864, 206.389, 
    206.3224,
  207.9002, 207.7984, 207.7141, 207.6098, 207.4816, 207.3797, 207.3019, 
    207.2167, 207.1349, 207.0435, 206.9207, 206.7646, 206.6067, 206.478, 
    206.3963,
  207.9695, 207.8606, 207.76, 207.6155, 207.4792, 207.3703, 207.2949, 
    207.2242, 207.149, 207.083, 207.0039, 206.8932, 206.748, 206.6073, 206.493,
  208.0006, 207.8755, 207.7729, 207.6496, 207.5402, 207.4316, 207.3452, 
    207.2613, 207.1942, 207.1236, 207.0487, 206.9784, 206.8803, 206.7631, 
    206.6457,
  207.9809, 207.8603, 207.7811, 207.6577, 207.5648, 207.5173, 207.4621, 
    207.39, 207.3195, 207.2419, 207.1473, 207.0639, 206.9736, 206.8833, 
    206.7911,
  207.981, 207.8564, 207.7666, 207.7089, 207.7006, 207.6931, 207.6277, 
    207.5308, 207.4753, 207.3608, 207.2457, 207.1534, 207.0723, 206.9927, 
    206.9253,
  206.1692, 206.1219, 206.122, 206.1454, 206.1783, 206.2177, 206.2589, 
    206.2851, 206.3123, 206.3432, 206.3668, 206.3814, 206.3883, 206.3805, 
    206.3722,
  206.33, 206.2909, 206.2511, 206.2445, 206.2596, 206.2836, 206.3118, 
    206.3301, 206.3591, 206.3927, 206.4313, 206.4631, 206.4912, 206.5068, 
    206.521,
  206.5225, 206.4602, 206.4095, 206.3768, 206.3642, 206.3638, 206.3632, 
    206.3614, 206.3799, 206.4133, 206.4615, 206.5175, 206.5679, 206.6038, 
    206.6359,
  206.6947, 206.6181, 206.5724, 206.5239, 206.4847, 206.4582, 206.4374, 
    206.4132, 206.4106, 206.4303, 206.4756, 206.5308, 206.5978, 206.6668, 
    206.7104,
  206.8845, 206.7931, 206.7264, 206.6575, 206.6143, 206.5788, 206.5421, 
    206.5062, 206.4781, 206.4792, 206.492, 206.5432, 206.6053, 206.6802, 
    206.7422,
  207.035, 206.9489, 206.8811, 206.8138, 206.7588, 206.7376, 206.7149, 
    206.6804, 206.6367, 206.5982, 206.5914, 206.6078, 206.6459, 206.7092, 
    206.7804,
  207.1804, 207.1009, 207.0247, 206.9627, 206.9384, 206.9394, 206.9409, 
    206.9084, 206.8593, 206.7888, 206.7398, 206.7286, 206.7328, 206.786, 
    206.8441,
  207.2836, 207.2206, 207.1646, 207.1267, 207.1435, 207.1685, 207.1748, 
    207.1346, 207.0533, 206.955, 206.8708, 206.8305, 206.8296, 206.8544, 
    206.9287,
  207.3859, 207.3395, 207.3279, 207.3193, 207.3316, 207.353, 207.3333, 
    207.2649, 207.1738, 207.0801, 206.9877, 206.9301, 206.9049, 206.9175, 
    206.9794,
  207.5068, 207.452, 207.4502, 207.475, 207.4958, 207.469, 207.3807, 
    207.3033, 207.2525, 207.2195, 207.1743, 207.1197, 207.0664, 207.0556, 
    207.067,
  207.9992, 208.0871, 208.1488, 208.2024, 208.2358, 208.2728, 208.2955, 
    208.3192, 208.3498, 208.3925, 208.4492, 208.4998, 208.5437, 208.5751, 
    208.605,
  207.9881, 208.0937, 208.1677, 208.2321, 208.2911, 208.3442, 208.384, 
    208.4199, 208.452, 208.5008, 208.558, 208.6075, 208.6493, 208.6864, 
    208.7233,
  208.0239, 208.1183, 208.1951, 208.2805, 208.3584, 208.416, 208.4596, 
    208.4949, 208.535, 208.6, 208.6594, 208.7115, 208.7579, 208.8029, 208.8588,
  208.0768, 208.1587, 208.2407, 208.3208, 208.3863, 208.4568, 208.5238, 
    208.5812, 208.6496, 208.7252, 208.7679, 208.8057, 208.8464, 208.8919, 
    208.9508,
  208.1877, 208.243, 208.2936, 208.3488, 208.4137, 208.4937, 208.5757, 
    208.6664, 208.7473, 208.8125, 208.8429, 208.8695, 208.8956, 208.9376, 
    209.0085,
  208.305, 208.3418, 208.3769, 208.4174, 208.4609, 208.538, 208.6416, 
    208.7411, 208.8149, 208.8635, 208.8786, 208.9112, 208.9639, 209.0394, 
    209.1133,
  208.4445, 208.4691, 208.4768, 208.487, 208.5421, 208.625, 208.7148, 
    208.7981, 208.8467, 208.8678, 208.9075, 208.9865, 209.0587, 209.112, 
    209.1649,
  208.5571, 208.5771, 208.5888, 208.5986, 208.6612, 208.7331, 208.8069, 
    208.851, 208.8539, 208.8618, 208.8802, 208.9794, 209.054, 209.1151, 
    209.1944,
  208.6609, 208.6753, 208.7099, 208.7131, 208.7695, 208.8511, 208.8932, 
    208.8936, 208.8714, 208.851, 208.9151, 209.0368, 209.0856, 209.1366, 
    209.2383,
  208.7538, 208.7639, 208.7901, 208.8363, 208.9166, 208.9672, 208.9631, 
    208.9378, 208.9276, 208.938, 209.0032, 209.0878, 209.1016, 209.1705, 
    209.2959,
  209.6112, 209.6082, 209.5835, 209.5699, 209.5736, 209.5919, 209.6071, 
    209.6261, 209.612, 209.6039, 209.6243, 209.6384, 209.6391, 209.591, 
    209.4806,
  209.6773, 209.6844, 209.6641, 209.6412, 209.6402, 209.6476, 209.6607, 
    209.6716, 209.6764, 209.7172, 209.7692, 209.8045, 209.7897, 209.6878, 
    209.5706,
  209.7486, 209.7619, 209.7448, 209.7351, 209.7416, 209.7487, 209.7586, 
    209.7605, 209.7718, 209.8328, 209.8956, 209.9467, 209.9154, 209.8024, 
    209.7171,
  209.7938, 209.8171, 209.8215, 209.8146, 209.8208, 209.8299, 209.8441, 
    209.8505, 209.8647, 209.9291, 209.9859, 210.0315, 209.9682, 209.8701, 
    209.8022,
  209.8467, 209.8843, 209.8934, 209.8889, 209.9009, 209.9138, 209.9326, 
    209.9337, 209.9419, 209.9999, 210.0758, 210.1254, 210.0746, 209.9982, 
    209.9247,
  209.8899, 209.9268, 209.9458, 209.9486, 209.9547, 209.9646, 209.9894, 
    209.9825, 209.9987, 210.0881, 210.1768, 210.2189, 210.1887, 210.1175, 
    210.0272,
  209.9321, 209.9478, 209.9656, 209.9603, 209.9858, 210.0029, 210.0181, 
    210.0121, 210.052, 210.1483, 210.2409, 210.297, 210.2708, 210.1831, 
    210.1065,
  209.9483, 209.9457, 209.9653, 209.9683, 209.9903, 210.0147, 210.0289, 
    210.0285, 210.0892, 210.1824, 210.2725, 210.3272, 210.2936, 210.2182, 
    210.1635,
  209.9436, 209.9361, 209.9599, 209.965, 209.9922, 210.0413, 210.0419, 
    210.0539, 210.1156, 210.1693, 210.2476, 210.3016, 210.2719, 210.2354, 
    210.2101,
  209.9459, 209.9323, 209.9467, 209.9924, 210.0511, 210.0715, 210.0688, 
    210.0566, 210.1048, 210.1423, 210.2145, 210.2938, 210.2816, 210.268, 
    210.2448,
  209.0096, 208.9784, 208.9358, 208.8984, 208.8666, 208.8589, 208.863, 
    208.8919, 208.9265, 208.9371, 208.9565, 208.9447, 208.8982, 208.8391, 
    208.7523,
  209.0148, 209.0131, 208.9648, 208.9232, 208.8925, 208.8898, 208.8962, 
    208.9256, 208.9438, 208.9594, 208.9831, 208.957, 208.9463, 208.9076, 
    208.8248,
  209.0242, 209.0417, 209.001, 208.983, 208.96, 208.9586, 208.9581, 208.9885, 
    208.9877, 209.0034, 209.0112, 208.9867, 209.0013, 208.9609, 208.9117,
  209.0415, 209.0686, 209.037, 209.0227, 209.0068, 209.0063, 209.0142, 
    209.0368, 209.0328, 209.0485, 209.0347, 209.0352, 209.0443, 209.0033, 
    208.9862,
  209.075, 209.0922, 209.0809, 209.074, 209.0671, 209.0633, 209.068, 
    209.0762, 209.0839, 209.1047, 209.1006, 209.1291, 209.141, 209.1211, 
    209.0936,
  209.1171, 209.1275, 209.1439, 209.1318, 209.11, 209.1036, 209.116, 
    209.1327, 209.1455, 209.1696, 209.1916, 209.2246, 209.2346, 209.2179, 
    209.1861,
  209.1749, 209.1725, 209.1812, 209.164, 209.1626, 209.1534, 209.1535, 
    209.1733, 209.1947, 209.2404, 209.279, 209.3132, 209.3256, 209.33, 209.307,
  209.2193, 209.2186, 209.2188, 209.2034, 209.1956, 209.1782, 209.1837, 
    209.2026, 209.2462, 209.3075, 209.3497, 209.3858, 209.4011, 209.4143, 
    209.4056,
  209.2625, 209.2621, 209.2646, 209.234, 209.2168, 209.2271, 209.2412, 
    209.2569, 209.3062, 209.36, 209.4188, 209.4538, 209.4602, 209.4804, 
    209.4954,
  209.3143, 209.2998, 209.3073, 209.3157, 209.3182, 209.336, 209.3273, 
    209.3281, 209.3912, 209.44, 209.4952, 209.5233, 209.5278, 209.5483, 
    209.5615,
  207.6964, 207.6329, 207.5654, 207.522, 207.4814, 207.4348, 207.3878, 
    207.3264, 207.2569, 207.1851, 207.1093, 207.0379, 206.9628, 206.8963, 
    206.8461,
  207.7677, 207.709, 207.6584, 207.6216, 207.5679, 207.5203, 207.475, 
    207.4189, 207.3557, 207.2847, 207.2193, 207.1541, 207.0749, 206.9932, 
    206.9362,
  207.8381, 207.7867, 207.7298, 207.6803, 207.6253, 207.5976, 207.5603, 
    207.5203, 207.4773, 207.4203, 207.3485, 207.271, 207.1743, 207.0848, 
    207.013,
  207.9193, 207.8725, 207.8087, 207.7395, 207.6907, 207.6586, 207.6314, 
    207.6036, 207.5617, 207.5005, 207.4344, 207.3623, 207.2748, 207.1866, 
    207.1048,
  208.0185, 207.9387, 207.874, 207.8143, 207.7673, 207.7241, 207.693, 
    207.6633, 207.6262, 207.5672, 207.5073, 207.4371, 207.3569, 207.2649, 
    207.1773,
  208.1236, 208.0273, 207.9696, 207.9004, 207.8189, 207.7878, 207.7662, 
    207.7288, 207.6872, 207.6386, 207.5794, 207.5111, 207.4352, 207.3357, 
    207.2242,
  208.2414, 208.1364, 208.0585, 207.9778, 207.9189, 207.8748, 207.8446, 
    207.8164, 207.7692, 207.7179, 207.6579, 207.5844, 207.4981, 207.3941, 
    207.2814,
  208.3688, 208.262, 208.1729, 208.0981, 208.0434, 207.9784, 207.939, 
    207.8978, 207.8446, 207.7976, 207.7381, 207.6738, 207.5871, 207.4814, 
    207.3741,
  208.4828, 208.3781, 208.2908, 208.1808, 208.11, 208.0739, 208.0488, 
    207.9899, 207.9294, 207.8751, 207.814, 207.7499, 207.649, 207.5426, 
    207.4403,
  208.6064, 208.4741, 208.3866, 208.2938, 208.2336, 208.195, 208.15, 
    208.0769, 208.029, 207.9633, 207.8914, 207.8081, 207.7022, 207.6095, 
    207.5352,
  206.9865, 206.9234, 206.8229, 206.7269, 206.6501, 206.5788, 206.5251, 
    206.4713, 206.4088, 206.335, 206.2453, 206.1628, 206.0931, 206.0366, 
    205.9873,
  207.1418, 207.0947, 206.9944, 206.9042, 206.8098, 206.7266, 206.6568, 
    206.5816, 206.511, 206.4261, 206.3379, 206.2553, 206.1836, 206.1196, 
    206.0581,
  207.3741, 207.3035, 207.1991, 207.0938, 206.9858, 206.8882, 206.8041, 
    206.7218, 206.6511, 206.5678, 206.476, 206.3818, 206.2979, 206.2265, 
    206.1665,
  207.5804, 207.5093, 207.4343, 207.3294, 207.2085, 207.0948, 206.9979, 
    206.9097, 206.827, 206.7429, 206.654, 206.5605, 206.473, 206.3974, 
    206.3311,
  207.782, 207.7034, 207.6416, 207.5566, 207.4531, 207.3292, 207.2214, 
    207.1255, 207.0373, 206.9594, 206.8655, 206.769, 206.6721, 206.5825, 
    206.5034,
  207.9292, 207.8745, 207.8313, 207.7639, 207.67, 207.5756, 207.4839, 
    207.3883, 207.2863, 207.1875, 207.0928, 206.9922, 206.8838, 206.7938, 
    206.714,
  208.0762, 208.0417, 207.9931, 207.9258, 207.8664, 207.7966, 207.728, 
    207.6501, 207.555, 207.447, 207.3383, 207.2265, 207.1198, 207.0098, 
    206.9178,
  208.2123, 208.1731, 208.1187, 208.0678, 208.0459, 207.9898, 207.9382, 
    207.8757, 207.7956, 207.6813, 207.5627, 207.4479, 207.3318, 207.2143, 
    207.1191,
  208.3326, 208.313, 208.2943, 208.23, 208.1699, 208.1421, 208.1228, 
    208.0578, 207.9816, 207.901, 207.8001, 207.6822, 207.5656, 207.4433, 
    207.3284,
  208.4693, 208.4325, 208.4097, 208.3741, 208.3496, 208.3368, 208.2865, 
    208.2198, 208.1642, 208.0779, 208.0092, 207.9188, 207.7989, 207.6604, 
    207.5322,
  206.2875, 206.2523, 206.23, 206.2272, 206.2304, 206.2388, 206.2509, 
    206.2685, 206.2904, 206.3099, 206.3166, 206.3251, 206.3238, 206.3244, 
    206.3195,
  206.3673, 206.3448, 206.3148, 206.2849, 206.2746, 206.2734, 206.278, 
    206.2914, 206.3106, 206.3282, 206.3423, 206.3548, 206.3702, 206.3742, 
    206.3736,
  206.4942, 206.4636, 206.4195, 206.3793, 206.3397, 206.3281, 206.3241, 
    206.3207, 206.3308, 206.3476, 206.3606, 206.3773, 206.3924, 206.4117, 
    206.4319,
  206.6398, 206.6081, 206.569, 206.5074, 206.4632, 206.4271, 206.4137, 
    206.3948, 206.3793, 206.3767, 206.385, 206.3955, 206.4124, 206.4319, 
    206.4538,
  206.8427, 206.7816, 206.7318, 206.6684, 206.6232, 206.5695, 206.5308, 
    206.4937, 206.4698, 206.4494, 206.4388, 206.4356, 206.4411, 206.4459, 
    206.4635,
  207.0598, 206.9973, 206.9476, 206.8808, 206.8035, 206.7457, 206.6953, 
    206.6478, 206.6009, 206.5598, 206.5323, 206.5075, 206.4914, 206.487, 
    206.4936,
  207.3122, 207.2424, 207.1721, 207.0917, 207.027, 206.9558, 206.8902, 
    206.8365, 206.7776, 206.7234, 206.6767, 206.6321, 206.5972, 206.5809, 
    206.5802,
  207.5916, 207.5059, 207.4158, 207.3336, 207.2959, 207.2259, 207.1587, 
    207.0753, 207.0009, 206.9395, 206.8764, 206.8117, 206.7753, 206.7444, 
    206.74,
  207.8291, 207.7628, 207.7012, 207.5914, 207.5153, 207.484, 207.4496, 
    207.3741, 207.2816, 207.2086, 207.1411, 207.0716, 207.0137, 206.9518, 
    206.9331,
  208.0502, 207.9634, 207.9184, 207.8603, 207.8101, 207.796, 207.7295, 
    207.6585, 207.6061, 207.5179, 207.4427, 207.3787, 207.3257, 207.2487, 
    207.203,
  206.3648, 206.3305, 206.3165, 206.3276, 206.3317, 206.3323, 206.34, 
    206.3563, 206.389, 206.4167, 206.4516, 206.4816, 206.5045, 206.5204, 
    206.5037,
  206.4511, 206.4463, 206.4167, 206.398, 206.388, 206.3722, 206.3787, 
    206.3972, 206.4274, 206.4574, 206.5001, 206.5262, 206.5439, 206.5601, 
    206.5505,
  206.5793, 206.5604, 206.5108, 206.4906, 206.4716, 206.4542, 206.4551, 
    206.4692, 206.4878, 206.5099, 206.5406, 206.5593, 206.5888, 206.6081, 
    206.6024,
  206.7109, 206.6731, 206.6405, 206.6279, 206.6076, 206.5823, 206.5716, 
    206.5759, 206.5775, 206.5886, 206.5995, 206.6137, 206.6223, 206.6333, 
    206.6467,
  206.8983, 206.8366, 206.7905, 206.7725, 206.7663, 206.7461, 206.7246, 
    206.7073, 206.6932, 206.6841, 206.6788, 206.6844, 206.6796, 206.6954, 
    206.7027,
  207.1243, 207.0587, 207.0097, 206.9847, 206.941, 206.9076, 206.8922, 
    206.8716, 206.859, 206.836, 206.8125, 206.7933, 206.786, 206.7916, 
    206.7824,
  207.3559, 207.3056, 207.2511, 207.2051, 207.1638, 207.1187, 207.073, 
    207.0486, 207.0384, 207.021, 206.9905, 206.9563, 206.9274, 206.9212, 
    206.9012,
  207.5987, 207.5698, 207.5044, 207.4581, 207.4534, 207.3792, 207.313, 
    207.2658, 207.2394, 207.241, 207.2271, 207.181, 207.1314, 207.1092, 
    207.0953,
  207.8562, 207.8145, 207.7931, 207.7341, 207.6667, 207.6589, 207.6241, 
    207.5469, 207.4853, 207.4618, 207.469, 207.445, 207.4016, 207.352, 
    207.3304,
  208.1657, 208.074, 208.0285, 208.0057, 207.9848, 207.9982, 207.9495, 
    207.8634, 207.8254, 207.7586, 207.7459, 207.7455, 207.7221, 207.6848, 
    207.6492,
  208.0751, 208.091, 208.0826, 208.0997, 208.0984, 208.0925, 208.1129, 
    208.1249, 208.1422, 208.1555, 208.1936, 208.2294, 208.2513, 208.2653, 
    208.2712,
  208.2131, 208.2414, 208.222, 208.2363, 208.2417, 208.2372, 208.2513, 
    208.2638, 208.2802, 208.2999, 208.325, 208.3567, 208.3789, 208.3938, 
    208.4041,
  208.3699, 208.3957, 208.3844, 208.4079, 208.4036, 208.4175, 208.4351, 
    208.451, 208.4699, 208.4835, 208.5144, 208.541, 208.5603, 208.5762, 
    208.5901,
  208.5206, 208.5309, 208.5402, 208.5615, 208.5687, 208.5917, 208.6167, 
    208.6383, 208.659, 208.6719, 208.6987, 208.7205, 208.7451, 208.758, 
    208.7769,
  208.7289, 208.7315, 208.7471, 208.7734, 208.8023, 208.8264, 208.8394, 
    208.8681, 208.8927, 208.9034, 208.9129, 208.9217, 208.9466, 208.959, 
    208.9619,
  208.9826, 208.9776, 209.0135, 209.0432, 209.0502, 209.0643, 209.0823, 
    209.1034, 209.1268, 209.1346, 209.1369, 209.1381, 209.1479, 209.1492, 
    209.1504,
  209.2526, 209.2464, 209.2815, 209.2998, 209.3517, 209.3713, 209.3724, 
    209.3861, 209.3957, 209.4085, 209.4057, 209.3954, 209.3866, 209.3736, 
    209.3762,
  209.4854, 209.5036, 209.5209, 209.5633, 209.6522, 209.6747, 209.692, 
    209.6924, 209.6895, 209.7012, 209.7029, 209.6878, 209.6644, 209.6453, 
    209.6406,
  209.6724, 209.7025, 209.7468, 209.7852, 209.8276, 209.9225, 209.9876, 
    209.9785, 209.977, 209.979, 209.9984, 209.9898, 209.9687, 209.9447, 
    209.9304,
  209.836, 209.8566, 209.8902, 209.9595, 210.0423, 210.1456, 210.1889, 
    210.1974, 210.2372, 210.2278, 210.2374, 210.251, 210.2436, 210.2378, 
    210.2248,
  207.8632, 207.882, 207.8657, 207.902, 207.9539, 207.9869, 208.0081, 
    208.0166, 208.0242, 208.0368, 208.0574, 208.0809, 208.0948, 208.0991, 
    208.1131,
  207.9619, 208.0021, 208.0027, 208.0474, 208.0972, 208.1243, 208.1467, 
    208.1556, 208.1701, 208.176, 208.1882, 208.2098, 208.228, 208.2609, 
    208.2872,
  208.1766, 208.2245, 208.2151, 208.2316, 208.2593, 208.2979, 208.3275, 
    208.3456, 208.3641, 208.3787, 208.3912, 208.3943, 208.4122, 208.4374, 
    208.464,
  208.3668, 208.3849, 208.377, 208.3941, 208.4321, 208.4904, 208.5208, 
    208.5517, 208.579, 208.59, 208.6034, 208.6061, 208.6237, 208.6327, 
    208.6546,
  208.6365, 208.6188, 208.6017, 208.6214, 208.6848, 208.7483, 208.8007, 
    208.8581, 208.8811, 208.8811, 208.8747, 208.8655, 208.87, 208.8823, 
    208.8885,
  208.9228, 208.8783, 208.8822, 208.8972, 208.9349, 208.9835, 209.0385, 
    209.0806, 209.1154, 209.1456, 209.1538, 209.1458, 209.1408, 209.1395, 
    209.1489,
  209.1519, 209.1351, 209.1337, 209.1464, 209.2222, 209.2979, 209.3575, 
    209.401, 209.4335, 209.4635, 209.4651, 209.4591, 209.46, 209.4554, 
    209.4552,
  209.3471, 209.3641, 209.3832, 209.4046, 209.4862, 209.5537, 209.6262, 
    209.6803, 209.7108, 209.7485, 209.7744, 209.7709, 209.7548, 209.7429, 
    209.7414,
  209.4964, 209.5451, 209.6064, 209.6176, 209.6345, 209.7356, 209.8214, 
    209.8653, 209.9023, 209.9367, 209.9809, 209.9942, 209.9816, 209.9501, 
    209.9448,
  209.6555, 209.7079, 209.7411, 209.7917, 209.8284, 209.8976, 209.9268, 
    209.9367, 210.0071, 210.0442, 210.0865, 210.1346, 210.137, 210.1241, 
    210.1161,
  207.5036, 207.5314, 207.5365, 207.5577, 207.5883, 207.6165, 207.6447, 
    207.6679, 207.6851, 207.689, 207.6904, 207.6812, 207.6671, 207.6522, 
    207.6409,
  207.6172, 207.6827, 207.6652, 207.69, 207.7286, 207.7506, 207.7863, 
    207.8122, 207.8377, 207.8401, 207.8352, 207.8255, 207.8268, 207.824, 
    207.8132,
  207.8214, 207.8654, 207.8533, 207.8839, 207.9085, 207.9472, 207.9935, 
    208.0433, 208.0804, 208.0957, 208.1028, 208.0937, 208.0718, 208.0341, 
    207.9915,
  208.021, 208.0078, 208.0184, 208.0458, 208.0752, 208.135, 208.1828, 
    208.2404, 208.2913, 208.3206, 208.3426, 208.3504, 208.3241, 208.2788, 
    208.2255,
  208.2295, 208.2099, 208.2429, 208.2832, 208.3331, 208.3716, 208.4187, 
    208.4887, 208.556, 208.6133, 208.6445, 208.6548, 208.632, 208.5808, 
    208.5104,
  208.4832, 208.4588, 208.485, 208.5211, 208.5526, 208.6039, 208.6633, 
    208.7393, 208.8281, 208.8955, 208.9365, 208.9631, 208.9464, 208.8972, 
    208.8141,
  208.7509, 208.7369, 208.7518, 208.766, 208.8333, 208.892, 208.9408, 
    209.0192, 209.1064, 209.1845, 209.2244, 209.2305, 209.2043, 209.1659, 
    209.1182,
  209.0134, 209.018, 209.0489, 209.0509, 209.1031, 209.1432, 209.2141, 
    209.2663, 209.3257, 209.3996, 209.4507, 209.4561, 209.4249, 209.3757, 
    209.3169,
  209.269, 209.2905, 209.333, 209.311, 209.3203, 209.3866, 209.4587, 
    209.4799, 209.5132, 209.542, 209.5956, 209.6057, 209.584, 209.5323, 
    209.4743,
  209.5216, 209.5234, 209.5412, 209.5463, 209.5724, 209.5984, 209.6197, 
    209.621, 209.6657, 209.6761, 209.6949, 209.7033, 209.6805, 209.6353, 
    209.5705,
  207.1199, 207.145, 207.1301, 207.112, 207.0784, 207.077, 207.1043, 
    207.1304, 207.1456, 207.1452, 207.1496, 207.1619, 207.202, 207.2318, 
    207.25,
  207.2702, 207.2619, 207.2116, 207.2099, 207.186, 207.1815, 207.1988, 
    207.2217, 207.2394, 207.2299, 207.2284, 207.232, 207.2695, 207.3051, 
    207.3358,
  207.4235, 207.38, 207.3479, 207.3517, 207.3091, 207.2824, 207.2889, 
    207.3254, 207.3591, 207.3608, 207.3696, 207.3894, 207.4225, 207.4571, 
    207.4954,
  207.5309, 207.4828, 207.4839, 207.4634, 207.4059, 207.3983, 207.4004, 
    207.4404, 207.4807, 207.4957, 207.5108, 207.5346, 207.5671, 207.6171, 
    207.6666,
  207.6714, 207.634, 207.6018, 207.5786, 207.5729, 207.5772, 207.578, 
    207.6063, 207.6422, 207.6673, 207.6822, 207.7167, 207.7633, 207.8307, 
    207.894,
  207.8673, 207.8316, 207.7853, 207.7699, 207.7499, 207.745, 207.7569, 
    207.7795, 207.8196, 207.8551, 207.8852, 207.9195, 207.9719, 208.0466, 
    208.1218,
  208.093, 208.0776, 208.0243, 207.9722, 207.956, 207.9585, 207.95, 207.9613, 
    207.9913, 208.0323, 208.0711, 208.1144, 208.1907, 208.2905, 208.3828,
  208.308, 208.3146, 208.2661, 208.2174, 208.202, 208.176, 208.1599, 
    208.1515, 208.1603, 208.2127, 208.2585, 208.3227, 208.418, 208.5208, 
    208.6227,
  208.5, 208.5115, 208.4915, 208.4496, 208.4039, 208.3946, 208.394, 208.3779, 
    208.3712, 208.3957, 208.4538, 208.5405, 208.6518, 208.7594, 208.8559,
  208.7019, 208.6915, 208.6661, 208.6401, 208.631, 208.6374, 208.6233, 
    208.5834, 208.5977, 208.6245, 208.6774, 208.7807, 208.8873, 208.9942, 
    209.0779,
  207.1485, 207.1393, 207.0935, 207.089, 207.1419, 207.1476, 207.1269, 
    207.0736, 207.0467, 207.0271, 206.9843, 206.928, 206.9303, 206.943, 
    206.9547,
  207.1697, 207.1952, 207.17, 207.1732, 207.2005, 207.1869, 207.1794, 
    207.1209, 207.1134, 207.1279, 207.1057, 207.0393, 206.995, 206.9715, 
    206.9869,
  207.2141, 207.2669, 207.2721, 207.2778, 207.2831, 207.3003, 207.3169, 
    207.2769, 207.269, 207.2561, 207.2262, 207.1586, 207.0911, 207.0627, 
    207.0712,
  207.2977, 207.3643, 207.3711, 207.3633, 207.3763, 207.39, 207.3898, 
    207.3573, 207.3325, 207.304, 207.2686, 207.2183, 207.1643, 207.1402, 
    207.1375,
  207.4039, 207.4135, 207.4152, 207.4341, 207.4381, 207.4337, 207.4305, 
    207.4373, 207.4285, 207.3968, 207.3461, 207.3008, 207.2655, 207.2423, 
    207.2265,
  207.5363, 207.5262, 207.5597, 207.5835, 207.5505, 207.5412, 207.551, 
    207.5576, 207.5463, 207.5152, 207.4716, 207.4318, 207.4102, 207.3908, 
    207.3715,
  207.6471, 207.6592, 207.6779, 207.6802, 207.6901, 207.6866, 207.6705, 
    207.6778, 207.6767, 207.6616, 207.6315, 207.5982, 207.5817, 207.5648, 
    207.5426,
  207.7089, 207.7368, 207.7612, 207.7911, 207.8361, 207.8467, 207.855, 
    207.8707, 207.8539, 207.8489, 207.8242, 207.7946, 207.7652, 207.7256, 
    207.6949,
  207.7745, 207.7836, 207.8295, 207.8583, 207.8681, 207.9337, 207.989, 
    208.0054, 208.0044, 207.9994, 207.996, 207.9615, 207.9194, 207.8666, 
    207.8234,
  207.868, 207.8548, 207.875, 207.9149, 207.9541, 208.0388, 208.0855, 
    208.0881, 208.1108, 208.1024, 208.0939, 208.0868, 208.049, 207.9955, 
    207.9418,
  207.275, 207.236, 207.2132, 207.2017, 207.1835, 207.1708, 207.1572, 
    207.1562, 207.1701, 207.1912, 207.213, 207.2307, 207.2575, 207.2902, 
    207.3329,
  207.3722, 207.3809, 207.3531, 207.3165, 207.2956, 207.2819, 207.2669, 
    207.2579, 207.2488, 207.2499, 207.2563, 207.2541, 207.2527, 207.2509, 
    207.251,
  207.4926, 207.5059, 207.476, 207.4591, 207.4386, 207.4186, 207.3967, 
    207.3708, 207.3473, 207.334, 207.3264, 207.3141, 207.298, 207.2758, 
    207.2601,
  207.6045, 207.5996, 207.595, 207.5904, 207.5729, 207.5531, 207.5308, 
    207.5042, 207.477, 207.4485, 207.4245, 207.3987, 207.3746, 207.3468, 
    207.3357,
  207.7443, 207.7234, 207.7163, 207.7014, 207.6986, 207.694, 207.6755, 
    207.6484, 207.6068, 207.5697, 207.5357, 207.5031, 207.4743, 207.4398, 
    207.418,
  207.8883, 207.8653, 207.8503, 207.8423, 207.8164, 207.8091, 207.7995, 
    207.7836, 207.7459, 207.7034, 207.6634, 207.6184, 207.5761, 207.5298, 
    207.5,
  208.0181, 207.9999, 207.976, 207.9481, 207.9434, 207.9344, 207.9213, 
    207.9146, 207.884, 207.8517, 207.8126, 207.7643, 207.7113, 207.6527, 
    207.5972,
  208.1181, 208.1082, 208.0807, 208.0478, 208.0644, 208.0531, 208.0492, 
    208.0346, 208.0037, 207.9858, 207.9522, 207.9211, 207.8666, 207.8023, 
    207.7313,
  208.2435, 208.235, 208.2236, 208.1936, 208.157, 208.1611, 208.1824, 
    208.1714, 208.1475, 208.118, 208.0959, 208.0712, 208.032, 207.9684, 
    207.8903,
  208.3921, 208.3567, 208.3295, 208.3174, 208.3196, 208.3585, 208.3562, 
    208.2986, 208.2924, 208.2659, 208.2264, 208.206, 208.1715, 208.121, 
    208.0462,
  207.949, 207.9116, 207.8504, 207.8243, 207.7755, 207.7272, 207.6839, 
    207.6584, 207.6281, 207.5914, 207.5522, 207.5158, 207.4923, 207.4733, 
    207.4641,
  208.0845, 208.0538, 207.9887, 207.9295, 207.8662, 207.8056, 207.7575, 
    207.7108, 207.681, 207.6494, 207.6118, 207.5678, 207.5274, 207.4958, 
    207.4748,
  208.1995, 208.1732, 208.1079, 208.0378, 207.971, 207.9091, 207.8481, 
    207.7969, 207.7552, 207.7135, 207.6746, 207.6307, 207.5824, 207.5437, 
    207.5118,
  208.2824, 208.2666, 208.2022, 208.1365, 208.0799, 208.0156, 207.9604, 
    207.9162, 207.8553, 207.802, 207.7505, 207.7075, 207.6589, 207.6149, 
    207.5763,
  208.3444, 208.3199, 208.2555, 208.1998, 208.1576, 208.1111, 208.0682, 
    208.0189, 207.9611, 207.9062, 207.8388, 207.7794, 207.736, 207.6929, 
    207.6505,
  208.3887, 208.352, 208.3002, 208.27, 208.2279, 208.1866, 208.1488, 
    208.1125, 208.0631, 208.0087, 207.937, 207.8705, 207.815, 207.7727, 
    207.7329,
  208.4851, 208.4337, 208.368, 208.3188, 208.3002, 208.2662, 208.229, 
    208.1938, 208.1531, 208.1097, 208.0516, 207.9704, 207.8967, 207.8406, 
    207.8015,
  208.5504, 208.503, 208.4458, 208.3871, 208.3694, 208.3374, 208.3031, 
    208.2669, 208.218, 208.188, 208.1384, 208.0763, 207.9907, 207.9125, 
    207.864,
  208.5922, 208.5519, 208.5406, 208.4798, 208.4122, 208.3963, 208.3877, 
    208.3554, 208.3136, 208.263, 208.2185, 208.1721, 208.0985, 208.0173, 
    207.942,
  208.6463, 208.5925, 208.5634, 208.5275, 208.5046, 208.5132, 208.4877, 
    208.4324, 208.414, 208.3662, 208.3167, 208.2716, 208.2198, 208.1514, 
    208.0644,
  207.8233, 207.7934, 207.7327, 207.694, 207.6718, 207.6491, 207.5988, 
    207.5483, 207.5036, 207.4698, 207.4382, 207.4131, 207.3868, 207.345, 
    207.3002,
  207.8785, 207.883, 207.8242, 207.7707, 207.7187, 207.6803, 207.659, 
    207.6281, 207.5704, 207.508, 207.4698, 207.4316, 207.3991, 207.3567, 
    207.3078,
  207.9435, 207.9658, 207.9306, 207.8856, 207.8053, 207.7596, 207.7354, 
    207.6849, 207.6273, 207.5676, 207.5157, 207.4593, 207.4096, 207.3649, 
    207.3136,
  208.0255, 208.0287, 207.9958, 207.971, 207.9176, 207.8611, 207.8272, 
    207.775, 207.7085, 207.6334, 207.5658, 207.5078, 207.4555, 207.4239, 
    207.367,
  208.1321, 208.0871, 208.045, 208.0288, 208.0117, 207.9686, 207.9271, 
    207.8772, 207.8014, 207.7173, 207.6514, 207.5946, 207.528, 207.4892, 
    207.4362,
  208.2311, 208.1736, 208.1293, 208.1132, 208.0861, 208.0447, 207.9918, 
    207.9545, 207.8895, 207.8106, 207.7264, 207.6636, 207.5965, 207.5324, 
    207.4733,
  208.2977, 208.2755, 208.2258, 208.1982, 208.1727, 208.1267, 208.0541, 
    208.0107, 207.9585, 207.8904, 207.8026, 207.7188, 207.6375, 207.5592, 
    207.4822,
  208.3411, 208.3625, 208.3349, 208.301, 208.2867, 208.2363, 208.1747, 
    208.1023, 208.0332, 207.9775, 207.8944, 207.7952, 207.6835, 207.5802, 
    207.4837,
  208.3837, 208.4159, 208.4453, 208.4124, 208.3522, 208.3405, 208.3093, 
    208.2449, 208.1679, 208.0825, 208.0129, 207.8959, 207.7802, 207.6464, 
    207.5298,
  208.4617, 208.4773, 208.505, 208.5089, 208.4911, 208.4959, 208.4451, 
    208.3646, 208.3128, 208.22, 208.1486, 208.0415, 207.9053, 207.7669, 
    207.6216,
  206.7876, 206.7607, 206.7154, 206.6869, 206.6678, 206.6451, 206.6182, 
    206.5916, 206.5772, 206.5488, 206.5051, 206.4886, 206.4494, 206.4083, 
    206.3604,
  206.7874, 206.7538, 206.6734, 206.6382, 206.6171, 206.5853, 206.5508, 
    206.5054, 206.4546, 206.4062, 206.3677, 206.3423, 206.3039, 206.2695, 
    206.2416,
  206.801, 206.7428, 206.64, 206.5985, 206.5479, 206.5099, 206.4717, 
    206.4138, 206.3493, 206.3022, 206.2633, 206.2212, 206.1775, 206.1471, 
    206.12,
  206.7943, 206.718, 206.6274, 206.57, 206.4983, 206.4518, 206.4058, 
    206.3562, 206.3012, 206.239, 206.1808, 206.1221, 206.0761, 206.0432, 
    206.0038,
  206.8375, 206.7364, 206.6436, 206.5716, 206.5108, 206.4485, 206.3796, 
    206.3195, 206.2594, 206.2011, 206.1414, 206.0808, 206.015, 205.9468, 
    205.8809,
  206.9251, 206.8, 206.7084, 206.6414, 206.5426, 206.4731, 206.4072, 
    206.3324, 206.2574, 206.1915, 206.1207, 206.036, 205.9435, 205.8418, 
    205.7573,
  207.0383, 206.9231, 206.807, 206.72, 206.6536, 206.5836, 206.4931, 
    206.4042, 206.3057, 206.2223, 206.1415, 206.0467, 205.9321, 205.8213, 
    205.708,
  207.1328, 207.0525, 206.9285, 206.8383, 206.7982, 206.7116, 206.6286, 
    206.5241, 206.3989, 206.3052, 206.2177, 206.1185, 205.995, 205.8621, 
    205.7375,
  207.2426, 207.1622, 207.0664, 206.9583, 206.8595, 206.8353, 206.795, 
    206.6937, 206.5725, 206.4392, 206.3408, 206.2431, 206.1197, 205.9766, 
    205.835,
  207.3809, 207.2655, 207.1851, 207.1068, 207.036, 207.0301, 206.9629, 
    206.848, 206.7643, 206.6167, 206.498, 206.4015, 206.2787, 206.1323, 
    205.9678,
  206.5122, 206.5005, 206.4841, 206.4633, 206.4365, 206.4305, 206.4155, 
    206.4093, 206.3985, 206.373, 206.3404, 206.3163, 206.2958, 206.2723, 
    206.2486,
  206.4227, 206.4379, 206.3958, 206.35, 206.326, 206.3156, 206.3106, 
    206.3031, 206.29, 206.2677, 206.2495, 206.2263, 206.2028, 206.1795, 
    206.1494,
  206.3876, 206.3886, 206.3233, 206.2829, 206.2504, 206.2326, 206.2282, 
    206.2215, 206.2082, 206.1833, 206.1657, 206.1488, 206.1268, 206.1089, 
    206.0776,
  206.3547, 206.3377, 206.2864, 206.248, 206.1957, 206.1725, 206.1595, 
    206.1507, 206.1335, 206.1001, 206.0723, 206.0518, 206.0412, 206.0339, 
    206.013,
  206.3319, 206.2796, 206.2262, 206.1966, 206.1629, 206.1414, 206.1202, 
    206.1041, 206.0773, 206.0416, 206.0067, 205.9746, 205.9582, 205.9496, 
    205.9353,
  206.3687, 206.3183, 206.2672, 206.2136, 206.1436, 206.1107, 206.0883, 
    206.0685, 206.0433, 206.0051, 205.9534, 205.9085, 205.8756, 205.8601, 
    205.8499,
  206.4525, 206.3896, 206.3037, 206.2353, 206.1761, 206.1272, 206.0875, 
    206.0574, 206.0263, 205.9919, 205.9296, 205.8729, 205.824, 205.7913, 
    205.7724,
  206.5298, 206.46, 206.3802, 206.3154, 206.2671, 206.2023, 206.1493, 
    206.0914, 206.0425, 206.0034, 205.9367, 205.8665, 205.7959, 205.7445, 
    205.7099,
  206.6269, 206.6105, 206.5496, 206.4527, 206.3651, 206.3189, 206.2593, 
    206.1799, 206.1065, 206.0406, 205.9743, 205.8941, 205.8113, 205.7382, 
    205.6772,
  206.7492, 206.712, 206.651, 206.5965, 206.5366, 206.4996, 206.4081, 
    206.2873, 206.2173, 206.1183, 206.0352, 205.9433, 205.8509, 205.7587, 
    205.6811,
  206.6533, 206.6513, 206.6474, 206.6392, 206.6279, 206.5905, 206.5714, 
    206.5444, 206.5078, 206.4624, 206.4138, 206.369, 206.3207, 206.2827, 
    206.2409,
  206.4424, 206.4797, 206.4515, 206.4387, 206.4059, 206.356, 206.339, 
    206.3351, 206.334, 206.3145, 206.2788, 206.2416, 206.1976, 206.1617, 
    206.1173,
  206.319, 206.3303, 206.2902, 206.2831, 206.2309, 206.194, 206.177, 
    206.1783, 206.1764, 206.1367, 206.1028, 206.0679, 206.0402, 206.0186, 
    206.0004,
  206.1692, 206.1764, 206.159, 206.1515, 206.1029, 206.0713, 206.0435, 
    206.0272, 206.0165, 205.9957, 205.9714, 205.9374, 205.9136, 205.8913, 
    205.8702,
  206.0836, 206.0338, 205.9965, 206.0235, 206.0521, 206.0567, 206.0572, 
    206.0485, 206.0252, 205.9828, 205.9261, 205.8805, 205.8553, 205.8212, 
    205.786,
  206.0292, 205.9605, 205.9521, 205.9816, 205.9704, 205.9852, 206.005, 
    205.9949, 205.9763, 205.9453, 205.9061, 205.867, 205.8447, 205.8211, 
    205.7731,
  206.0098, 205.9654, 205.9386, 205.9218, 205.895, 205.881, 205.856, 
    205.8514, 205.8699, 205.8933, 205.8784, 205.8323, 205.7894, 205.7505, 
    205.7158,
  206.0132, 205.9675, 205.9138, 205.8774, 205.8658, 205.8549, 205.8585, 
    205.8282, 205.797, 205.8041, 205.794, 205.7639, 205.7283, 205.6979, 
    205.6858,
  205.9956, 205.9838, 205.9628, 205.8795, 205.8096, 205.8354, 205.8575, 
    205.8217, 205.7643, 205.7629, 205.7836, 205.7721, 205.7365, 205.6867, 
    205.6676,
  206.0538, 206.0382, 205.9919, 205.9759, 205.9572, 205.98, 205.9694, 
    205.9073, 205.8652, 205.8217, 205.8093, 205.7947, 205.7707, 205.7419, 
    205.7165,
  207.6517, 207.6042, 207.5621, 207.5446, 207.5284, 207.5089, 207.4965, 
    207.4706, 207.4237, 207.362, 207.3047, 207.2565, 207.2118, 207.1593, 
    207.0984,
  207.3331, 207.3179, 207.252, 207.2168, 207.1989, 207.1766, 207.1519, 
    207.1212, 207.0934, 207.0623, 207.0337, 207.0047, 206.968, 206.9315, 
    206.8793,
  207.151, 207.0993, 207.0228, 206.9963, 206.9621, 206.9305, 206.9021, 
    206.8713, 206.849, 206.8294, 206.8092, 206.7774, 206.742, 206.6935, 
    206.6417,
  206.9967, 206.9273, 206.8713, 206.8384, 206.7896, 206.7551, 206.7267, 
    206.7025, 206.687, 206.6706, 206.6488, 206.6082, 206.5535, 206.5041, 
    206.4688,
  206.9364, 206.8355, 206.7757, 206.7361, 206.6904, 206.6509, 206.6203, 
    206.6025, 206.5882, 206.57, 206.5378, 206.4804, 206.4299, 206.3938, 
    206.3638,
  206.9249, 206.814, 206.7671, 206.707, 206.6222, 206.5797, 206.5576, 
    206.5418, 206.5253, 206.5035, 206.4714, 206.4215, 206.3716, 206.3402, 
    206.3219,
  206.938, 206.8391, 206.7615, 206.6644, 206.6072, 206.5536, 206.5176, 
    206.5011, 206.479, 206.469, 206.4479, 206.4146, 206.3754, 206.3574, 
    206.3452,
  206.9697, 206.8952, 206.7947, 206.7006, 206.6403, 206.5726, 206.5376, 
    206.5032, 206.4716, 206.4604, 206.4384, 206.4194, 206.3978, 206.3667, 
    206.348,
  207.0465, 206.9851, 206.9021, 206.7741, 206.6434, 206.6259, 206.6026, 
    206.5558, 206.519, 206.4811, 206.4673, 206.4612, 206.4585, 206.4222, 
    206.3746,
  207.1852, 207.0706, 206.9738, 206.8696, 206.7988, 206.787, 206.7271, 
    206.6507, 206.6323, 206.583, 206.5349, 206.5369, 206.5462, 206.5319, 
    206.5054,
  207.8778, 207.802, 207.7245, 207.6691, 207.6263, 207.5839, 207.5513, 
    207.5233, 207.4964, 207.4784, 207.4603, 207.4498, 207.4462, 207.4285, 
    207.4301,
  207.6888, 207.6555, 207.5348, 207.4458, 207.3778, 207.3204, 207.2858, 
    207.2512, 207.2166, 207.1875, 207.1627, 207.1565, 207.1478, 207.1335, 
    207.1208,
  207.5899, 207.5135, 207.3767, 207.2927, 207.1996, 207.1309, 207.0838, 
    207.0437, 207.0053, 206.9721, 206.9445, 206.9378, 206.9191, 206.9141, 
    206.8996,
  207.5264, 207.4238, 207.2986, 207.2065, 207.102, 207.0157, 206.957, 
    206.9102, 206.8651, 206.8244, 206.7888, 206.7667, 206.7506, 206.7432, 
    206.7339,
  207.5609, 207.3996, 207.2568, 207.1687, 207.0726, 206.9815, 206.8932, 
    206.8375, 206.7882, 206.7396, 206.6976, 206.6667, 206.6501, 206.6444, 
    206.6408,
  207.6188, 207.4429, 207.306, 207.215, 207.0717, 206.9666, 206.8828, 
    206.8176, 206.7607, 206.7086, 206.6626, 206.6171, 206.5917, 206.5851, 
    206.5894,
  207.6835, 207.5346, 207.3685, 207.2324, 207.1229, 207.0157, 206.9076, 
    206.8334, 206.7606, 206.7108, 206.6593, 206.6111, 206.574, 206.5611, 
    206.5618,
  207.758, 207.6391, 207.4726, 207.3314, 207.2352, 207.108, 206.9972, 
    206.9013, 206.8101, 206.7589, 206.7, 206.6514, 206.6042, 206.5789, 
    206.5785,
  207.848, 207.7408, 207.6214, 207.4792, 207.3068, 207.2055, 207.1245, 
    207.0158, 206.9236, 206.8378, 206.7702, 206.7212, 206.6769, 206.6512, 
    206.6376,
  207.9824, 207.8371, 207.7034, 207.6029, 207.4794, 207.411, 207.3001, 
    207.1424, 207.0883, 206.9945, 206.907, 206.8595, 206.8207, 206.7973, 
    206.7724,
  208.6486, 208.6031, 208.543, 208.4675, 208.4039, 208.3493, 208.3038, 
    208.2488, 208.1802, 208.0984, 208.0042, 207.9151, 207.8298, 207.7404, 
    207.6467,
  208.5612, 208.5366, 208.5001, 208.4552, 208.4062, 208.3494, 208.2943, 
    208.2416, 208.1773, 208.093, 207.996, 207.8944, 207.8056, 207.7233, 
    207.6452,
  208.5345, 208.5194, 208.4728, 208.4009, 208.3117, 208.2459, 208.206, 
    208.1688, 208.1252, 208.0515, 207.9609, 207.8558, 207.7526, 207.6597, 
    207.5798,
  208.5495, 208.534, 208.4849, 208.4462, 208.3826, 208.3112, 208.226, 
    208.1491, 208.0617, 207.9776, 207.8944, 207.7976, 207.6932, 207.5952, 
    207.5081,
  208.5962, 208.5713, 208.546, 208.5084, 208.4467, 208.369, 208.2656, 
    208.1709, 208.036, 207.8997, 207.7917, 207.7077, 207.6188, 207.5262, 
    207.425,
  208.6342, 208.5425, 208.4355, 208.4014, 208.3529, 208.2912, 208.2399, 
    208.1615, 208.0358, 207.87, 207.7466, 207.6505, 207.5606, 207.4645, 
    207.3543,
  208.547, 208.4579, 208.3656, 208.3774, 208.382, 208.2969, 208.2229, 
    208.1532, 208.0617, 207.9189, 207.7745, 207.641, 207.5288, 207.4136, 
    207.2914,
  208.5497, 208.4977, 208.4263, 208.3474, 208.2718, 208.2003, 208.1594, 
    208.1075, 208.0327, 207.9345, 207.8177, 207.6898, 207.5612, 207.4298, 
    207.2967,
  208.6118, 208.5317, 208.44, 208.3425, 208.2202, 208.1975, 208.1688, 
    208.1038, 208.0096, 207.9093, 207.8272, 207.7335, 207.6251, 207.4919, 
    207.357,
  208.6238, 208.5321, 208.446, 208.3812, 208.2945, 208.2616, 208.2032, 
    208.1117, 208.0427, 207.9349, 207.8497, 207.7859, 207.7128, 207.6132, 
    207.4794,
  207.2157, 207.0726, 206.9534, 206.8367, 206.7454, 206.6622, 206.5863, 
    206.5209, 206.4594, 206.3952, 206.3179, 206.2424, 206.1608, 206.0722, 
    205.974,
  207.3809, 207.2872, 207.1583, 207.0061, 206.9001, 206.8161, 206.7584, 
    206.7051, 206.6499, 206.5884, 206.523, 206.4445, 206.373, 206.2841, 
    206.1903,
  207.5763, 207.4657, 207.3297, 207.1973, 207.0829, 207.0008, 206.9354, 
    206.8755, 206.823, 206.7742, 206.7114, 206.6429, 206.5703, 206.496, 
    206.414,
  207.7598, 207.6412, 207.521, 207.3994, 207.2624, 207.1755, 207.12, 
    207.0619, 206.9989, 206.9418, 206.8851, 206.8354, 206.7749, 206.7074, 
    206.6379,
  207.9374, 207.8301, 207.7212, 207.5872, 207.4736, 207.3847, 207.3079, 
    207.2451, 207.1814, 207.1207, 207.0657, 207.0158, 206.9672, 206.9166, 
    206.8668,
  208.067, 207.9808, 207.8949, 207.7919, 207.6686, 207.5831, 207.5152, 
    207.4475, 207.3746, 207.3041, 207.2455, 207.2089, 207.1772, 207.1455, 
    207.1044,
  208.1818, 208.1051, 208.0184, 207.9124, 207.8205, 207.7567, 207.6858, 
    207.6361, 207.5764, 207.5267, 207.47, 207.4176, 207.3852, 207.3608, 
    207.3429,
  208.2575, 208.1909, 208.107, 208.0306, 207.9762, 207.9167, 207.8518, 
    207.7826, 207.7305, 207.7186, 207.6732, 207.6222, 207.5846, 207.5551, 
    207.5377,
  208.3092, 208.2503, 208.2205, 208.1341, 208.0197, 207.978, 207.9507, 
    207.9125, 207.8592, 207.843, 207.8385, 207.8006, 207.7574, 207.7245, 
    207.6956,
  208.3926, 208.3146, 208.2655, 208.2108, 208.137, 208.1332, 208.0885, 
    208.0283, 208.0029, 207.9655, 207.9609, 207.951, 207.9223, 207.8768, 
    207.8324,
  207.7669, 207.7853, 207.6972, 207.5933, 207.4725, 207.3395, 207.2079, 
    207.0751, 206.956, 206.8402, 206.738, 206.6395, 206.553, 206.4693, 
    206.4061,
  207.7594, 207.7992, 207.7735, 207.715, 207.6004, 207.4706, 207.3405, 
    207.2158, 207.0953, 206.9879, 206.8867, 206.7937, 206.7234, 206.6494, 
    206.5848,
  207.6774, 207.7485, 207.7721, 207.7531, 207.6786, 207.6087, 207.514, 
    207.4004, 207.2669, 207.1386, 207.0233, 206.9139, 206.8308, 206.7508, 
    206.6836,
  207.6162, 207.6561, 207.6985, 207.7097, 207.6647, 207.6271, 207.5611, 
    207.4781, 207.3562, 207.2249, 207.1035, 206.9964, 206.9137, 206.8289, 
    206.748,
  207.688, 207.6721, 207.6712, 207.6617, 207.639, 207.6158, 207.5589, 
    207.497, 207.4004, 207.3012, 207.1967, 207.1101, 207.0207, 206.9406, 
    206.8621,
  207.8772, 207.8073, 207.7537, 207.7257, 207.6806, 207.6383, 207.5873, 
    207.532, 207.459, 207.3768, 207.2944, 207.2095, 207.1267, 207.0436, 
    206.953,
  208.1587, 208.0627, 207.9663, 207.8873, 207.8219, 207.7582, 207.6921, 
    207.6426, 207.5854, 207.525, 207.4567, 207.3744, 207.2758, 207.1836, 
    207.0801,
  208.4238, 208.3404, 208.2191, 208.108, 208.0479, 207.9618, 207.8741, 
    207.8115, 207.7482, 207.6967, 207.6282, 207.5469, 207.4465, 207.3376, 
    207.2275,
  208.7157, 208.6283, 208.5273, 208.4135, 208.2902, 208.191, 208.1137, 
    208.0382, 207.9631, 207.8866, 207.8209, 207.7415, 207.6454, 207.5335, 
    207.4187,
  209.0137, 208.9072, 208.7947, 208.6953, 208.5832, 208.5179, 208.4274, 
    208.31, 208.2364, 208.1362, 208.0456, 207.9736, 207.8784, 207.7845, 
    207.6817,
  207.1093, 207.0723, 207.0499, 207.0336, 207.0173, 207.0004, 206.9956, 
    207.0083, 207.0281, 207.0449, 207.0638, 207.0757, 207.0845, 207.0823, 
    207.0894,
  207.2665, 207.2406, 207.193, 207.17, 207.1579, 207.1302, 207.1241, 
    207.1319, 207.1541, 207.1733, 207.206, 207.2388, 207.2635, 207.2848, 
    207.2924,
  207.4406, 207.4278, 207.3937, 207.3694, 207.3566, 207.338, 207.3356, 
    207.3441, 207.3719, 207.4013, 207.4326, 207.4642, 207.4951, 207.5235, 
    207.5494,
  207.5884, 207.5768, 207.5413, 207.5187, 207.5128, 207.5033, 207.5106, 
    207.5383, 207.5718, 207.603, 207.618, 207.6392, 207.6695, 207.7231, 
    207.7738,
  207.7755, 207.7366, 207.6957, 207.676, 207.6799, 207.6783, 207.6857, 
    207.7189, 207.7619, 207.8025, 207.8215, 207.8426, 207.8748, 207.9291, 
    207.9912,
  208.0072, 207.9537, 207.9088, 207.8921, 207.8675, 207.8473, 207.8449, 
    207.8692, 207.9062, 207.948, 207.9826, 208.0185, 208.0665, 208.1212, 
    208.1821,
  208.3025, 208.2296, 208.1501, 208.0927, 208.066, 208.0431, 208.0223, 
    208.0344, 208.0543, 208.0879, 208.1302, 208.1814, 208.2354, 208.28, 
    208.3155,
  208.6897, 208.5879, 208.4815, 208.3924, 208.3543, 208.3082, 208.2698, 
    208.2617, 208.2528, 208.267, 208.2914, 208.3283, 208.3713, 208.4056, 
    208.4362,
  209.1208, 209.0014, 208.8977, 208.7946, 208.6782, 208.6098, 208.5758, 
    208.5544, 208.5355, 208.52, 208.5154, 208.5313, 208.5694, 208.6005, 
    208.6264,
  209.6369, 209.4927, 209.3405, 209.2254, 209.1071, 209.0357, 208.9826, 
    208.8984, 208.8753, 208.8556, 208.8257, 208.8192, 208.824, 208.8425, 
    208.862,
  208.8835, 208.8253, 208.7606, 208.7052, 208.6567, 208.6102, 208.5767, 
    208.5516, 208.5284, 208.4999, 208.4805, 208.4673, 208.4649, 208.4608, 
    208.4522,
  209.0711, 209.0155, 208.9535, 208.8993, 208.8478, 208.7952, 208.7567, 
    208.7283, 208.7032, 208.6797, 208.6576, 208.6443, 208.6375, 208.6315, 
    208.6202,
  209.3062, 209.2574, 209.1928, 209.1299, 209.0655, 209.0109, 208.96, 
    208.9246, 208.8942, 208.8668, 208.8465, 208.8295, 208.8173, 208.801, 
    208.7783,
  209.5485, 209.4904, 209.4175, 209.3474, 209.2816, 209.2168, 209.1566, 
    209.1124, 209.0784, 209.0449, 209.0198, 208.9983, 208.9804, 208.9555, 
    208.922,
  209.7953, 209.718, 209.6357, 209.5677, 209.5007, 209.4372, 209.3805, 
    209.3336, 209.2931, 209.2573, 209.2181, 209.1862, 209.1456, 209.1138, 
    209.0788,
  210.0335, 209.9511, 209.8715, 209.8118, 209.7265, 209.6488, 209.596, 
    209.555, 209.5219, 209.4793, 209.431, 209.3684, 209.3166, 209.2758, 
    209.2661,
  210.2832, 210.2117, 210.1279, 210.0476, 209.9745, 209.8985, 209.832, 
    209.7879, 209.7491, 209.7063, 209.6572, 209.5933, 209.5336, 209.5021, 
    209.4938,
  210.5578, 210.4987, 210.4171, 210.3223, 210.2528, 210.1642, 210.0884, 
    210.03, 209.9675, 209.9195, 209.8781, 209.8299, 209.7831, 209.7458, 
    209.7229,
  210.8209, 210.7676, 210.7088, 210.6355, 210.5191, 210.4311, 210.3754, 
    210.3165, 210.2494, 210.1747, 210.1264, 210.0824, 210.0405, 209.9908, 
    209.9459,
  211.1152, 211.0668, 210.9872, 210.9209, 210.8282, 210.7745, 210.7253, 
    210.627, 210.5662, 210.4952, 210.4147, 210.373, 210.3275, 210.2775, 
    210.2203,
  211.3463, 211.2988, 211.2202, 211.1429, 211.0598, 210.9868, 210.9241, 
    210.8694, 210.8161, 210.764, 210.7127, 210.6651, 210.6262, 210.5897, 
    210.5555,
  211.5007, 211.4663, 211.3928, 211.3138, 211.2262, 211.1453, 211.0716, 
    211.0066, 210.9451, 210.8867, 210.8244, 210.7667, 210.7135, 210.6639, 
    210.6157,
  211.6781, 211.667, 211.5991, 211.5295, 211.4398, 211.3586, 211.2812, 
    211.2088, 211.1372, 211.0645, 210.9909, 210.9211, 210.8565, 210.7945, 
    210.7363,
  211.829, 211.8252, 211.7711, 211.7122, 211.6324, 211.5503, 211.4759, 
    211.4051, 211.3305, 211.2509, 211.1672, 211.0864, 211.0079, 210.9364, 
    210.8675,
  211.9536, 211.9624, 211.9259, 211.8775, 211.8087, 211.7427, 211.6759, 
    211.6159, 211.5464, 211.4683, 211.38, 211.2898, 211.2031, 211.1229, 
    211.0468,
  212.0384, 212.0623, 212.0443, 212.0215, 211.9576, 211.8948, 211.838, 
    211.7889, 211.7316, 211.6661, 211.5839, 211.4962, 211.4085, 211.326, 
    211.2482,
  212.0621, 212.1059, 212.109, 212.093, 212.049, 212.0123, 211.9659, 
    211.9311, 211.8866, 211.8322, 211.7653, 211.6888, 211.6063, 211.5253, 
    211.4465,
  212.0482, 212.1079, 212.1269, 212.1194, 212.1019, 212.0782, 212.0495, 
    212.0236, 211.9845, 211.9435, 211.892, 211.8294, 211.757, 211.6808, 
    211.6053,
  211.9778, 212.0448, 212.0822, 212.0968, 212.0571, 212.0499, 212.0574, 
    212.0577, 212.0315, 211.9881, 211.9409, 211.8914, 211.832, 211.7686, 
    211.7009,
  211.8991, 211.9577, 211.9826, 212.009, 211.9993, 212.0228, 212.0457, 
    212.0229, 212.0116, 211.975, 211.9227, 211.8823, 211.8313, 211.7833, 
    211.7227,
  211.2546, 211.269, 211.2503, 211.2474, 211.2403, 211.2489, 211.2674, 
    211.2926, 211.3138, 211.3281, 211.3334, 211.3403, 211.3456, 211.3436, 
    211.3372,
  211.1445, 211.1931, 211.1719, 211.1645, 211.151, 211.1595, 211.175, 
    211.2042, 211.2321, 211.2519, 211.2607, 211.2675, 211.273, 211.2731, 
    211.2683,
  211.0512, 211.1145, 211.0912, 211.0885, 211.0672, 211.0649, 211.0764, 
    211.1045, 211.1294, 211.149, 211.1591, 211.1646, 211.1734, 211.1786, 
    211.1789,
  210.9529, 210.9952, 210.9809, 210.9854, 210.9604, 210.9507, 210.9563, 
    210.9824, 211.0083, 211.0264, 211.0368, 211.0406, 211.0474, 211.0589, 
    211.063,
  210.8508, 210.8788, 210.8588, 210.862, 210.847, 210.8461, 210.8434, 
    210.8647, 210.8901, 210.9034, 210.905, 210.9081, 210.9129, 210.9222, 
    210.9358,
  210.7392, 210.755, 210.7431, 210.7502, 210.7045, 210.6921, 210.6981, 
    210.7231, 210.7509, 210.7672, 210.772, 210.7682, 210.7751, 210.7887, 
    210.8123,
  210.6093, 210.6215, 210.6004, 210.5778, 210.5442, 210.5389, 210.5324, 
    210.5628, 210.5902, 210.6167, 210.6231, 210.6292, 210.6356, 210.6574, 
    210.683,
  210.4722, 210.4937, 210.4588, 210.4181, 210.3976, 210.3765, 210.3846, 
    210.4078, 210.4245, 210.4552, 210.4761, 210.493, 210.5078, 210.5358, 
    210.5655,
  210.3327, 210.3389, 210.3166, 210.2811, 210.1923, 210.1949, 210.2378, 
    210.2691, 210.278, 210.2849, 210.3152, 210.3498, 210.3804, 210.4178, 
    210.4468,
  210.2013, 210.1665, 210.1289, 210.1125, 210.0803, 210.1063, 210.1105, 
    210.0964, 210.1375, 210.1463, 210.161, 210.2115, 210.2551, 210.3011, 
    210.3316,
  209.5386, 209.5751, 209.5947, 209.624, 209.6522, 209.6841, 209.714, 
    209.7512, 209.7825, 209.8023, 209.8034, 209.8328, 209.8869, 209.9373, 
    209.9836,
  209.3353, 209.4282, 209.4335, 209.4441, 209.4506, 209.4938, 209.5213, 
    209.5738, 209.6345, 209.6745, 209.6698, 209.6847, 209.7359, 209.7973, 
    209.8501,
  209.1726, 209.2599, 209.2534, 209.2914, 209.3154, 209.3492, 209.3785, 
    209.4403, 209.5005, 209.5425, 209.535, 209.547, 209.6033, 209.678, 
    209.7388,
  208.9937, 209.0634, 209.0823, 209.1597, 209.1842, 209.1997, 209.2342, 
    209.3114, 209.3858, 209.4201, 209.4138, 209.4362, 209.5018, 209.5877, 
    209.6565,
  208.8362, 208.8915, 208.9164, 208.9967, 209.0329, 209.08, 209.1296, 
    209.2092, 209.2801, 209.3039, 209.3041, 209.3456, 209.4225, 209.5133, 
    209.5829,
  208.6802, 208.7327, 208.807, 208.9022, 208.9073, 208.9596, 209.023, 
    209.1078, 209.1721, 209.2039, 209.2298, 209.2754, 209.351, 209.4386, 
    209.5107,
  208.5523, 208.6318, 208.701, 208.7543, 208.7937, 208.8475, 208.9056, 
    208.9999, 209.0689, 209.1297, 209.1755, 209.2249, 209.287, 209.3611, 
    209.4272,
  208.447, 208.5476, 208.5997, 208.6523, 208.7183, 208.7702, 208.8411, 
    208.9174, 208.9642, 209.0594, 209.1264, 209.1968, 209.2464, 209.3023, 
    209.3567,
  208.3563, 208.4724, 208.5591, 208.5879, 208.5817, 208.6802, 208.7984, 
    208.8733, 208.9263, 208.9925, 209.0781, 209.1582, 209.2152, 209.2576, 
    209.2979,
  208.314, 208.3804, 208.4437, 208.5213, 208.5862, 208.7103, 208.7675, 
    208.8057, 208.9, 208.9438, 209.0089, 209.1035, 209.1642, 209.2133, 
    209.2365,
  208.7237, 208.8041, 208.7935, 208.7425, 208.685, 208.6465, 208.6522, 
    208.6851, 208.7087, 208.7241, 208.7327, 208.7132, 208.6895, 208.6719, 
    208.6705,
  208.4886, 208.691, 208.7718, 208.7755, 208.7096, 208.6513, 208.6393, 
    208.6397, 208.6611, 208.6821, 208.6728, 208.6378, 208.5942, 208.581, 
    208.5929,
  208.4915, 208.6458, 208.7001, 208.6998, 208.6385, 208.6057, 208.5874, 
    208.5776, 208.6022, 208.6196, 208.6125, 208.5713, 208.5193, 208.5109, 
    208.5274,
  208.4796, 208.5397, 208.6369, 208.6346, 208.5729, 208.5539, 208.536, 
    208.5509, 208.5616, 208.5766, 208.5757, 208.5323, 208.4804, 208.464, 
    208.4792,
  208.4613, 208.5038, 208.534, 208.5043, 208.4823, 208.4641, 208.4653, 
    208.4957, 208.5117, 208.5267, 208.5059, 208.4606, 208.4124, 208.394, 
    208.42,
  208.427, 208.4453, 208.4832, 208.4376, 208.3734, 208.3751, 208.409, 
    208.4458, 208.4546, 208.4461, 208.414, 208.3749, 208.337, 208.3274, 
    208.3486,
  208.4136, 208.4221, 208.4062, 208.3416, 208.323, 208.3189, 208.3236, 
    208.3545, 208.3704, 208.3559, 208.3111, 208.263, 208.2275, 208.2236, 
    208.2294,
  208.3918, 208.3989, 208.3524, 208.2921, 208.2875, 208.2724, 208.2907, 
    208.2989, 208.2862, 208.2742, 208.2438, 208.2055, 208.1535, 208.1234, 
    208.1049,
  208.3953, 208.3954, 208.3694, 208.2668, 208.2112, 208.2643, 208.2858, 
    208.2771, 208.2409, 208.2064, 208.1915, 208.152, 208.0956, 208.0548, 
    208.0486,
  208.4269, 208.3658, 208.352, 208.2941, 208.2832, 208.3099, 208.2647, 
    208.2499, 208.2433, 208.1624, 208.1353, 208.0955, 208.0556, 208.0347, 
    208.0258,
  208.3918, 208.4903, 208.5357, 208.5624, 208.5461, 208.513, 208.476, 
    208.4418, 208.3971, 208.3461, 208.284, 208.2233, 208.1778, 208.1251, 
    208.071,
  208.2239, 208.3925, 208.4509, 208.4957, 208.5172, 208.5228, 208.5193, 
    208.4884, 208.4475, 208.3993, 208.3403, 208.2819, 208.234, 208.1799, 
    208.1288,
  208.1729, 208.3008, 208.3544, 208.4242, 208.4497, 208.4657, 208.4832, 
    208.4872, 208.4821, 208.4528, 208.3942, 208.3268, 208.2662, 208.2094, 
    208.1577,
  208.0492, 208.1353, 208.2391, 208.3318, 208.3488, 208.3865, 208.423, 
    208.4508, 208.4657, 208.4438, 208.4006, 208.3495, 208.2989, 208.2464, 
    208.1891,
  207.9525, 208.0177, 208.095, 208.1598, 208.2273, 208.2781, 208.3282, 
    208.3761, 208.4088, 208.3945, 208.3649, 208.3294, 208.2909, 208.245, 
    208.1929,
  207.8479, 207.8712, 207.9272, 207.9902, 208.0472, 208.1293, 208.2073, 
    208.2776, 208.324, 208.3259, 208.3031, 208.272, 208.241, 208.2143, 
    208.1797,
  207.7627, 207.7753, 207.7928, 207.8166, 207.8955, 207.9639, 208.0328, 
    208.1075, 208.1592, 208.1843, 208.1691, 208.1437, 208.1236, 208.105, 
    208.0773,
  207.6721, 207.696, 207.6935, 207.7007, 207.7499, 207.7889, 207.8535, 
    207.9053, 207.9487, 207.9922, 207.9955, 207.9877, 207.9693, 207.9525, 
    207.9233,
  207.5958, 207.6203, 207.619, 207.6019, 207.6025, 207.671, 207.7303, 
    207.7544, 207.7773, 207.7976, 207.8306, 207.8295, 207.8143, 207.7893, 
    207.7679,
  207.5409, 207.5276, 207.529, 207.5321, 207.5333, 207.5756, 207.5753, 
    207.5985, 207.639, 207.629, 207.664, 207.678, 207.6811, 207.6618, 207.6404,
  209.3607, 209.4769, 209.5174, 209.4929, 209.4047, 209.3062, 209.1972, 
    209.0722, 208.8915, 208.6881, 208.5014, 208.3378, 208.1855, 208.0424, 
    207.8983,
  209.0816, 209.2405, 209.3271, 209.3726, 209.381, 209.3522, 209.2993, 
    209.2146, 209.1049, 208.9574, 208.7785, 208.5925, 208.4285, 208.2755, 
    208.1415,
  208.7938, 208.9867, 209.0855, 209.1795, 209.2355, 209.2629, 209.2602, 
    209.2206, 209.1619, 209.0645, 208.9394, 208.7973, 208.6586, 208.5335, 
    208.4137,
  208.4781, 208.6427, 208.7625, 208.8849, 208.9594, 209.0316, 209.094, 
    209.1158, 209.1095, 209.0656, 208.9813, 208.8759, 208.7632, 208.6597, 
    208.5513,
  208.1806, 208.3031, 208.4424, 208.5655, 208.6815, 208.7927, 208.8708, 
    208.938, 208.9584, 208.9483, 208.9042, 208.8381, 208.7587, 208.6793, 
    208.5927,
  207.9139, 208.0058, 208.129, 208.2397, 208.3404, 208.4426, 208.5527, 
    208.6573, 208.731, 208.7596, 208.7498, 208.7101, 208.6664, 208.6172, 
    208.5657,
  207.6859, 207.7705, 207.8576, 207.9316, 208.0519, 208.1717, 208.2679, 
    208.3746, 208.4624, 208.519, 208.5357, 208.5193, 208.4997, 208.4901, 
    208.4745,
  207.4892, 207.5754, 207.6398, 207.7049, 207.8301, 207.9177, 208.0029, 
    208.0958, 208.1711, 208.2462, 208.2896, 208.3031, 208.3068, 208.3207, 
    208.3204,
  207.3512, 207.4354, 207.51, 207.5447, 207.5768, 207.6809, 207.807, 
    207.8824, 207.9387, 208.0026, 208.0595, 208.1004, 208.1259, 208.1388, 
    208.1385,
  207.2917, 207.3301, 207.3881, 207.4365, 207.4908, 207.5915, 207.654, 
    207.6883, 207.7643, 207.8052, 207.8707, 207.9329, 207.9738, 207.9921, 
    207.9968,
  208.0551, 207.9024, 207.6305, 207.2708, 206.8784, 206.5204, 206.2018, 
    205.9042, 205.6281, 205.364, 205.1221, 204.9225, 204.7419, 204.5466, 
    204.3253,
  208.2993, 208.1771, 208.0182, 207.775, 207.4754, 207.1196, 206.7773, 
    206.4467, 206.1463, 205.8662, 205.6083, 205.3758, 205.1766, 205.0011, 
    204.8383,
  208.4899, 208.4273, 208.3024, 208.1248, 207.9227, 207.6574, 207.3596, 
    207.0376, 206.7214, 206.4218, 206.1468, 205.8996, 205.6756, 205.4808, 
    205.3094,
  208.4988, 208.5587, 208.5362, 208.3999, 208.2388, 208.0581, 207.8476, 
    207.5976, 207.3185, 207.0326, 206.7485, 206.4818, 206.2456, 206.0293, 
    205.8442,
  208.3496, 208.4465, 208.5361, 208.5365, 208.4549, 208.334, 208.187, 
    208.0222, 207.8193, 207.5715, 207.3192, 207.0674, 206.837, 206.6264, 
    206.4379,
  208.1223, 208.2679, 208.4216, 208.4937, 208.4881, 208.4461, 208.3786, 
    208.3006, 208.1904, 208.0315, 207.8123, 207.5832, 207.3663, 207.1732, 
    206.9942,
  207.8744, 208.0332, 208.1849, 208.3011, 208.3652, 208.3894, 208.3902, 
    208.3799, 208.3502, 208.2861, 208.1818, 208.0257, 207.8408, 207.6502, 
    207.487,
  207.6113, 207.7599, 207.8926, 208.0011, 208.1295, 208.2216, 208.2903, 
    208.3223, 208.3299, 208.3212, 208.2943, 208.2333, 208.1386, 208.0188, 
    207.8927,
  207.3148, 207.4758, 207.6429, 207.7378, 207.7881, 207.9118, 208.0582, 
    208.1452, 208.1866, 208.2052, 208.2169, 208.2114, 208.175, 208.1084, 
    208.0394,
  207.0872, 207.204, 207.3445, 207.4599, 207.5399, 207.6832, 207.8347, 
    207.9034, 207.9806, 208.0107, 208.0325, 208.073, 208.0845, 208.0714, 
    208.0346,
  207.8125, 207.9366, 207.9198, 207.8008, 207.6246, 207.4029, 207.1635, 
    206.916, 206.7057, 206.554, 206.4483, 206.3729, 206.3155, 206.2382, 
    206.1315,
  207.7966, 207.9233, 207.9915, 208.0009, 207.9396, 207.8187, 207.6604, 
    207.4828, 207.267, 207.048, 206.845, 206.6748, 206.5364, 206.4283, 
    206.3285,
  207.775, 207.8988, 208.0156, 208.0696, 208.0896, 208.0723, 208.0039, 
    207.8995, 207.7612, 207.5771, 207.3689, 207.1504, 206.9454, 206.7649, 
    206.6128,
  207.6905, 207.8234, 207.9497, 208.0342, 208.0939, 208.1325, 208.1387, 
    208.1147, 208.0491, 207.9429, 207.7996, 207.6213, 207.4247, 207.2195, 
    207.0255,
  207.636, 207.751, 207.8718, 207.9607, 208.0446, 208.1256, 208.1824, 
    208.2155, 208.2184, 208.1773, 208.0987, 207.9823, 207.8339, 207.6592, 
    207.4744,
  207.627, 207.7177, 207.8316, 207.9159, 207.9925, 208.0648, 208.1352, 
    208.2028, 208.2445, 208.2613, 208.2378, 208.1919, 208.1105, 208.0045, 
    207.865,
  207.6406, 207.7149, 207.8077, 207.8905, 207.9719, 208.0426, 208.1103, 
    208.1711, 208.2245, 208.2666, 208.283, 208.2665, 208.2359, 208.1794, 
    208.1085,
  207.6676, 207.7336, 207.8001, 207.8589, 207.9633, 208.0433, 208.1166, 
    208.1753, 208.216, 208.2661, 208.3081, 208.3185, 208.3047, 208.2786, 
    208.2434,
  207.6765, 207.7316, 207.8013, 207.8503, 207.8849, 207.9755, 208.095, 
    208.1933, 208.2383, 208.2839, 208.3388, 208.377, 208.3799, 208.3649, 
    208.3406,
  207.7136, 207.7419, 207.7886, 207.8367, 207.8783, 207.9708, 208.0799, 
    208.178, 208.2493, 208.2978, 208.3573, 208.4251, 208.4675, 208.47, 
    208.4517,
  207.3704, 207.3935, 207.3914, 207.3617, 207.3156, 207.2577, 207.2101, 
    207.1687, 207.1334, 207.0877, 207.0321, 206.9699, 206.9188, 206.8833, 
    206.8539,
  207.4925, 207.5373, 207.5343, 207.49, 207.4489, 207.4019, 207.3695, 
    207.3416, 207.3112, 207.2743, 207.229, 207.1707, 207.1116, 207.0708, 
    207.0365,
  207.5566, 207.649, 207.6734, 207.6374, 207.5953, 207.5572, 207.5429, 
    207.5313, 207.5241, 207.5027, 207.4645, 207.4122, 207.3535, 207.3021, 
    207.2595,
  207.6294, 207.7098, 207.7365, 207.7115, 207.6889, 207.6656, 207.6608, 
    207.6654, 207.6728, 207.6669, 207.6476, 207.6085, 207.5681, 207.5194, 
    207.4756,
  207.6563, 207.7401, 207.7697, 207.7581, 207.7581, 207.7615, 207.7725, 
    207.7939, 207.8106, 207.8193, 207.8008, 207.7857, 207.759, 207.7347, 
    207.7063,
  207.6877, 207.7621, 207.7924, 207.7938, 207.7906, 207.7946, 207.828, 
    207.8678, 207.9022, 207.9238, 207.9159, 207.903, 207.8916, 207.893, 
    207.8913,
  207.7293, 207.7952, 207.8218, 207.8191, 207.8187, 207.8301, 207.8569, 
    207.8956, 207.9458, 207.9792, 207.9892, 207.9782, 207.9724, 207.9848, 
    208.0075,
  207.8037, 207.8514, 207.8663, 207.8529, 207.8535, 207.8558, 207.8819, 
    207.9152, 207.9497, 207.9891, 208.0149, 208.0158, 208.013, 208.0255, 
    208.0568,
  207.8979, 207.9285, 207.9462, 207.9315, 207.8807, 207.8701, 207.9115, 
    207.9493, 207.9692, 207.9849, 208.0048, 208.0217, 208.0243, 208.0377, 
    208.065,
  208.0405, 208.0503, 208.0453, 208.0212, 207.9906, 207.9862, 207.9954, 
    207.9974, 208.0132, 208.0088, 207.9947, 208.0134, 208.0272, 208.04, 
    208.0539,
  207.4019, 207.375, 207.3037, 207.2255, 207.1466, 207.074, 207.0392, 
    207.0401, 207.056, 207.0664, 207.062, 207.0472, 207.0438, 207.0439, 
    207.0561,
  207.5987, 207.5829, 207.5249, 207.4396, 207.3512, 207.2804, 207.2453, 
    207.2471, 207.2622, 207.2803, 207.2783, 207.2638, 207.2533, 207.2566, 
    207.2655,
  207.8098, 207.8144, 207.7692, 207.6898, 207.5963, 207.5185, 207.4857, 
    207.4807, 207.502, 207.5155, 207.5188, 207.5021, 207.4921, 207.499, 
    207.5108,
  207.9872, 207.996, 207.9672, 207.8958, 207.8191, 207.7495, 207.7142, 
    207.7164, 207.7395, 207.7601, 207.7656, 207.7557, 207.7493, 207.7575, 
    207.7729,
  208.0993, 208.1246, 208.1159, 208.0589, 208.0135, 207.9689, 207.9507, 
    207.9617, 207.9891, 208.0109, 208.0144, 208.0038, 208.0022, 208.0132, 
    208.0352,
  208.1393, 208.1784, 208.1822, 208.1551, 208.1287, 208.1031, 208.108, 
    208.133, 208.1802, 208.2079, 208.2141, 208.203, 208.1998, 208.2192, 
    208.2443,
  208.1423, 208.1978, 208.2116, 208.2019, 208.1899, 208.1862, 208.2043, 
    208.2439, 208.3009, 208.3421, 208.3564, 208.3468, 208.3436, 208.3633, 
    208.3941,
  208.1407, 208.2004, 208.2149, 208.2086, 208.213, 208.2276, 208.2646, 
    208.3158, 208.3637, 208.4122, 208.4403, 208.4436, 208.445, 208.4668, 
    208.4958,
  208.1556, 208.2042, 208.2296, 208.2265, 208.2039, 208.2344, 208.2974, 
    208.3702, 208.4143, 208.4429, 208.4705, 208.4916, 208.5106, 208.5322, 
    208.567,
  208.2019, 208.2284, 208.229, 208.239, 208.2345, 208.2865, 208.3437, 
    208.3995, 208.4499, 208.4694, 208.483, 208.5073, 208.5416, 208.5727, 
    208.6108,
  208.1829, 208.2244, 208.233, 208.2359, 208.2307, 208.2309, 208.233, 
    208.245, 208.2512, 208.2457, 208.237, 208.2245, 208.219, 208.2266, 
    208.2434,
  208.2344, 208.2958, 208.3111, 208.3097, 208.3014, 208.3044, 208.323, 
    208.3382, 208.35, 208.3464, 208.343, 208.3416, 208.3401, 208.3538, 
    208.3714,
  208.2716, 208.3635, 208.3903, 208.4059, 208.405, 208.4186, 208.4481, 
    208.4725, 208.4905, 208.4951, 208.4931, 208.4932, 208.4962, 208.5061, 
    208.5189,
  208.319, 208.3938, 208.4237, 208.4491, 208.4568, 208.4788, 208.5166, 
    208.5606, 208.5901, 208.6055, 208.6006, 208.6014, 208.6045, 208.6135, 
    208.6264,
  208.3782, 208.4359, 208.4601, 208.4798, 208.4935, 208.5308, 208.5739, 
    208.6304, 208.667, 208.6847, 208.6795, 208.6827, 208.6888, 208.705, 
    208.7283,
  208.441, 208.4901, 208.5009, 208.5139, 208.5134, 208.5459, 208.594, 
    208.6584, 208.7058, 208.729, 208.7222, 208.7149, 208.7173, 208.7348, 
    208.7697,
  208.4913, 208.5418, 208.5355, 208.5302, 208.5216, 208.5512, 208.5926, 
    208.6552, 208.71, 208.7425, 208.7465, 208.737, 208.7381, 208.7523, 
    208.7929,
  208.5495, 208.5838, 208.5698, 208.539, 208.528, 208.5424, 208.583, 
    208.6388, 208.6793, 208.7159, 208.7352, 208.734, 208.7344, 208.7475, 
    208.7822,
  208.6039, 208.6159, 208.6035, 208.5627, 208.5103, 208.5135, 208.5636, 
    208.6234, 208.6534, 208.6646, 208.6829, 208.6964, 208.7074, 208.7191, 
    208.7376,
  208.6453, 208.6395, 208.606, 208.5656, 208.5293, 208.55, 208.5825, 
    208.6085, 208.6386, 208.6351, 208.6284, 208.6425, 208.6552, 208.6656, 
    208.678,
  208.9631, 209.0172, 209.032, 209.0685, 209.0755, 209.0737, 209.076, 
    209.0807, 209.0725, 209.0616, 209.0372, 209.0076, 208.9685, 208.9308, 
    208.8976,
  208.8618, 208.969, 208.9855, 209.011, 209.0169, 209.0053, 209.0065, 
    209.0124, 209.0159, 209.0093, 208.994, 208.9631, 208.9267, 208.8883, 
    208.8563,
  208.7409, 208.8797, 208.8927, 208.9312, 208.9234, 208.9277, 208.9383, 
    208.9604, 208.9726, 208.9696, 208.9512, 208.9267, 208.8953, 208.8626, 
    208.832,
  208.665, 208.779, 208.7989, 208.8465, 208.8503, 208.8621, 208.8735, 
    208.891, 208.909, 208.9088, 208.8929, 208.8719, 208.8462, 208.8131, 
    208.7802,
  208.6341, 208.7294, 208.7349, 208.7609, 208.7802, 208.7964, 208.8087, 
    208.8232, 208.8467, 208.8429, 208.82, 208.7932, 208.7669, 208.738, 208.707,
  208.6222, 208.6873, 208.6811, 208.7155, 208.724, 208.7431, 208.772, 
    208.792, 208.8187, 208.8065, 208.7717, 208.7234, 208.688, 208.6495, 
    208.6227,
  208.5983, 208.6581, 208.6596, 208.6844, 208.6833, 208.7042, 208.7233, 
    208.7485, 208.7704, 208.7631, 208.7298, 208.6772, 208.6293, 208.5897, 
    208.5686,
  208.5964, 208.6355, 208.6498, 208.6564, 208.6556, 208.6661, 208.6872, 
    208.714, 208.716, 208.716, 208.6912, 208.652, 208.603, 208.5634, 208.5372,
  208.5917, 208.6266, 208.6534, 208.6524, 208.6299, 208.6343, 208.6554, 
    208.6724, 208.6665, 208.6486, 208.6322, 208.6151, 208.5795, 208.5461, 
    208.514,
  208.6247, 208.6679, 208.6567, 208.6571, 208.6549, 208.6574, 208.6536, 
    208.6346, 208.634, 208.614, 208.5829, 208.5734, 208.5527, 208.5287, 
    208.4928,
  208.6742, 208.6864, 208.6494, 208.6385, 208.6161, 208.6134, 208.6265, 
    208.657, 208.6944, 208.7241, 208.7574, 208.7925, 208.8315, 208.8546, 
    208.855,
  208.5452, 208.6355, 208.573, 208.5327, 208.4863, 208.4743, 208.4839, 
    208.5117, 208.5334, 208.5479, 208.5636, 208.5857, 208.6148, 208.6395, 
    208.6519,
  208.4535, 208.5676, 208.4974, 208.4651, 208.4084, 208.3879, 208.3867, 
    208.4054, 208.4336, 208.4522, 208.4644, 208.4676, 208.4742, 208.483, 
    208.4907,
  208.3733, 208.4508, 208.3995, 208.3685, 208.2982, 208.2586, 208.2547, 
    208.2892, 208.3258, 208.3407, 208.334, 208.3188, 208.3079, 208.3125, 
    208.3274,
  208.3249, 208.3825, 208.3356, 208.2976, 208.2205, 208.1852, 208.1761, 
    208.2013, 208.2244, 208.233, 208.2169, 208.1928, 208.179, 208.1792, 
    208.1886,
  208.2923, 208.3188, 208.2836, 208.2488, 208.1543, 208.0953, 208.0728, 
    208.0932, 208.1235, 208.1417, 208.1265, 208.0906, 208.0568, 208.037, 
    208.0308,
  208.2402, 208.2686, 208.2422, 208.1894, 208.0949, 208.0428, 207.9987, 
    208.0102, 208.0293, 208.0374, 208.0246, 207.9848, 207.9367, 207.9084, 
    207.898,
  208.16, 208.1973, 208.1635, 208.1066, 208.0353, 207.983, 207.9505, 
    207.9464, 207.91, 207.9073, 207.8985, 207.8804, 207.8412, 207.8081, 
    207.7812,
  208.0891, 208.084, 208.0791, 208.0153, 207.88, 207.8416, 207.8571, 
    207.8667, 207.8206, 207.7661, 207.7343, 207.7217, 207.6982, 207.6764, 
    207.6573,
  208.0345, 208.0105, 207.9849, 207.9324, 207.8119, 207.8035, 207.7858, 
    207.7552, 207.7289, 207.6427, 207.571, 207.5478, 207.5465, 207.5583, 
    207.5531,
  207.6696, 207.7024, 207.7799, 207.8735, 207.9154, 207.9544, 207.9924, 
    208.0396, 208.0877, 208.1365, 208.1808, 208.2231, 208.2665, 208.3034, 
    208.3402,
  207.4065, 207.53, 207.5631, 207.6203, 207.6523, 207.6911, 207.7352, 
    207.7915, 207.8513, 207.9041, 207.951, 207.9895, 208.0299, 208.0712, 
    208.114,
  207.2627, 207.3735, 207.389, 207.4393, 207.4539, 207.4863, 207.5333, 
    207.5958, 207.6671, 207.7304, 207.7829, 207.8242, 207.8663, 207.9097, 
    207.9588,
  207.123, 207.2039, 207.235, 207.2849, 207.2835, 207.2929, 207.3229, 
    207.3799, 207.4462, 207.516, 207.5651, 207.6054, 207.641, 207.6906, 
    207.742,
  207.0696, 207.0866, 207.1165, 207.1473, 207.1579, 207.1687, 207.1767, 
    207.2241, 207.2794, 207.3352, 207.3751, 207.4007, 207.4272, 207.4669, 
    207.5173,
  207.0338, 207.0276, 207.0639, 207.089, 207.0567, 207.0409, 207.049, 
    207.0828, 207.1195, 207.157, 207.1846, 207.1983, 207.2098, 207.2403, 
    207.2822,
  207.0038, 206.9984, 207.0151, 207.0057, 206.98, 206.9795, 206.9813, 
    207.0176, 207.0392, 207.0508, 207.062, 207.073, 207.0829, 207.1018, 
    207.1231,
  206.9411, 206.9436, 206.9382, 206.9341, 206.9571, 206.9334, 206.9296, 
    206.9646, 206.9788, 206.9958, 207, 207.0132, 207.0223, 207.0188, 207.0218,
  206.8804, 206.9107, 206.9324, 206.8871, 206.8361, 206.8596, 206.91, 
    206.944, 206.9559, 206.9697, 206.9734, 206.9789, 206.9792, 206.9844, 
    206.9777,
  206.8712, 206.8502, 206.8602, 206.8407, 206.8214, 206.8919, 206.8821, 
    206.8554, 206.9073, 206.9129, 206.9032, 206.9036, 206.91, 206.9367, 
    206.9562,
  206.3681, 206.3753, 206.4313, 206.5191, 206.59, 206.6541, 206.707, 
    206.7669, 206.8274, 206.8884, 206.9545, 207.032, 207.1076, 207.1794, 
    207.2405,
  206.2259, 206.3053, 206.3415, 206.3972, 206.4547, 206.5155, 206.5614, 
    206.6217, 206.6813, 206.737, 206.7957, 206.8566, 206.9182, 206.978, 
    207.0272,
  206.1359, 206.2248, 206.2554, 206.2991, 206.3311, 206.3761, 206.4275, 
    206.4893, 206.5542, 206.6109, 206.6655, 206.7197, 206.7789, 206.8307, 
    206.884,
  206.0875, 206.157, 206.2033, 206.246, 206.2663, 206.3, 206.3516, 206.4193, 
    206.4869, 206.5472, 206.6001, 206.6533, 206.7094, 206.7569, 206.8141,
  206.1079, 206.1541, 206.1768, 206.2138, 206.2543, 206.3017, 206.3486, 
    206.4164, 206.4844, 206.5438, 206.5942, 206.6384, 206.6864, 206.7461, 
    206.8147,
  206.1398, 206.166, 206.2045, 206.2554, 206.2441, 206.2776, 206.3413, 
    206.419, 206.4952, 206.5602, 206.6108, 206.6514, 206.6904, 206.7532, 
    206.8238,
  206.2072, 206.2361, 206.2526, 206.2545, 206.271, 206.2996, 206.3393, 
    206.4121, 206.4844, 206.5455, 206.599, 206.6337, 206.6743, 206.7338, 
    206.8133,
  206.2884, 206.3051, 206.2695, 206.275, 206.3454, 206.3291, 206.3483, 
    206.3872, 206.4245, 206.4944, 206.5327, 206.5807, 206.6231, 206.6789, 
    206.741,
  206.3574, 206.3758, 206.3672, 206.33, 206.277, 206.3119, 206.3734, 
    206.3909, 206.3934, 206.4109, 206.445, 206.4929, 206.5399, 206.5805, 
    206.6245,
  206.4465, 206.401, 206.3857, 206.3715, 206.3608, 206.4166, 206.3947, 
    206.3476, 206.3944, 206.3713, 206.3791, 206.4097, 206.4338, 206.4713, 
    206.4884,
  206.8451, 206.8351, 206.847, 206.8891, 206.9313, 206.9833, 207.0384, 
    207.09, 207.1375, 207.1754, 207.208, 207.24, 207.2702, 207.2984, 207.3314,
  206.7314, 206.747, 206.7378, 206.7545, 206.7773, 206.8129, 206.8623, 
    206.9181, 206.9666, 207.0123, 207.0461, 207.0779, 207.1034, 207.1291, 
    207.1624,
  206.7027, 206.7081, 206.6851, 206.6637, 206.6476, 206.6632, 206.6918, 
    206.7313, 206.7719, 206.8101, 206.8407, 206.8721, 206.8962, 206.9228, 
    206.9509,
  206.6842, 206.6967, 206.6698, 206.6362, 206.6084, 206.5948, 206.5871, 
    206.5993, 206.6184, 206.6413, 206.6646, 206.6897, 206.713, 206.7419, 
    206.7685,
  206.6633, 206.6503, 206.6371, 206.5972, 206.582, 206.5799, 206.5676, 
    206.5682, 206.5657, 206.5655, 206.5604, 206.5705, 206.5857, 206.6108, 
    206.6346,
  206.6429, 206.627, 206.6218, 206.6071, 206.5501, 206.5241, 206.525, 
    206.5271, 206.5291, 206.52, 206.506, 206.4962, 206.4979, 206.5165, 
    206.5393,
  206.5972, 206.5891, 206.5772, 206.5612, 206.5327, 206.4966, 206.471, 
    206.4765, 206.4892, 206.4912, 206.4791, 206.4572, 206.4433, 206.4513, 
    206.4697,
  206.5309, 206.5388, 206.5077, 206.4881, 206.4918, 206.4412, 206.4095, 
    206.398, 206.3889, 206.4169, 206.4257, 206.4133, 206.393, 206.3906, 
    206.4087,
  206.471, 206.4812, 206.4928, 206.4544, 206.3375, 206.3284, 206.3535, 
    206.3627, 206.3403, 206.3305, 206.3608, 206.3699, 206.3664, 206.3586, 
    206.3624,
  206.4819, 206.4357, 206.4169, 206.4023, 206.372, 206.3831, 206.3481, 
    206.2981, 206.3183, 206.2923, 206.2879, 206.3266, 206.3347, 206.3415, 
    206.3413,
  206.9469, 206.9324, 206.9044, 206.8862, 206.8699, 206.8643, 206.8771, 
    206.8958, 206.918, 206.9462, 206.9693, 206.9989, 207.0127, 207.0306, 
    207.0447,
  206.8872, 206.9155, 206.8983, 206.8771, 206.8576, 206.8527, 206.8607, 
    206.8834, 206.908, 206.9358, 206.9573, 206.9782, 206.9895, 206.995, 
    207.0035,
  206.8867, 206.9332, 206.9301, 206.9157, 206.8894, 206.8754, 206.8771, 
    206.8799, 206.8914, 206.9036, 206.9121, 206.925, 206.9372, 206.9508, 
    206.9697,
  206.862, 206.9043, 206.912, 206.9079, 206.8956, 206.8925, 206.8942, 
    206.8992, 206.9042, 206.9081, 206.9019, 206.8961, 206.8908, 206.8895, 
    206.8957,
  206.813, 206.8524, 206.887, 206.8937, 206.8988, 206.9148, 206.9236, 
    206.9411, 206.952, 206.9557, 206.9523, 206.9426, 206.9324, 206.925, 
    206.9273,
  206.759, 206.793, 206.828, 206.8704, 206.8707, 206.8796, 206.91, 206.9386, 
    206.9632, 206.9723, 206.9689, 206.9584, 206.9548, 206.951, 206.9544,
  206.7117, 206.734, 206.7618, 206.7835, 206.8013, 206.8233, 206.8543, 
    206.8978, 206.9417, 206.9736, 206.9901, 206.9948, 206.9989, 207.0107, 
    207.0245,
  206.6564, 206.6767, 206.6918, 206.6918, 206.7251, 206.742, 206.7706, 
    206.8204, 206.8597, 206.908, 206.9402, 206.9627, 206.98, 207.0073, 
    207.0319,
  206.6125, 206.6129, 206.6344, 206.6385, 206.6058, 206.6225, 206.6716, 
    206.7236, 206.7673, 206.7956, 206.8445, 206.8884, 206.9243, 206.9577, 
    206.9926,
  206.6172, 206.5953, 206.5862, 206.5842, 206.5948, 206.6404, 206.6629, 
    206.6502, 206.6931, 206.7041, 206.7217, 206.7651, 206.8038, 206.8446, 
    206.8779,
  207.2068, 207.2636, 207.2686, 207.2567, 207.2205, 207.1866, 207.1625, 
    207.1641, 207.1702, 207.1806, 207.1797, 207.1791, 207.1798, 207.1756, 
    207.1711,
  207.2701, 207.3341, 207.3474, 207.32, 207.2843, 207.2455, 207.2294, 
    207.2208, 207.2346, 207.2394, 207.2314, 207.2204, 207.2066, 207.1942, 
    207.1781,
  207.3333, 207.4291, 207.4511, 207.43, 207.3996, 207.3675, 207.353, 
    207.3471, 207.3481, 207.346, 207.3318, 207.3149, 207.2943, 207.2798, 
    207.263,
  207.3523, 207.4471, 207.4802, 207.4783, 207.4514, 207.4333, 207.4252, 
    207.442, 207.4494, 207.4519, 207.4275, 207.3911, 207.3575, 207.3312, 
    207.3153,
  207.296, 207.385, 207.4395, 207.4547, 207.4572, 207.4713, 207.4933, 207.53, 
    207.566, 207.586, 207.5789, 207.5532, 207.5234, 207.497, 207.4742,
  207.2295, 207.2949, 207.3426, 207.3702, 207.3732, 207.3924, 207.4451, 
    207.5102, 207.5773, 207.6157, 207.6298, 207.622, 207.6086, 207.6038, 
    207.6083,
  207.1659, 207.2138, 207.2489, 207.2613, 207.2697, 207.2979, 207.3443, 
    207.4197, 207.5001, 207.5614, 207.5951, 207.6091, 207.6225, 207.6384, 
    207.6597,
  207.1307, 207.1654, 207.1841, 207.1681, 207.1765, 207.2007, 207.2427, 
    207.3111, 207.3704, 207.4301, 207.4684, 207.4939, 207.5168, 207.5499, 
    207.5926,
  207.1086, 207.1213, 207.1306, 207.1164, 207.0848, 207.0916, 207.1399, 
    207.1991, 207.2478, 207.2763, 207.3159, 207.347, 207.3851, 207.4299, 
    207.4757,
  207.1257, 207.1128, 207.0951, 207.0772, 207.0673, 207.0856, 207.1118, 
    207.1189, 207.1494, 207.1583, 207.1577, 207.1866, 207.2117, 207.2564, 
    207.3014,
  206.7062, 206.708, 206.7132, 206.7438, 206.7811, 206.8165, 206.8445, 
    206.8713, 206.9031, 206.9364, 206.9678, 206.9959, 207.0188, 207.0387, 
    207.047,
  206.7516, 206.7547, 206.7467, 206.7463, 206.7618, 206.7854, 206.8189, 
    206.8497, 206.8916, 206.9326, 206.9767, 207.0131, 207.0459, 207.0738, 
    207.092,
  206.8385, 206.8547, 206.8463, 206.8335, 206.8304, 206.8336, 206.8546, 
    206.8835, 206.9304, 206.9787, 207.0377, 207.0874, 207.1314, 207.1665, 
    207.1902,
  206.9273, 206.9229, 206.907, 206.8867, 206.8765, 206.8688, 206.8733, 
    206.8997, 206.9396, 206.9907, 207.0466, 207.1003, 207.1487, 207.1921, 
    207.2243,
  206.9823, 206.9819, 206.9772, 206.9679, 206.9721, 206.9784, 206.9826, 
    207.011, 207.0462, 207.0865, 207.1215, 207.1584, 207.1988, 207.2395, 
    207.2775,
  207.0394, 207.0387, 207.0367, 207.0468, 207.0417, 207.0501, 207.0691, 
    207.1066, 207.1475, 207.1872, 207.2115, 207.2312, 207.2525, 207.2901, 
    207.3276,
  207.0977, 207.0978, 207.0977, 207.097, 207.108, 207.1229, 207.1426, 
    207.1774, 207.2259, 207.2745, 207.3096, 207.3326, 207.3496, 207.3795, 
    207.4179,
  207.1699, 207.1725, 207.1684, 207.15, 207.1696, 207.1782, 207.1903, 
    207.2228, 207.2426, 207.2939, 207.3365, 207.3724, 207.3973, 207.4268, 
    207.4704,
  207.2389, 207.2375, 207.2429, 207.2349, 207.2117, 207.2083, 207.2355, 
    207.2658, 207.2805, 207.2959, 207.3318, 207.3757, 207.4128, 207.4436, 
    207.4837,
  207.353, 207.3326, 207.3151, 207.3035, 207.2925, 207.306, 207.3149, 
    207.3101, 207.322, 207.3174, 207.3262, 207.3609, 207.3956, 207.4261, 
    207.4564,
  207.5669, 207.5684, 207.5482, 207.5267, 207.5193, 207.4972, 207.4714, 
    207.4378, 207.401, 207.3613, 207.3252, 207.2952, 207.28, 207.2689, 
    207.2551,
  207.6864, 207.7108, 207.6786, 207.6491, 207.625, 207.6026, 207.5824, 
    207.5502, 207.5213, 207.4829, 207.4528, 207.429, 207.4098, 207.3939, 
    207.3754,
  207.8067, 207.8579, 207.8249, 207.807, 207.7808, 207.7636, 207.744, 
    207.7171, 207.6915, 207.6578, 207.6308, 207.6054, 207.5808, 207.5616, 
    207.5358,
  207.939, 207.966, 207.9375, 207.9268, 207.9105, 207.8916, 207.8701, 
    207.843, 207.814, 207.7739, 207.7396, 207.7077, 207.6957, 207.6816, 
    207.6569,
  208.0416, 208.0584, 208.0342, 208.0333, 208.0421, 208.0511, 208.0343, 
    208.0078, 207.9697, 207.921, 207.8776, 207.8443, 207.829, 207.8176, 
    207.7986,
  208.1171, 208.1362, 208.1217, 208.1431, 208.1413, 208.1465, 208.1412, 
    208.1302, 208.1145, 208.0911, 208.0517, 208.006, 207.973, 207.9456, 
    207.9256,
  208.181, 208.2182, 208.2004, 208.2015, 208.2149, 208.2318, 208.2315, 
    208.2398, 208.246, 208.239, 208.2168, 208.1773, 208.1358, 208.0991, 
    208.0747,
  208.2424, 208.2863, 208.2685, 208.2598, 208.2811, 208.298, 208.2989, 
    208.3089, 208.3085, 208.3203, 208.3234, 208.3092, 208.2745, 208.2469, 
    208.2286,
  208.307, 208.3385, 208.346, 208.3455, 208.3159, 208.322, 208.3574, 
    208.3816, 208.3817, 208.3711, 208.3833, 208.3914, 208.3897, 208.3793, 
    208.3647,
  208.3972, 208.4212, 208.4091, 208.4037, 208.3891, 208.4211, 208.4585, 
    208.4477, 208.4515, 208.4374, 208.4249, 208.4495, 208.461, 208.4718, 
    208.4607,
  209.0135, 208.9866, 208.923, 208.8563, 208.7843, 208.7113, 208.6418, 
    208.5798, 208.5143, 208.4538, 208.402, 208.344, 208.2928, 208.2402, 
    208.2008,
  209.1017, 209.1294, 209.0642, 208.994, 208.9029, 208.8273, 208.7647, 
    208.7102, 208.6571, 208.5987, 208.5441, 208.4787, 208.4262, 208.3787, 
    208.3318,
  209.2169, 209.2683, 209.1974, 209.138, 209.044, 208.9588, 208.9001, 
    208.8574, 208.823, 208.7698, 208.7133, 208.6502, 208.6026, 208.5475, 
    208.4955,
  209.3182, 209.3506, 209.2944, 209.2525, 209.1706, 209.0831, 209.0129, 
    208.9702, 208.9414, 208.9021, 208.8525, 208.796, 208.7442, 208.6966, 
    208.6551,
  209.3631, 209.3821, 209.3233, 209.2918, 209.2335, 209.1736, 209.1067, 
    209.0637, 209.0434, 209.0183, 208.9659, 208.9045, 208.8511, 208.8125, 
    208.7959,
  209.368, 209.3867, 209.3335, 209.325, 209.2653, 209.2099, 209.1642, 
    209.1371, 209.1239, 209.0949, 209.0467, 208.9851, 208.9319, 208.8946, 
    208.8931,
  209.3275, 209.3731, 209.3287, 209.3035, 209.2659, 209.241, 209.1996, 
    209.1815, 209.1701, 209.1575, 209.1238, 209.0762, 209.0204, 208.9943, 
    208.9833,
  209.3083, 209.3648, 209.3311, 209.2971, 209.2833, 209.2593, 209.2377, 
    209.2284, 209.2093, 209.2058, 209.1888, 209.1647, 209.1329, 209.1005, 
    209.0798,
  209.3009, 209.3453, 209.3512, 209.341, 209.2695, 209.2401, 209.2672, 
    209.2738, 209.2524, 209.2256, 209.2156, 209.2094, 209.1885, 209.1739, 
    209.1636,
  209.3232, 209.3608, 209.344, 209.3481, 209.301, 209.3107, 209.3365, 
    209.303, 209.293, 209.275, 209.2391, 209.237, 209.2363, 209.2439, 209.2395,
  210.696, 210.7136, 210.7354, 210.76, 210.7437, 210.7192, 210.6954, 
    210.6826, 210.682, 210.6845, 210.6804, 210.6763, 210.6756, 210.6781, 
    210.6669,
  210.6324, 210.6832, 210.6736, 210.6779, 210.6722, 210.6546, 210.6234, 
    210.61, 210.615, 210.63, 210.6303, 210.6248, 210.6157, 210.6083, 210.5974,
  210.615, 210.6849, 210.6733, 210.6915, 210.7031, 210.6744, 210.6288, 
    210.5962, 210.5926, 210.5982, 210.5917, 210.5794, 210.5654, 210.5568, 
    210.5509,
  210.6062, 210.6691, 210.6823, 210.7216, 210.7402, 210.7128, 210.6523, 
    210.6292, 210.6193, 210.623, 210.5943, 210.5726, 210.5522, 210.5461, 
    210.5375,
  210.5961, 210.6618, 210.6667, 210.6763, 210.6925, 210.6904, 210.6381, 
    210.6193, 210.6105, 210.6113, 210.5907, 210.5727, 210.5605, 210.5639, 
    210.561,
  210.5552, 210.6295, 210.6255, 210.6653, 210.696, 210.7222, 210.6906, 
    210.645, 210.6234, 210.6231, 210.6082, 210.5804, 210.5537, 210.5394, 
    210.5376,
  210.4268, 210.5218, 210.5267, 210.5561, 210.6134, 210.6761, 210.652, 
    210.6063, 210.5876, 210.5961, 210.5904, 210.5554, 210.506, 210.473, 
    210.4584,
  210.2695, 210.3485, 210.3493, 210.3638, 210.4072, 210.4618, 210.4617, 
    210.4497, 210.4358, 210.4525, 210.4502, 210.419, 210.3717, 210.3312, 
    210.3149,
  210.0903, 210.1607, 210.1718, 210.191, 210.1609, 210.1913, 210.2096, 
    210.2313, 210.2393, 210.2438, 210.2359, 210.2233, 210.1962, 210.1754, 
    210.161,
  209.968, 210.0326, 210.004, 210.0175, 210.0131, 210.0351, 210.0332, 
    210.0186, 210.039, 210.043, 210.0264, 210.029, 210.0231, 210.0202, 
    210.0098,
  211.5618, 211.5157, 211.5323, 211.5639, 211.5582, 211.5559, 211.5717, 
    211.5806, 211.5678, 211.5359, 211.4835, 211.4281, 211.3593, 211.2857, 
    211.2289,
  211.4277, 211.4216, 211.405, 211.4527, 211.434, 211.4201, 211.4124, 
    211.3999, 211.3931, 211.3462, 211.2967, 211.2577, 211.2031, 211.1298, 
    211.0618,
  211.2957, 211.2629, 211.2358, 211.2922, 211.2753, 211.256, 211.2125, 
    211.2071, 211.2026, 211.1493, 211.0987, 211.0583, 211.0191, 210.9513, 
    210.8691,
  211.1184, 211.1048, 211.1208, 211.1809, 211.1407, 211.0698, 210.9778, 
    210.9899, 210.9915, 210.9486, 210.9003, 210.8539, 210.8259, 210.7807, 
    210.7077,
  210.8784, 210.916, 210.9019, 210.925, 210.9151, 210.8469, 210.7881, 
    210.8046, 210.8021, 210.7653, 210.7033, 210.6524, 210.624, 210.5986, 
    210.5395,
  210.6706, 210.7048, 210.6712, 210.6949, 210.6962, 210.6433, 210.6462, 
    210.6709, 210.6853, 210.6395, 210.5576, 210.4933, 210.4677, 210.4426, 
    210.4011,
  210.5101, 210.5322, 210.4978, 210.5017, 210.4814, 210.4327, 210.4368, 
    210.4782, 210.5136, 210.5058, 210.459, 210.386, 210.3433, 210.2872, 
    210.2628,
  210.3447, 210.3526, 210.3074, 210.3271, 210.3315, 210.2771, 210.2575, 
    210.276, 210.2895, 210.3267, 210.325, 210.2583, 210.1912, 210.1102, 
    210.0786,
  210.135, 210.1506, 210.1627, 210.2414, 210.2242, 210.1933, 210.166, 
    210.1597, 210.1437, 210.1354, 210.14, 210.0889, 210.0278, 209.9504, 
    209.9344,
  209.9638, 209.9699, 209.9524, 210.0624, 210.1475, 210.1385, 210.101, 
    210.0697, 210.0284, 209.9584, 209.9121, 209.8863, 209.8569, 209.8208, 
    209.8401,
  211.9987, 212.102, 212.1747, 212.2271, 212.2352, 212.2492, 212.246, 
    212.2666, 212.3141, 212.3342, 212.3406, 212.3222, 212.2649, 212.216, 
    212.1493,
  211.5833, 211.7122, 211.8039, 211.8722, 211.8983, 211.9412, 211.9286, 
    211.9616, 212.01, 212.0189, 212.0531, 212.0492, 212.0046, 211.9419, 
    211.8692,
  211.1582, 211.3097, 211.4097, 211.4884, 211.5336, 211.5706, 211.5508, 
    211.6124, 211.6707, 211.7105, 211.7401, 211.7031, 211.6771, 211.6404, 
    211.6038,
  210.7191, 210.8539, 210.9524, 211.0616, 211.1372, 211.1882, 211.2235, 
    211.2947, 211.3149, 211.3343, 211.35, 211.3619, 211.3915, 211.3705, 
    211.3333,
  210.2679, 210.3876, 210.4861, 210.6172, 210.7019, 210.8036, 210.8742, 
    210.9478, 210.9815, 210.9921, 210.996, 211.0172, 211.0397, 211.0123, 
    210.9729,
  209.8013, 209.9365, 210.0623, 210.1876, 210.205, 210.2729, 210.3614, 
    210.4592, 210.5275, 210.5211, 210.4929, 210.4918, 210.5432, 210.5974, 
    210.6156,
  209.4106, 209.5276, 209.617, 209.7135, 209.789, 209.8641, 209.9059, 
    209.9888, 210.0618, 210.0726, 210.0751, 210.0717, 210.1182, 210.1975, 
    210.233,
  209.1069, 209.1891, 209.2545, 209.3686, 209.4568, 209.4984, 209.5046, 
    209.5413, 209.5981, 209.6606, 209.7176, 209.7258, 209.7478, 209.8279, 
    209.851,
  208.7351, 208.8219, 208.9545, 209.0237, 209.0097, 209.0996, 209.1747, 
    209.1909, 209.2087, 209.2489, 209.385, 209.4608, 209.4903, 209.5229, 
    209.4869,
  208.418, 208.4763, 208.5703, 208.6863, 208.7536, 208.7953, 208.817, 
    208.8305, 208.8839, 208.9089, 209.044, 209.149, 209.1885, 209.1912, 
    209.1477,
  211.0585, 211.2291, 211.3827, 211.5213, 211.6382, 211.7451, 211.8427, 
    211.9276, 211.9922, 212.0462, 212.0692, 212.0639, 212.0421, 211.9987, 
    211.9462,
  210.5896, 210.7422, 210.8802, 210.9963, 211.1087, 211.2251, 211.349, 
    211.47, 211.5754, 211.6637, 211.7229, 211.7528, 211.7594, 211.7478, 
    211.7243,
  210.1822, 210.3263, 210.4517, 210.568, 210.6678, 210.7784, 210.9005, 
    211.0264, 211.1436, 211.2498, 211.3297, 211.3902, 211.424, 211.4419, 
    211.4463,
  209.7756, 209.8978, 210.0212, 210.1309, 210.2308, 210.3433, 210.4658, 
    210.5978, 210.7222, 210.8229, 210.9072, 210.9806, 211.0445, 211.0975, 
    211.1361,
  209.4032, 209.5152, 209.6301, 209.7216, 209.8347, 209.9656, 210.0867, 
    210.2225, 210.3461, 210.4378, 210.5104, 210.5897, 210.6731, 210.752, 
    210.8143,
  209.0623, 209.1546, 209.2621, 209.3594, 209.4545, 209.574, 209.7128, 
    209.8532, 209.9824, 210.0738, 210.1418, 210.2153, 210.3149, 210.4106, 
    210.4852,
  208.7402, 208.8257, 208.914, 209.0083, 209.1277, 209.2404, 209.3613, 
    209.502, 209.6265, 209.7415, 209.8104, 209.8843, 209.9638, 210.0635, 
    210.1574,
  208.4395, 208.5278, 208.5988, 208.7041, 208.8323, 208.9244, 209.0404, 
    209.1558, 209.2689, 209.3922, 209.4906, 209.5591, 209.6345, 209.7329, 
    209.831,
  208.1518, 208.2493, 208.3514, 208.4448, 208.4849, 208.6146, 208.7631, 
    208.8755, 208.9547, 209.046, 209.172, 209.2645, 209.3364, 209.404, 
    209.4956,
  207.9089, 207.9982, 208.0967, 208.1991, 208.2937, 208.3992, 208.4644, 
    208.5576, 208.6575, 208.715, 208.8234, 208.9615, 209.0465, 209.1001, 
    209.1761,
  210.717, 210.6995, 210.7863, 210.8017, 210.836, 210.8264, 210.8147, 
    210.7748, 210.7199, 210.6461, 210.562, 210.4768, 210.3947, 210.3162, 
    210.2538,
  210.3065, 210.4811, 210.6108, 210.6258, 210.6672, 210.6443, 210.658, 
    210.636, 210.6097, 210.5666, 210.5224, 210.4709, 210.4183, 210.372, 
    210.3379,
  210.011, 210.2372, 210.3415, 210.4061, 210.4619, 210.4559, 210.4979, 
    210.509, 210.5174, 210.4969, 210.4773, 210.4487, 210.4241, 210.3958, 
    210.3785,
  209.7191, 209.8793, 210.081, 210.1734, 210.2334, 210.2475, 210.2871, 
    210.3119, 210.3306, 210.3273, 210.3263, 210.326, 210.3278, 210.3326, 
    210.3374,
  209.476, 209.6026, 209.7905, 209.8916, 209.9647, 210.0002, 210.049, 
    210.0889, 210.1243, 210.1347, 210.1464, 210.1539, 210.1766, 210.1967, 
    210.2132,
  209.2473, 209.3457, 209.4859, 209.6078, 209.6877, 209.7389, 209.8005, 
    209.8345, 209.8717, 209.8833, 209.8932, 209.9121, 209.9393, 209.9731, 
    210.0058,
  209.007, 209.0974, 209.1832, 209.2831, 209.3851, 209.4504, 209.5074, 
    209.551, 209.5859, 209.6062, 209.6244, 209.6465, 209.6758, 209.7096, 
    209.7483,
  208.7695, 208.8528, 208.9118, 209.0016, 209.0911, 209.146, 209.2048, 
    209.2491, 209.2759, 209.3094, 209.3327, 209.3593, 209.3831, 209.4248, 
    209.4567,
  208.4991, 208.5797, 208.6397, 208.7007, 208.7554, 208.8374, 208.9145, 
    208.9536, 208.9765, 209.0028, 209.0381, 209.0685, 209.0978, 209.1239, 
    209.1484,
  208.2621, 208.3068, 208.3684, 208.4458, 208.5045, 208.5696, 208.6101, 
    208.6384, 208.6831, 208.7008, 208.7347, 208.772, 208.8018, 208.819, 
    208.8378,
  209.3749, 209.3293, 209.3063, 209.2877, 209.2706, 209.246, 209.1801, 
    209.079, 208.955, 208.8225, 208.6966, 208.585, 208.4884, 208.3961, 
    208.3097,
  209.3396, 209.2939, 209.2317, 209.1837, 209.1701, 209.1466, 209.1216, 
    209.0585, 208.9727, 208.8624, 208.7543, 208.6451, 208.5472, 208.4596, 
    208.3832,
  209.3007, 209.2814, 209.2229, 209.1538, 209.1134, 209.0744, 209.0482, 
    208.9955, 208.9374, 208.8591, 208.7735, 208.6926, 208.6122, 208.5283, 
    208.4492,
  209.1706, 209.1708, 209.154, 209.11, 209.0492, 208.996, 208.9617, 208.9215, 
    208.8758, 208.8161, 208.7523, 208.6854, 208.6197, 208.5404, 208.4568,
  209.0106, 209.0199, 209.0398, 209.0213, 208.986, 208.9361, 208.8938, 
    208.8463, 208.7963, 208.7351, 208.6757, 208.6148, 208.5571, 208.4877, 
    208.4132,
  208.8131, 208.8285, 208.8787, 208.8986, 208.8625, 208.8186, 208.7886, 
    208.7512, 208.7025, 208.6428, 208.5773, 208.5129, 208.449, 208.3865, 
    208.32,
  208.587, 208.6204, 208.6817, 208.6999, 208.6978, 208.6759, 208.6547, 
    208.6268, 208.5846, 208.5252, 208.4608, 208.389, 208.3265, 208.2687, 
    208.2099,
  208.3703, 208.4178, 208.4585, 208.4861, 208.5195, 208.5002, 208.4779, 
    208.4612, 208.4168, 208.3962, 208.3424, 208.289, 208.2218, 208.1674, 
    208.1154,
  208.161, 208.2332, 208.27, 208.2842, 208.262, 208.2803, 208.3069, 208.2953, 
    208.2625, 208.2381, 208.2104, 208.1749, 208.1282, 208.0784, 208.0343,
  207.9897, 208.0278, 208.0513, 208.0903, 208.0967, 208.1494, 208.1427, 
    208.1015, 208.1067, 208.0739, 208.062, 208.049, 208.0164, 207.9814, 
    207.9374,
  208.3125, 208.3261, 208.3684, 208.3987, 208.443, 208.4733, 208.4655, 
    208.3904, 208.2473, 208.0765, 207.8994, 207.7281, 207.57, 207.4124, 
    207.2754,
  208.3798, 208.4032, 208.4271, 208.4618, 208.4904, 208.5212, 208.5348, 
    208.4955, 208.4083, 208.2679, 208.0982, 207.9179, 207.7424, 207.573, 
    207.4182,
  208.4695, 208.4981, 208.4999, 208.5182, 208.5346, 208.5581, 208.5728, 
    208.5681, 208.5219, 208.4167, 208.2674, 208.0934, 207.9135, 207.739, 
    207.5808,
  208.5569, 208.5704, 208.5634, 208.5703, 208.5852, 208.5937, 208.6046, 
    208.607, 208.579, 208.516, 208.4, 208.2466, 208.0702, 207.8878, 207.713,
  208.6416, 208.6461, 208.6406, 208.625, 208.6309, 208.6274, 208.619, 
    208.6191, 208.5956, 208.5508, 208.4699, 208.349, 208.1945, 208.0234, 
    207.8434,
  208.7045, 208.6951, 208.692, 208.6843, 208.6642, 208.653, 208.6424, 
    208.6226, 208.5981, 208.5567, 208.49, 208.3892, 208.2579, 208.1028, 
    207.9353,
  208.7436, 208.74, 208.73, 208.7065, 208.688, 208.6707, 208.6489, 208.627, 
    208.598, 208.5608, 208.5043, 208.4212, 208.3012, 208.1553, 207.9944,
  208.7313, 208.7423, 208.7348, 208.7195, 208.7183, 208.6902, 208.661, 
    208.6312, 208.5958, 208.5651, 208.5155, 208.4405, 208.3374, 208.2049, 
    208.0512,
  208.6948, 208.7195, 208.7355, 208.7225, 208.6864, 208.668, 208.6581, 
    208.6296, 208.5957, 208.5587, 208.5213, 208.4595, 208.3676, 208.2482, 
    208.1064,
  208.6063, 208.6489, 208.6663, 208.685, 208.6757, 208.676, 208.6403, 
    208.6011, 208.5771, 208.5353, 208.5013, 208.4585, 208.3868, 208.2875, 
    208.1635,
  207.1225, 207.1287, 207.1491, 207.1676, 207.2047, 207.2299, 207.2311, 
    207.1885, 207.1163, 207.0146, 206.8907, 206.7612, 206.6246, 206.491, 
    206.3636,
  207.1692, 207.1813, 207.2003, 207.2202, 207.2613, 207.303, 207.3271, 
    207.3414, 207.3186, 207.2606, 207.1663, 207.0413, 206.9019, 206.7523, 
    206.606,
  207.281, 207.2689, 207.2783, 207.2869, 207.3249, 207.3716, 207.414, 
    207.4395, 207.4539, 207.4479, 207.4003, 207.3214, 207.2023, 207.0544, 
    206.9002,
  207.3905, 207.3913, 207.3979, 207.4027, 207.434, 207.4643, 207.5053, 
    207.5404, 207.5602, 207.5744, 207.5733, 207.532, 207.4668, 207.3513, 
    207.2078,
  207.475, 207.5061, 207.5166, 207.5191, 207.5479, 207.579, 207.6068, 
    207.6466, 207.6716, 207.6952, 207.7133, 207.7074, 207.6733, 207.6124, 
    207.5012,
  207.548, 207.601, 207.6266, 207.6462, 207.6581, 207.6847, 207.7165, 
    207.7444, 207.7724, 207.7939, 207.8255, 207.8457, 207.8472, 207.8227, 
    207.7632,
  207.6294, 207.6859, 207.7205, 207.7484, 207.7641, 207.7889, 207.8114, 
    207.8363, 207.8634, 207.8898, 207.9106, 207.9461, 207.9751, 207.9897, 
    207.9645,
  207.7396, 207.7887, 207.8228, 207.8486, 207.8681, 207.8849, 207.9076, 
    207.9241, 207.935, 207.9604, 207.9772, 208.005, 208.0436, 208.0804, 
    208.1079,
  207.8479, 207.9017, 207.9484, 207.9582, 207.9665, 207.9882, 208.0028, 
    208.0075, 208.0072, 208.0149, 208.0251, 208.0468, 208.0717, 208.107, 
    208.157,
  207.9466, 208.0033, 208.0441, 208.0795, 208.1227, 208.1273, 208.1114, 
    208.1014, 208.1006, 208.0856, 208.0806, 208.0823, 208.0824, 208.1128, 
    208.1462,
  206.7917, 206.7933, 206.7976, 206.7859, 206.7916, 206.8163, 206.8466, 
    206.8766, 206.9023, 206.9167, 206.9195, 206.91, 206.8866, 206.8708, 
    206.8605,
  206.7927, 206.8103, 206.795, 206.7692, 206.772, 206.7936, 206.8315, 
    206.8674, 206.8953, 206.9176, 206.935, 206.9388, 206.9448, 206.9451, 
    206.9499,
  206.8523, 206.8433, 206.8034, 206.7773, 206.7728, 206.7995, 206.8398, 
    206.8814, 206.9181, 206.9428, 206.9635, 206.9816, 207.0045, 207.0247, 
    207.0474,
  206.9312, 206.8965, 206.8531, 206.8124, 206.801, 206.8258, 206.8634, 
    206.9094, 206.9486, 206.9759, 207.0052, 207.0305, 207.0638, 207.0986, 
    207.1394,
  207.0172, 206.9805, 206.9228, 206.8705, 206.863, 206.888, 206.9206, 
    206.9675, 207.0057, 207.0347, 207.064, 207.0968, 207.1346, 207.1722, 
    207.2143,
  207.1056, 207.0635, 206.998, 206.9635, 206.9484, 206.966, 207.0033, 
    207.044, 207.0814, 207.1142, 207.1485, 207.1719, 207.2091, 207.2501, 
    207.3006,
  207.2019, 207.1417, 207.0681, 207.0367, 207.0415, 207.063, 207.0988, 
    207.1356, 207.1723, 207.2128, 207.2397, 207.2687, 207.2989, 207.3373, 
    207.3873,
  207.2856, 207.2084, 207.1542, 207.1313, 207.1279, 207.151, 207.2016, 
    207.2334, 207.2575, 207.2988, 207.3396, 207.3709, 207.4039, 207.439, 
    207.4885,
  207.3503, 207.2798, 207.2453, 207.2068, 207.2151, 207.2653, 207.2854, 
    207.3174, 207.341, 207.3734, 207.425, 207.4708, 207.5109, 207.5446, 
    207.5852,
  207.423, 207.3718, 207.3114, 207.3108, 207.3705, 207.3722, 207.3771, 
    207.4058, 207.4363, 207.4693, 207.5112, 207.5595, 207.604, 207.6404, 
    207.6798,
  207.8504, 207.7839, 207.6936, 207.5966, 207.4974, 207.4118, 207.342, 
    207.2725, 207.1974, 207.1163, 207.0281, 206.9341, 206.8374, 206.7433, 
    206.6551,
  207.9707, 207.9026, 207.8048, 207.6977, 207.5828, 207.4795, 207.3875, 
    207.3016, 207.2086, 207.107, 207.0023, 206.8949, 206.7909, 206.6952, 
    206.6131,
  208.103, 208.0395, 207.9464, 207.8303, 207.7024, 207.5843, 207.4751, 
    207.3676, 207.2593, 207.1397, 207.0221, 206.9096, 206.8062, 206.7128, 
    206.6332,
  208.2246, 208.158, 208.0641, 207.9448, 207.8257, 207.7083, 207.5956, 
    207.4814, 207.3593, 207.2246, 207.0895, 206.9689, 206.8633, 206.7728, 
    206.6967,
  208.335, 208.2739, 208.1802, 208.0655, 207.9529, 207.8402, 207.7259, 
    207.6135, 207.4886, 207.3526, 207.2111, 207.0829, 206.974, 206.8819, 
    206.8044,
  208.4221, 208.3714, 208.2881, 208.1828, 208.0739, 207.9631, 207.8564, 
    207.7492, 207.6303, 207.499, 207.362, 207.2294, 207.118, 207.0249, 
    206.9509,
  208.4892, 208.4379, 208.358, 208.2675, 208.1786, 208.0852, 207.9821, 
    207.8769, 207.7647, 207.6452, 207.5186, 207.3913, 207.2785, 207.1824, 
    207.1074,
  208.5447, 208.4982, 208.4262, 208.3486, 208.267, 208.1797, 208.0893, 
    207.9964, 207.8886, 207.7863, 207.6721, 207.5579, 207.4437, 207.3482, 
    207.2617,
  208.5863, 208.5442, 208.4871, 208.4099, 208.3283, 208.2577, 208.179, 
    208.0992, 207.9995, 207.8998, 207.8018, 207.7037, 207.6015, 207.5038, 
    207.4158,
  208.6185, 208.5779, 208.5124, 208.4542, 208.4008, 208.3326, 208.2494, 
    208.1792, 208.1012, 208.0049, 207.9095, 207.8208, 207.7293, 207.6382, 
    207.5468,
  207.7256, 207.7303, 207.6721, 207.5704, 207.4406, 207.3136, 207.2254, 
    207.1806, 207.171, 207.1768, 207.1828, 207.1659, 207.1241, 207.071, 
    207.0201,
  207.8893, 207.9066, 207.8719, 207.7809, 207.6665, 207.5485, 207.464, 
    207.4066, 207.3803, 207.3613, 207.3457, 207.3163, 207.2821, 207.2461, 
    207.214,
  208.0597, 208.0863, 208.0644, 207.9862, 207.8866, 207.7809, 207.7133, 
    207.6663, 207.6352, 207.606, 207.5675, 207.5211, 207.4733, 207.4342, 
    207.4068,
  208.2525, 208.2542, 208.2213, 208.1384, 208.051, 207.9646, 207.915, 
    207.8847, 207.8586, 207.8249, 207.771, 207.7117, 207.6519, 207.6046, 
    207.5717,
  208.4672, 208.4501, 208.4039, 208.3084, 208.2134, 208.136, 208.0926, 
    208.0747, 208.0553, 208.0156, 207.9537, 207.8865, 207.8235, 207.774, 
    207.7373,
  208.6624, 208.6361, 208.5777, 208.4831, 208.381, 208.2982, 208.2581, 
    208.2442, 208.2296, 208.1935, 208.1339, 208.0668, 208.0084, 207.962, 
    207.9287,
  208.7887, 208.7593, 208.6993, 208.6144, 208.5291, 208.4557, 208.4138, 
    208.3954, 208.3765, 208.3417, 208.2848, 208.218, 208.1622, 208.1233, 
    208.0982,
  208.8196, 208.7916, 208.7568, 208.6918, 208.6173, 208.5592, 208.5324, 
    208.5178, 208.4888, 208.4568, 208.4065, 208.348, 208.2964, 208.2617, 
    208.2394,
  208.7761, 208.7689, 208.7609, 208.705, 208.6394, 208.6247, 208.603, 
    208.5995, 208.57, 208.5376, 208.4968, 208.4486, 208.4054, 208.3688, 
    208.3439,
  208.7267, 208.7265, 208.7043, 208.6579, 208.6592, 208.6546, 208.6278, 
    208.6266, 208.601, 208.5652, 208.5254, 208.4874, 208.4544, 208.4221, 
    208.3967,
  209.336, 209.2871, 209.1868, 209.0721, 208.9437, 208.8224, 208.7195, 
    208.632, 208.5518, 208.4704, 208.3838, 208.2957, 208.2027, 208.1108, 
    208.0227,
  209.4872, 209.4458, 209.3496, 209.2485, 209.1275, 209.0151, 208.9191, 
    208.836, 208.7599, 208.6808, 208.5977, 208.5112, 208.4249, 208.3418, 
    208.2607,
  209.567, 209.5439, 209.4658, 209.3829, 209.2758, 209.1856, 209.1053, 
    209.0361, 208.9666, 208.8928, 208.8123, 208.7286, 208.6456, 208.5652, 
    208.4894,
  209.5956, 209.5812, 209.5199, 209.439, 209.3467, 209.27, 209.204, 209.1516, 
    209.0934, 209.0257, 208.948, 208.8685, 208.7891, 208.7126, 208.637,
  209.5714, 209.5562, 209.5087, 209.4337, 209.3624, 209.3037, 209.2492, 
    209.2101, 209.1658, 209.104, 209.027, 208.9463, 208.8689, 208.7975, 
    208.7271,
  209.4854, 209.4701, 209.4355, 209.382, 209.3257, 209.2818, 209.2422, 
    209.2152, 209.182, 209.1313, 209.0601, 208.9807, 208.9061, 208.8398, 
    208.777,
  209.3551, 209.3432, 209.3119, 209.2684, 209.2311, 209.2095, 209.1883, 
    209.1771, 209.1581, 209.1226, 209.0658, 208.9915, 208.9227, 208.8608, 
    208.8073,
  209.2041, 209.1927, 209.1733, 209.147, 209.1202, 209.1082, 209.1095, 
    209.1149, 209.1023, 209.0819, 209.043, 208.9863, 208.9283, 208.875, 208.83,
  209.0333, 209.0285, 209.0324, 209.0114, 208.9858, 208.9964, 209.008, 
    209.0289, 209.0284, 209.0136, 208.9959, 208.9616, 208.9176, 208.8696, 
    208.8301,
  208.8665, 208.8732, 208.8656, 208.8612, 208.8655, 208.8908, 208.8955, 
    208.9159, 208.925, 208.9165, 208.9064, 208.8928, 208.8673, 208.8344, 
    208.8021,
  210.8037, 210.8282, 210.835, 210.8116, 210.7758, 210.7359, 210.7055, 
    210.6881, 210.6764, 210.6705, 210.6637, 210.6521, 210.6315, 210.6044, 
    210.564,
  210.874, 210.9161, 210.9337, 210.9275, 210.9037, 210.8759, 210.8613, 
    210.8551, 210.861, 210.8585, 210.8511, 210.8335, 210.805, 210.7644, 
    210.7123,
  211.0145, 211.0515, 211.0756, 211.0822, 211.0574, 211.0431, 211.0408, 
    211.0556, 211.0708, 211.0735, 211.0632, 211.0417, 211.0086, 210.9672, 
    210.9191,
  211.0789, 211.1221, 211.1449, 211.1432, 211.1397, 211.1373, 211.1462, 
    211.1689, 211.1877, 211.1918, 211.1808, 211.1518, 211.1192, 211.078, 
    211.0293,
  211.0435, 211.1016, 211.1231, 211.1342, 211.141, 211.1531, 211.1676, 
    211.1942, 211.212, 211.2146, 211.1957, 211.1646, 211.1303, 211.0917, 
    211.0495,
  210.9256, 210.9737, 210.9974, 211.0127, 211.0053, 211.0162, 211.0389, 
    211.0728, 211.0956, 211.1013, 211.0766, 211.0416, 211.0004, 210.9598, 
    210.9129,
  210.6958, 210.7471, 210.7663, 210.7693, 210.7623, 210.7751, 210.7877, 
    210.8124, 210.8283, 210.8275, 210.8034, 210.7642, 210.7185, 210.6766, 
    210.6296,
  210.4159, 210.4627, 210.4695, 210.4661, 210.4464, 210.4418, 210.441, 
    210.4582, 210.4623, 210.4598, 210.4379, 210.4011, 210.3564, 210.3067, 
    210.262,
  210.1163, 210.1516, 210.1589, 210.1509, 210.0974, 210.0905, 210.0921, 
    210.0974, 210.0975, 210.0829, 210.0704, 210.0472, 210.0097, 209.9607, 
    209.9193,
  209.8306, 209.8572, 209.8558, 209.8512, 209.8118, 209.8191, 209.798, 
    209.7864, 209.7955, 209.7761, 209.7523, 209.7325, 209.7036, 209.6632, 
    209.6236,
  210.828, 210.8932, 210.9173, 210.9489, 210.9705, 211.0005, 211.0526, 
    211.1037, 211.1392, 211.1556, 211.159, 211.1546, 211.1463, 211.135, 
    211.1196,
  210.5579, 210.6493, 210.6838, 210.718, 210.7256, 210.7516, 210.7931, 
    210.843, 210.8865, 210.9149, 210.9255, 210.9311, 210.9276, 210.9232, 
    210.9178,
  210.3438, 210.4409, 210.4683, 210.4826, 210.4792, 210.5035, 210.5377, 
    210.5851, 210.6357, 210.6774, 210.7051, 210.7243, 210.7409, 210.7576, 
    210.7728,
  210.1048, 210.1644, 210.1763, 210.1879, 210.177, 210.1952, 210.2223, 
    210.2734, 210.3198, 210.3591, 210.3931, 210.4162, 210.4428, 210.4687, 
    210.499,
  209.8521, 209.8894, 209.8863, 209.8909, 209.8703, 209.8893, 209.9155, 
    209.962, 210.0065, 210.052, 210.0825, 210.1059, 210.1362, 210.1736, 
    210.2168,
  209.6124, 209.6255, 209.6118, 209.6082, 209.5679, 209.5743, 209.5989, 
    209.6429, 209.6893, 209.7318, 209.7599, 209.7874, 209.8186, 209.8666, 
    209.9183,
  209.3676, 209.3702, 209.3411, 209.3141, 209.2861, 209.2936, 209.311, 
    209.3544, 209.4061, 209.4501, 209.48, 209.5031, 209.5318, 209.5747, 
    209.6251,
  209.1749, 209.1595, 209.1118, 209.078, 209.0492, 209.0392, 209.0554, 
    209.098, 209.1372, 209.1759, 209.2072, 209.2307, 209.2573, 209.2992, 
    209.3454,
  209.0189, 208.9725, 208.9213, 208.8872, 208.8206, 208.8219, 208.852, 
    208.877, 208.9115, 208.9345, 208.9616, 208.9895, 209.0157, 209.0516, 
    209.0845,
  208.9194, 208.8537, 208.7784, 208.7379, 208.7032, 208.7085, 208.702, 
    208.7019, 208.7273, 208.7401, 208.7463, 208.7721, 208.7982, 208.8307, 
    208.8545,
  209.3409, 209.3626, 209.3649, 209.3711, 209.3727, 209.3895, 209.4117, 
    209.4336, 209.4559, 209.477, 209.491, 209.5069, 209.5188, 209.5223, 
    209.5215,
  209.1609, 209.2443, 209.2508, 209.2587, 209.2559, 209.269, 209.2944, 
    209.3129, 209.3285, 209.341, 209.3481, 209.3564, 209.3666, 209.375, 
    209.3775,
  209.0156, 209.0959, 209.0963, 209.1118, 209.1082, 209.1264, 209.1479, 
    209.1716, 209.1867, 209.197, 209.2035, 209.207, 209.2119, 209.2215, 
    209.2318,
  208.9362, 208.9845, 208.9813, 208.9797, 208.9697, 208.9802, 208.9986, 
    209.027, 209.0451, 209.0582, 209.0649, 209.066, 209.0683, 209.0772, 
    209.0834,
  208.879, 208.9111, 208.8983, 208.8813, 208.8725, 208.8809, 208.8933, 
    208.9113, 208.9297, 208.938, 208.9436, 208.9459, 208.9455, 208.9477, 
    208.9523,
  208.8519, 208.8697, 208.8517, 208.8387, 208.8163, 208.8131, 208.8199, 
    208.8315, 208.8363, 208.8379, 208.8355, 208.8253, 208.8151, 208.8087, 
    208.8111,
  208.7767, 208.7983, 208.7832, 208.7652, 208.746, 208.7432, 208.7393, 
    208.7407, 208.7391, 208.7271, 208.7123, 208.6905, 208.6763, 208.6651, 
    208.6595,
  208.7157, 208.7392, 208.7249, 208.7045, 208.6889, 208.6754, 208.6717, 
    208.6676, 208.6537, 208.6401, 208.6168, 208.5986, 208.5788, 208.5671, 
    208.5606,
  208.6443, 208.6658, 208.6642, 208.6451, 208.6008, 208.5901, 208.5893, 
    208.5926, 208.578, 208.5495, 208.5291, 208.5174, 208.5077, 208.4993, 
    208.4925,
  208.6135, 208.6184, 208.6023, 208.5877, 208.5669, 208.5613, 208.5452, 
    208.5177, 208.5087, 208.4877, 208.4587, 208.448, 208.4417, 208.4395, 
    208.4329,
  208.3173, 208.2535, 208.2165, 208.2289, 208.245, 208.268, 208.2797, 
    208.2834, 208.2881, 208.3042, 208.3353, 208.3722, 208.4091, 208.441, 
    208.4732,
  208.1658, 208.1697, 208.1226, 208.1213, 208.1244, 208.1424, 208.1562, 
    208.1687, 208.1834, 208.2066, 208.2459, 208.2953, 208.3464, 208.3969, 
    208.4409,
  208.0893, 208.0922, 208.0394, 208.0458, 208.0404, 208.0602, 208.0787, 
    208.1005, 208.1234, 208.1566, 208.2059, 208.2731, 208.3333, 208.3907, 
    208.4361,
  208.0106, 208.0141, 207.9814, 207.989, 207.975, 207.9991, 208.0176, 
    208.0472, 208.0716, 208.1105, 208.163, 208.2347, 208.2993, 208.3588, 
    208.4051,
  207.9609, 207.9477, 207.9159, 207.9151, 207.9229, 207.9496, 207.969, 
    207.9979, 208.0259, 208.0673, 208.1242, 208.1968, 208.2653, 208.3277, 
    208.377,
  207.9618, 207.9298, 207.8892, 207.8985, 207.8927, 207.914, 207.9405, 
    207.9686, 207.9989, 208.0407, 208.098, 208.1587, 208.2308, 208.29, 
    208.3486,
  207.9979, 207.949, 207.8984, 207.885, 207.8834, 207.9011, 207.9154, 
    207.9445, 207.979, 208.0253, 208.0818, 208.1409, 208.2027, 208.2587, 
    208.3162,
  208.0785, 208.0286, 207.9676, 207.9355, 207.9353, 207.9274, 207.9334, 
    207.9548, 207.9786, 208.033, 208.0922, 208.1496, 208.2016, 208.2502, 
    208.299,
  208.1915, 208.1397, 208.0875, 208.036, 207.9892, 207.9694, 207.9859, 
    208.0008, 208.02, 208.0552, 208.1122, 208.17, 208.2137, 208.2538, 208.2924,
  208.3458, 208.2921, 208.2191, 208.1729, 208.1325, 208.1187, 208.0985, 
    208.0763, 208.1011, 208.1134, 208.1433, 208.1933, 208.2272, 208.2565, 
    208.2865,
  208.6668, 208.6266, 208.6033, 208.5978, 208.5884, 208.5873, 208.5757, 
    208.567, 208.5524, 208.5519, 208.5641, 208.5939, 208.6303, 208.6713, 
    208.7106,
  208.4642, 208.4692, 208.4438, 208.4249, 208.4122, 208.4023, 208.3963, 
    208.3953, 208.4009, 208.4104, 208.4254, 208.4492, 208.4811, 208.5137, 
    208.5493,
  208.4265, 208.4148, 208.3783, 208.3595, 208.3375, 208.3152, 208.2991, 
    208.2848, 208.2794, 208.2815, 208.2883, 208.298, 208.3098, 208.3287, 
    208.3466,
  208.418, 208.3934, 208.3565, 208.3386, 208.3002, 208.2606, 208.2225, 
    208.1913, 208.1687, 208.1571, 208.1507, 208.1517, 208.1552, 208.1602, 
    208.1688,
  208.4553, 208.4203, 208.388, 208.3511, 208.3167, 208.2755, 208.2211, 
    208.1692, 208.1246, 208.0868, 208.056, 208.034, 208.0201, 208.0092, 
    208.0011,
  208.5151, 208.4875, 208.4469, 208.4074, 208.3564, 208.2956, 208.2299, 
    208.1663, 208.102, 208.0437, 207.9922, 207.9478, 207.912, 207.8855, 
    207.8659,
  208.5878, 208.563, 208.5114, 208.4526, 208.3972, 208.3315, 208.2453, 
    208.1789, 208.1038, 208.0417, 207.979, 207.9229, 207.8648, 207.8228, 
    207.7902,
  208.6281, 208.6285, 208.5868, 208.5257, 208.4799, 208.4077, 208.3221, 
    208.2483, 208.164, 208.0976, 208.0322, 207.9658, 207.8943, 207.8352, 
    207.7885,
  208.636, 208.6483, 208.6376, 208.5982, 208.5132, 208.4498, 208.4051, 
    208.3465, 208.2774, 208.2052, 208.1369, 208.0694, 207.9924, 207.9168, 
    207.8519,
  208.6462, 208.6425, 208.6319, 208.6166, 208.5709, 208.5462, 208.5001, 
    208.4203, 208.3839, 208.3177, 208.2484, 208.184, 208.1059, 208.0238, 
    207.9445,
  208.2828, 208.3506, 208.4303, 208.5361, 208.6289, 208.7061, 208.7579, 
    208.8004, 208.8323, 208.8518, 208.8635, 208.8698, 208.8699, 208.8696, 
    208.864,
  208.0872, 208.1864, 208.2523, 208.3353, 208.4177, 208.4985, 208.5674, 
    208.6251, 208.6682, 208.7043, 208.7269, 208.7461, 208.7553, 208.7613, 
    208.7616,
  207.9563, 208.0421, 208.0953, 208.1589, 208.2093, 208.2748, 208.3395, 
    208.4023, 208.4594, 208.5081, 208.5446, 208.5726, 208.5969, 208.6149, 
    208.6253,
  207.9118, 207.9761, 207.9977, 208.0229, 208.0517, 208.0918, 208.1318, 
    208.1783, 208.2242, 208.2671, 208.306, 208.3439, 208.3804, 208.4123, 
    208.4307,
  207.9334, 207.9411, 207.9451, 207.9514, 207.9698, 207.9951, 208.0123, 
    208.0347, 208.0563, 208.0786, 208.0961, 208.1188, 208.1467, 208.1783, 
    208.2071,
  207.9908, 207.9962, 207.9916, 207.995, 207.9752, 207.9637, 207.9656, 
    207.9717, 207.978, 207.9775, 207.9724, 207.9603, 207.9594, 207.9706, 
    207.9881,
  208.0954, 208.0832, 208.0569, 208.0309, 208.0223, 208.0045, 207.9797, 
    207.9677, 207.9605, 207.9516, 207.9322, 207.9082, 207.8777, 207.8638, 
    207.8562,
  208.1992, 208.1636, 208.1294, 208.1067, 208.1059, 208.0809, 208.0394, 
    208.0099, 207.9712, 207.9536, 207.9282, 207.8979, 207.854, 207.8167, 
    207.7859,
  208.2745, 208.234, 208.2282, 208.1982, 208.1218, 208.1066, 208.11, 
    208.0789, 208.0325, 207.9816, 207.9502, 207.9179, 207.8766, 207.8315, 
    207.7871,
  208.3342, 208.3068, 208.2793, 208.2566, 208.2227, 208.2283, 208.202, 
    208.1218, 208.0823, 208.0218, 207.9632, 207.929, 207.8879, 207.8435, 
    207.7977,
  208.1151, 208.1532, 208.1611, 208.1568, 208.1395, 208.1102, 208.0667, 
    208.0193, 207.9701, 207.9245, 207.8788, 207.832, 207.7814, 207.7239, 
    207.6604,
  208.1067, 208.1307, 208.1269, 208.1255, 208.1197, 208.0955, 208.0603, 
    208.0223, 207.9839, 207.9512, 207.9222, 207.8934, 207.8577, 207.8175, 
    207.7698,
  208.067, 208.1002, 208.0958, 208.097, 208.0871, 208.0695, 208.0471, 
    208.0202, 207.9929, 207.9664, 207.9469, 207.9288, 207.9139, 207.8913, 
    207.865,
  207.9972, 208.0208, 208.0149, 208.0152, 208.0073, 207.9963, 207.9811, 
    207.9732, 207.968, 207.9606, 207.953, 207.9443, 207.9339, 207.9255, 
    207.9075,
  207.9168, 207.9159, 207.9136, 207.9281, 207.9349, 207.9455, 207.9319, 
    207.9269, 207.9259, 207.9304, 207.9297, 207.9296, 207.9298, 207.9284, 
    207.919,
  207.8556, 207.8494, 207.8472, 207.8732, 207.8752, 207.8811, 207.8819, 
    207.8873, 207.8873, 207.8913, 207.8906, 207.8915, 207.8952, 207.8978, 
    207.8885,
  207.8196, 207.8264, 207.8048, 207.8023, 207.8407, 207.8735, 207.8681, 
    207.8628, 207.8577, 207.8665, 207.8646, 207.8591, 207.8451, 207.8407, 
    207.8309,
  207.8024, 207.7988, 207.768, 207.7565, 207.8072, 207.8556, 207.8469, 
    207.8664, 207.845, 207.8538, 207.8508, 207.8435, 207.814, 207.7821, 
    207.7546,
  207.7945, 207.7547, 207.7691, 207.7545, 207.7211, 207.7957, 207.8296, 
    207.8591, 207.8342, 207.8139, 207.8071, 207.7989, 207.7654, 207.7234, 
    207.6754,
  207.8268, 207.774, 207.7718, 207.7499, 207.7536, 207.8206, 207.8219, 
    207.8297, 207.818, 207.7984, 207.7617, 207.752, 207.719, 207.6756, 
    207.6119,
  208.6704, 208.6699, 208.6831, 208.6995, 208.7217, 208.7454, 208.7714, 
    208.8032, 208.8391, 208.8785, 208.9153, 208.9436, 208.966, 208.976, 
    208.9809,
  208.6139, 208.6279, 208.6461, 208.6483, 208.6611, 208.6676, 208.6776, 
    208.6964, 208.7204, 208.7529, 208.786, 208.8218, 208.8483, 208.8687, 
    208.8808,
  208.5868, 208.6236, 208.6448, 208.6526, 208.6621, 208.6639, 208.6603, 
    208.6611, 208.6646, 208.6786, 208.7002, 208.7293, 208.759, 208.7897, 
    208.8152,
  208.5376, 208.5713, 208.6018, 208.6246, 208.6385, 208.6391, 208.6313, 
    208.6195, 208.6139, 208.6084, 208.617, 208.6292, 208.6558, 208.6874, 
    208.7243,
  208.483, 208.5289, 208.5666, 208.5973, 208.6227, 208.6433, 208.6444, 
    208.6306, 208.6218, 208.609, 208.6028, 208.6023, 208.6183, 208.6436, 
    208.6751,
  208.4342, 208.4812, 208.5281, 208.5764, 208.5921, 208.6093, 208.6253, 
    208.6246, 208.6183, 208.6018, 208.5825, 208.5646, 208.5592, 208.5709, 
    208.5879,
  208.3988, 208.4661, 208.5202, 208.5515, 208.576, 208.5988, 208.6091, 
    208.6225, 208.6272, 208.6211, 208.6032, 208.577, 208.5523, 208.5394, 
    208.5394,
  208.3893, 208.4799, 208.5217, 208.5502, 208.5986, 208.612, 208.6152, 
    208.6138, 208.5986, 208.5895, 208.573, 208.5473, 208.5133, 208.4828, 
    208.4662,
  208.3912, 208.4649, 208.549, 208.5968, 208.6049, 208.6323, 208.6765, 
    208.6822, 208.6561, 208.6102, 208.5822, 208.5567, 208.5223, 208.4809, 
    208.4504,
  208.403, 208.4635, 208.5495, 208.6135, 208.6658, 208.7396, 208.7755, 
    208.7687, 208.7701, 208.7266, 208.6817, 208.6547, 208.6239, 208.5814, 
    208.544,
  208.4617, 208.5202, 208.5966, 208.6799, 208.7625, 208.8332, 208.8941, 
    208.9495, 209, 209.0524, 209.1008, 209.1447, 209.1791, 209.2037, 209.2185,
  208.2965, 208.3725, 208.4436, 208.5031, 208.5815, 208.6551, 208.7258, 
    208.7941, 208.8611, 208.9281, 208.9916, 209.0503, 209.0975, 209.1357, 
    209.1671,
  208.1261, 208.2168, 208.3073, 208.3782, 208.4518, 208.5219, 208.5973, 
    208.6681, 208.7397, 208.8119, 208.8847, 208.9572, 209.0233, 209.0779, 
    209.1257,
  208.0139, 208.0588, 208.1459, 208.2246, 208.3044, 208.3674, 208.4366, 
    208.502, 208.5708, 208.6358, 208.7063, 208.7802, 208.8569, 208.923, 
    208.9812,
  207.9189, 207.9364, 208.0118, 208.0799, 208.1649, 208.239, 208.3056, 
    208.3683, 208.4307, 208.4918, 208.5554, 208.6263, 208.6959, 208.7639, 
    208.8228,
  207.8479, 207.864, 207.9056, 207.9729, 208.0329, 208.0915, 208.1543, 
    208.2133, 208.2673, 208.3203, 208.3704, 208.4322, 208.4975, 208.5695, 
    208.633,
  207.7756, 207.7938, 207.8145, 207.8501, 207.9223, 207.9792, 208.0277, 
    208.0776, 208.1225, 208.1635, 208.2045, 208.2512, 208.3042, 208.3687, 
    208.4333,
  207.7328, 207.7449, 207.7617, 207.771, 207.813, 207.8894, 207.9191, 
    207.9624, 207.9845, 208.0231, 208.054, 208.0906, 208.1257, 208.172, 
    208.2265,
  207.6943, 207.7055, 207.7345, 207.7388, 207.7296, 207.788, 207.8346, 
    207.8797, 207.8924, 207.9104, 207.9377, 207.9664, 207.9903, 208.0186, 
    208.0531,
  207.6804, 207.6866, 207.6979, 207.7115, 207.7153, 207.7577, 207.7955, 
    207.801, 207.8177, 207.8213, 207.8284, 207.8549, 207.8693, 207.8841, 
    207.9008,
  207.9067, 207.9407, 208.0155, 208.0947, 208.1717, 208.2426, 208.309, 
    208.3742, 208.4318, 208.4647, 208.4865, 208.4986, 208.4931, 208.4611, 
    208.4101,
  207.8371, 207.8711, 207.9171, 207.9697, 208.0393, 208.108, 208.1735, 
    208.2371, 208.3018, 208.3546, 208.3922, 208.4176, 208.4327, 208.4346, 
    208.4269,
  207.7826, 207.8122, 207.8403, 207.8882, 207.9455, 208.0007, 208.0684, 
    208.1366, 208.2019, 208.2678, 208.3221, 208.3636, 208.3978, 208.4198, 
    208.4307,
  207.756, 207.7581, 207.7734, 207.8148, 207.8617, 207.9036, 207.95, 
    208.0049, 208.0685, 208.1337, 208.1947, 208.2504, 208.2971, 208.34, 
    208.3719,
  207.7421, 207.7292, 207.7421, 207.7671, 207.8074, 207.8516, 207.8879, 
    207.9228, 207.9724, 208.0283, 208.0852, 208.1452, 208.2008, 208.2586, 
    208.3054,
  207.7567, 207.7337, 207.731, 207.7519, 207.7766, 207.7989, 207.835, 
    207.8653, 207.8967, 207.935, 207.9744, 208.0233, 208.0771, 208.1454, 
    208.207,
  207.7746, 207.7675, 207.7472, 207.7412, 207.7593, 207.7677, 207.7861, 
    207.8145, 207.8485, 207.8872, 207.9203, 207.9522, 207.9881, 208.0432, 
    208.1083,
  207.808, 207.7961, 207.779, 207.7475, 207.7503, 207.762, 207.7699, 
    207.7803, 207.7895, 207.8256, 207.8662, 207.9027, 207.9305, 207.9675, 
    208.0169,
  207.8222, 207.8221, 207.827, 207.7963, 207.7374, 207.737, 207.7636, 
    207.7912, 207.7958, 207.8012, 207.8342, 207.8699, 207.9002, 207.92, 
    207.9494,
  207.8443, 207.8595, 207.8469, 207.8287, 207.7835, 207.7905, 207.8071, 
    207.8073, 207.8125, 207.8127, 207.8173, 207.8496, 207.8769, 207.8963, 
    207.9056,
  208.6782, 208.7276, 208.7878, 208.8471, 208.899, 208.9353, 208.9534, 
    208.958, 208.9573, 208.9544, 208.9519, 208.9482, 208.9444, 208.9457, 
    208.9447,
  208.4612, 208.5354, 208.5905, 208.6285, 208.6661, 208.7011, 208.7283, 
    208.7441, 208.7508, 208.7505, 208.7504, 208.7512, 208.7541, 208.7584, 
    208.7629,
  208.3294, 208.4085, 208.4458, 208.4815, 208.5079, 208.5325, 208.5554, 
    208.5723, 208.5822, 208.5878, 208.5904, 208.5919, 208.5974, 208.6056, 
    208.6153,
  208.2515, 208.2932, 208.3158, 208.349, 208.364, 208.3797, 208.393, 
    208.4084, 208.4196, 208.4231, 208.4239, 208.4256, 208.4339, 208.4452, 
    208.4548,
  208.1828, 208.2164, 208.2323, 208.253, 208.2653, 208.2769, 208.2818, 
    208.2901, 208.2976, 208.3022, 208.3033, 208.3017, 208.3089, 208.3204, 
    208.3332,
  208.1282, 208.1513, 208.1536, 208.1722, 208.173, 208.1761, 208.1765, 
    208.1837, 208.1912, 208.1961, 208.1953, 208.1924, 208.1928, 208.2016, 
    208.2151,
  208.0545, 208.0764, 208.0808, 208.0849, 208.0902, 208.0893, 208.0881, 
    208.1007, 208.1131, 208.1265, 208.1295, 208.1251, 208.1214, 208.1213, 
    208.1306,
  207.9945, 208.0168, 208.0171, 208.006, 208.0062, 208.004, 208.0094, 
    208.0279, 208.0349, 208.0576, 208.0732, 208.0809, 208.0751, 208.0685, 
    208.0676,
  207.9224, 207.9545, 207.9749, 207.9606, 207.9247, 207.9161, 207.9441, 
    207.9793, 207.9938, 208.0039, 208.0222, 208.046, 208.055, 208.0492, 
    208.0413,
  207.87, 207.9048, 207.9068, 207.903, 207.8894, 207.8947, 207.9229, 
    207.9388, 207.96, 207.9679, 207.9672, 207.9951, 208.0115, 208.0146, 
    208.0058,
  207.8558, 207.881, 207.9139, 207.9527, 207.9825, 208.0205, 208.0692, 
    208.1233, 208.1785, 208.2301, 208.2775, 208.319, 208.359, 208.3955, 
    208.4327,
  207.7514, 207.803, 207.8469, 207.8912, 207.9256, 207.9601, 208.0046, 
    208.0596, 208.1213, 208.1779, 208.2314, 208.2766, 208.3247, 208.3709, 
    208.4176,
  207.7077, 207.7653, 207.7968, 207.8302, 207.855, 207.8788, 207.9134, 
    207.9633, 208.0255, 208.0816, 208.1357, 208.1846, 208.2356, 208.288, 
    208.3451,
  207.6897, 207.7285, 207.7471, 207.7683, 207.7741, 207.7873, 207.8094, 
    207.8561, 207.9146, 207.9705, 208.0182, 208.0613, 208.1095, 208.1652, 
    208.2291,
  207.6521, 207.6984, 207.7236, 207.7391, 207.7376, 207.7437, 207.7475, 
    207.7772, 207.8201, 207.8721, 207.9134, 207.9515, 207.9903, 208.0422, 
    208.1045,
  207.6285, 207.672, 207.693, 207.7062, 207.7066, 207.7046, 207.7, 207.7173, 
    207.7512, 207.789, 207.822, 207.844, 207.8667, 207.9044, 207.9616,
  207.5762, 207.625, 207.6492, 207.6584, 207.6669, 207.6703, 207.6701, 
    207.679, 207.6983, 207.7306, 207.752, 207.7631, 207.766, 207.7823, 
    207.8257,
  207.5144, 207.556, 207.578, 207.5815, 207.5939, 207.5979, 207.6029, 
    207.6219, 207.6279, 207.6503, 207.6729, 207.6801, 207.6742, 207.6735, 
    207.7014,
  207.4431, 207.482, 207.5098, 207.5194, 207.4926, 207.5177, 207.5542, 
    207.5922, 207.6093, 207.6234, 207.6512, 207.6729, 207.6883, 207.697, 
    207.7191,
  207.4014, 207.4249, 207.4375, 207.4406, 207.4286, 207.4802, 207.5509, 
    207.5953, 207.6167, 207.6248, 207.6322, 207.6623, 207.6965, 207.7196, 
    207.7424,
  208.2027, 208.2953, 208.3661, 208.4202, 208.4286, 208.4228, 208.4254, 
    208.4585, 208.5154, 208.5841, 208.6445, 208.6807, 208.6943, 208.6938, 
    208.6892,
  208.2071, 208.3192, 208.4065, 208.4564, 208.4678, 208.4711, 208.485, 
    208.5306, 208.6037, 208.6854, 208.7495, 208.7854, 208.7979, 208.7964, 
    208.7911,
  208.2214, 208.3498, 208.4432, 208.4925, 208.503, 208.4964, 208.5079, 
    208.5535, 208.625, 208.7095, 208.7764, 208.8105, 208.822, 208.8224, 
    208.8235,
  208.2427, 208.3436, 208.422, 208.4638, 208.4704, 208.4745, 208.4911, 
    208.5439, 208.6205, 208.7044, 208.7666, 208.7984, 208.811, 208.8166, 
    208.8293,
  208.2627, 208.3415, 208.4132, 208.4427, 208.4456, 208.4553, 208.4764, 
    208.5358, 208.6161, 208.6995, 208.7588, 208.7865, 208.7918, 208.7953, 
    208.8118,
  208.3095, 208.3643, 208.4006, 208.4074, 208.392, 208.388, 208.4158, 
    208.4836, 208.5691, 208.6508, 208.7077, 208.7305, 208.7371, 208.7474, 
    208.7761,
  208.3673, 208.401, 208.4061, 208.3866, 208.358, 208.337, 208.358, 208.417, 
    208.4999, 208.5764, 208.6288, 208.6442, 208.6447, 208.6566, 208.6894,
  208.4326, 208.4414, 208.4312, 208.3944, 208.3454, 208.3143, 208.3184, 
    208.3626, 208.4225, 208.4819, 208.5194, 208.5329, 208.5289, 208.5374, 
    208.5657,
  208.4609, 208.4664, 208.4541, 208.4145, 208.3511, 208.3253, 208.3271, 
    208.3537, 208.3907, 208.4155, 208.4289, 208.4285, 208.4192, 208.4181, 
    208.4286,
  208.4947, 208.4913, 208.4602, 208.4164, 208.3768, 208.3603, 208.3563, 
    208.3605, 208.3688, 208.3663, 208.3548, 208.3426, 208.3348, 208.3316, 
    208.3382,
  208.0653, 208.0984, 208.1032, 208.0936, 208.0725, 208.0621, 208.0772, 
    208.1077, 208.147, 208.1819, 208.2055, 208.2145, 208.2139, 208.2097, 
    208.2117,
  208.1359, 208.1816, 208.1827, 208.1462, 208.1171, 208.0981, 208.1113, 
    208.1476, 208.1933, 208.2342, 208.2622, 208.2791, 208.2864, 208.2908, 
    208.2967,
  208.2057, 208.2863, 208.2954, 208.2639, 208.229, 208.2117, 208.2278, 
    208.263, 208.3045, 208.3366, 208.3532, 208.3606, 208.3624, 208.3675, 
    208.3764,
  208.3048, 208.368, 208.3668, 208.3283, 208.2842, 208.2707, 208.2836, 
    208.3273, 208.3683, 208.3943, 208.4012, 208.4006, 208.398, 208.4035, 
    208.4156,
  208.385, 208.4542, 208.461, 208.4116, 208.3596, 208.3442, 208.3601, 
    208.4021, 208.4486, 208.4744, 208.4753, 208.4664, 208.4621, 208.4718, 
    208.491,
  208.4672, 208.5262, 208.5218, 208.4781, 208.4228, 208.3916, 208.4067, 
    208.445, 208.4855, 208.507, 208.5007, 208.4831, 208.4747, 208.4852, 
    208.5061,
  208.5264, 208.5688, 208.5581, 208.5143, 208.4747, 208.4496, 208.4608, 
    208.4951, 208.5324, 208.5525, 208.5419, 208.5182, 208.503, 208.5126, 
    208.5377,
  208.5585, 208.5882, 208.5797, 208.5448, 208.5042, 208.4831, 208.5053, 
    208.5401, 208.5562, 208.5638, 208.5508, 208.5264, 208.5082, 208.5083, 
    208.5259,
  208.5235, 208.552, 208.5729, 208.5535, 208.5118, 208.5257, 208.5543, 
    208.5935, 208.6124, 208.5974, 208.5817, 208.5636, 208.5506, 208.5454, 
    208.5513,
  208.4743, 208.5093, 208.5148, 208.504, 208.5314, 208.5674, 208.5823, 
    208.613, 208.6373, 208.6317, 208.6074, 208.5975, 208.5958, 208.597, 
    208.5945,
  208.0984, 208.1346, 208.1296, 208.0977, 208.0675, 208.0609, 208.0704, 
    208.088, 208.106, 208.1235, 208.1361, 208.1496, 208.1641, 208.1773, 
    208.1939,
  208.0735, 208.1467, 208.1428, 208.0891, 208.0476, 208.033, 208.0424, 
    208.0613, 208.0755, 208.0829, 208.0826, 208.086, 208.0917, 208.1036, 
    208.1189,
  208.034, 208.1565, 208.1691, 208.1241, 208.0755, 208.0536, 208.0667, 
    208.0914, 208.1078, 208.106, 208.0907, 208.073, 208.0623, 208.0625, 
    208.0716,
  208.0228, 208.127, 208.1428, 208.0988, 208.0474, 208.0294, 208.0504, 
    208.0872, 208.1144, 208.1149, 208.0903, 208.0598, 208.0353, 208.0232, 
    208.022,
  208.0173, 208.114, 208.1381, 208.0892, 208.0355, 208.0208, 208.0451, 
    208.0931, 208.1371, 208.1486, 208.1296, 208.0983, 208.0746, 208.063, 
    208.0616,
  208.0191, 208.0971, 208.1202, 208.0742, 208.0149, 207.9848, 208.0105, 
    208.062, 208.113, 208.1355, 208.1214, 208.0966, 208.0785, 208.079, 
    208.0871,
  207.9946, 208.0691, 208.0849, 208.052, 207.9993, 207.9745, 207.998, 
    208.0481, 208.1043, 208.1349, 208.1282, 208.1052, 208.0947, 208.1043, 
    208.1294,
  207.9588, 208.0443, 208.0532, 208.0246, 207.9765, 207.9467, 207.9839, 
    208.0393, 208.0873, 208.1191, 208.123, 208.1094, 208.1026, 208.1178, 
    208.1492,
  207.9203, 207.9959, 208.0302, 208.0022, 207.9504, 207.9361, 207.9721, 
    208.0347, 208.0849, 208.1061, 208.1196, 208.1251, 208.1293, 208.1509, 
    208.1861,
  207.896, 207.9652, 207.9803, 207.9641, 207.959, 207.9679, 207.9831, 
    208.0348, 208.0819, 208.0993, 208.1045, 208.1189, 208.1393, 208.164, 
    208.1983,
  207.4053, 207.4387, 207.4679, 207.5149, 207.58, 207.6505, 207.7105, 
    207.755, 207.7935, 207.836, 207.8918, 207.9611, 208.0338, 208.1017, 
    208.1589,
  207.3666, 207.4394, 207.4799, 207.4972, 207.551, 207.6125, 207.6762, 
    207.7255, 207.7657, 207.8055, 207.8561, 207.9195, 207.989, 208.0553, 
    208.1114,
  207.3592, 207.4772, 207.5319, 207.5423, 207.5728, 207.6195, 207.6853, 
    207.7434, 207.7949, 207.8402, 207.8941, 207.9562, 208.0222, 208.0824, 
    208.1322,
  207.3576, 207.4713, 207.5263, 207.5338, 207.5538, 207.5938, 207.6597, 
    207.7328, 207.7982, 207.8557, 207.9103, 207.9753, 208.0406, 208.1025, 
    208.1499,
  207.3378, 207.4627, 207.5274, 207.5397, 207.5601, 207.5959, 207.6575, 
    207.7396, 207.8195, 207.8898, 207.9504, 208.0163, 208.0823, 208.1441, 
    208.1964,
  207.3211, 207.4438, 207.5032, 207.5171, 207.5281, 207.5532, 207.6117, 
    207.6943, 207.7804, 207.8583, 207.9222, 207.9804, 208.043, 208.1076, 
    208.168,
  207.2843, 207.4085, 207.4647, 207.4826, 207.4944, 207.5212, 207.5708, 
    207.6492, 207.7379, 207.8171, 207.8801, 207.9307, 207.9832, 208.047, 
    208.1124,
  207.2388, 207.3554, 207.414, 207.4308, 207.4395, 207.4594, 207.5087, 
    207.5858, 207.664, 207.7385, 207.7992, 207.8448, 207.8885, 207.9464, 
    208.0132,
  207.1599, 207.2751, 207.35, 207.3824, 207.3735, 207.3964, 207.453, 
    207.5356, 207.6096, 207.6676, 207.7234, 207.7722, 207.8171, 207.8747, 
    207.9392,
  207.1221, 207.2249, 207.2796, 207.324, 207.3446, 207.3845, 207.4357, 
    207.5054, 207.5818, 207.6318, 207.6739, 207.7227, 207.7711, 207.827, 
    207.8897,
  207.6242, 207.6384, 207.6256, 207.6221, 207.6497, 207.704, 207.7623, 
    207.8317, 207.8889, 207.9329, 207.9673, 208.0106, 208.0797, 208.1652, 
    208.2478,
  207.6192, 207.6602, 207.6601, 207.6208, 207.6052, 207.6374, 207.7027, 
    207.7795, 207.8501, 207.8908, 207.925, 207.9653, 208.0231, 208.1014, 
    208.1759,
  207.5914, 207.715, 207.7491, 207.7205, 207.6874, 207.687, 207.7312, 
    207.7984, 207.8602, 207.8969, 207.9143, 207.9389, 207.9788, 208.0419, 
    208.1102,
  207.5743, 207.6934, 207.7298, 207.7104, 207.6727, 207.6658, 207.7053, 
    207.7688, 207.8375, 207.8828, 207.9094, 207.9249, 207.9549, 208.0002, 
    208.0637,
  207.4855, 207.6245, 207.6888, 207.7032, 207.6834, 207.6836, 207.7233, 
    207.784, 207.8557, 207.908, 207.9377, 207.9547, 207.9772, 208.0156, 
    208.0746,
  207.3928, 207.5282, 207.6024, 207.6288, 207.6171, 207.6151, 207.6587, 
    207.7303, 207.8089, 207.8766, 207.9152, 207.9349, 207.9554, 207.9875, 
    208.0484,
  207.305, 207.4387, 207.5219, 207.5565, 207.5554, 207.5626, 207.6034, 
    207.6767, 207.7645, 207.8457, 207.8949, 207.9239, 207.9488, 207.9853, 
    208.0464,
  207.2736, 207.3946, 207.4702, 207.4968, 207.4958, 207.4942, 207.5247, 
    207.5942, 207.6747, 207.7543, 207.8137, 207.8473, 207.8768, 207.9165, 
    207.9782,
  207.2521, 207.3696, 207.4603, 207.4983, 207.4676, 207.4488, 207.4896, 
    207.5662, 207.6441, 207.7001, 207.7472, 207.7835, 207.8145, 207.8546, 
    207.9068,
  207.2608, 207.3596, 207.4359, 207.4841, 207.4753, 207.4688, 207.4976, 
    207.5412, 207.6136, 207.6635, 207.6803, 207.7078, 207.7354, 207.7696, 
    207.8095,
  208.1269, 208.1611, 208.1422, 208.138, 208.1092, 208.0733, 208.043, 
    208.0416, 208.0692, 208.1035, 208.1234, 208.1153, 208.0917, 208.0754, 
    208.0695,
  208.0094, 208.1347, 208.1624, 208.1369, 208.0764, 208.0222, 207.989, 
    207.9986, 208.0452, 208.1021, 208.1451, 208.1579, 208.1408, 208.122, 
    208.1091,
  207.8732, 208.0384, 208.118, 208.1356, 208.0711, 208.0045, 207.969, 
    207.9818, 208.0384, 208.1083, 208.1713, 208.2034, 208.2113, 208.2106, 
    208.216,
  207.7798, 207.9106, 207.9924, 208.0376, 207.9705, 207.8979, 207.8545, 
    207.8665, 207.9278, 208.0105, 208.086, 208.1303, 208.1527, 208.1674, 
    208.1926,
  207.6784, 207.8113, 207.894, 207.9543, 207.9004, 207.8378, 207.7937, 
    207.8086, 207.8704, 207.9599, 208.0355, 208.0796, 208.0984, 208.1162, 
    208.1462,
  207.6371, 207.7423, 207.8029, 207.8541, 207.8033, 207.7375, 207.6932, 
    207.7137, 207.7808, 207.8726, 207.9437, 207.9784, 207.9885, 208, 208.0324,
  207.5939, 207.6953, 207.7427, 207.7788, 207.7249, 207.6656, 207.6199, 
    207.6407, 207.7112, 207.8018, 207.8683, 207.8892, 207.8864, 207.8857, 
    207.9103,
  207.5644, 207.6515, 207.6898, 207.706, 207.6497, 207.5889, 207.5538, 
    207.5751, 207.6332, 207.71, 207.7597, 207.7687, 207.7536, 207.7465, 
    207.761,
  207.5335, 207.6091, 207.6473, 207.6606, 207.5838, 207.5182, 207.4984, 
    207.5339, 207.5908, 207.6423, 207.6707, 207.668, 207.6478, 207.6395, 
    207.6487,
  207.5239, 207.5829, 207.6006, 207.6103, 207.548, 207.4971, 207.472, 
    207.4939, 207.5425, 207.5834, 207.5834, 207.5671, 207.5439, 207.5376, 
    207.5482,
  207.9353, 207.9177, 207.8877, 207.8904, 207.8886, 207.881, 207.8785, 
    207.8992, 207.9369, 207.9876, 208.0308, 208.0658, 208.082, 208.0787, 
    208.0615,
  207.8991, 207.972, 207.9465, 207.8906, 207.8411, 207.7781, 207.7481, 
    207.7592, 207.7971, 207.8507, 207.9007, 207.9388, 207.96, 207.9613, 
    207.9531,
  207.8683, 208.0014, 208.037, 207.9997, 207.9268, 207.8296, 207.7638, 
    207.7507, 207.7712, 207.8178, 207.8654, 207.9048, 207.931, 207.9376, 
    207.9346,
  207.8729, 207.9721, 208.0062, 207.9904, 207.9231, 207.8254, 207.7528, 
    207.7258, 207.7335, 207.7657, 207.7952, 207.8127, 207.821, 207.821, 
    207.8187,
  207.8418, 207.9385, 207.9783, 207.9746, 207.9232, 207.8529, 207.7865, 
    207.7567, 207.7622, 207.7925, 207.8058, 207.7955, 207.7731, 207.7516, 
    207.7417,
  207.8176, 207.901, 207.9361, 207.9477, 207.9052, 207.8486, 207.7931, 
    207.7698, 207.7823, 207.8111, 207.8108, 207.7756, 207.7346, 207.7036, 
    207.6918,
  207.7847, 207.8634, 207.8897, 207.9142, 207.8936, 207.8541, 207.7982, 
    207.7762, 207.7939, 207.8199, 207.819, 207.7731, 207.7208, 207.6864, 
    207.6776,
  207.7628, 207.8321, 207.8461, 207.8635, 207.8538, 207.8215, 207.7791, 
    207.7659, 207.7752, 207.7946, 207.7922, 207.7507, 207.698, 207.6646, 
    207.6543,
  207.7065, 207.7697, 207.7958, 207.8107, 207.7816, 207.75, 207.7202, 
    207.7227, 207.7278, 207.7303, 207.7348, 207.7224, 207.6948, 207.6721, 
    207.6681,
  207.6413, 207.6874, 207.6901, 207.7087, 207.6895, 207.6724, 207.6444, 
    207.6354, 207.6473, 207.6487, 207.6456, 207.6452, 207.6422, 207.6396, 
    207.6531,
  208.6039, 208.5604, 208.5425, 208.5715, 208.5655, 208.5172, 208.4537, 
    208.392, 208.3594, 208.3591, 208.3752, 208.3984, 208.4117, 208.4099, 
    208.393,
  208.6419, 208.6648, 208.6464, 208.6206, 208.559, 208.4803, 208.3965, 
    208.327, 208.2855, 208.2769, 208.2832, 208.2954, 208.2953, 208.2816, 
    208.2586,
  208.6357, 208.7596, 208.8107, 208.8157, 208.731, 208.6117, 208.487, 
    208.3962, 208.3508, 208.3405, 208.3444, 208.3418, 208.3193, 208.2843, 
    208.2436,
  208.6057, 208.7383, 208.8326, 208.8789, 208.8083, 208.6786, 208.5291, 
    208.4201, 208.3729, 208.3597, 208.363, 208.3518, 208.3153, 208.2585, 
    208.2038,
  208.4964, 208.6673, 208.8099, 208.8903, 208.843, 208.729, 208.5914, 
    208.4944, 208.4618, 208.4594, 208.4672, 208.4477, 208.3948, 208.3236, 
    208.256,
  208.3864, 208.5658, 208.7121, 208.8093, 208.761, 208.6511, 208.5379, 
    208.4713, 208.4637, 208.483, 208.493, 208.4655, 208.3918, 208.3005, 
    208.2234,
  208.2237, 208.4169, 208.5522, 208.6479, 208.6198, 208.5351, 208.4411, 
    208.4036, 208.4229, 208.4662, 208.4926, 208.4676, 208.3851, 208.2863, 
    208.2098,
  208.0849, 208.2673, 208.3789, 208.4379, 208.4114, 208.3458, 208.2764, 
    208.2643, 208.2942, 208.3597, 208.3951, 208.3697, 208.2841, 208.194, 
    208.1348,
  207.9094, 208.0671, 208.1762, 208.2211, 208.1532, 208.0913, 208.0649, 
    208.1024, 208.1618, 208.2237, 208.2603, 208.2404, 208.1776, 208.105, 
    208.067,
  207.749, 207.8691, 207.9501, 207.9854, 207.9375, 207.9072, 207.9025, 
    207.9306, 208.0045, 208.0662, 208.0715, 208.0544, 208.019, 207.984, 
    207.9742,
  207.1084, 207.1922, 207.2856, 207.3833, 207.4298, 207.4286, 207.4243, 
    207.435, 207.482, 207.5638, 207.6567, 207.7447, 207.8215, 207.8874, 
    207.9538,
  207.0738, 207.1867, 207.2928, 207.3656, 207.3925, 207.3856, 207.378, 
    207.404, 207.4758, 207.5757, 207.6876, 207.7868, 207.8621, 207.9237, 
    207.9838,
  207.0885, 207.2856, 207.4429, 207.5427, 207.5435, 207.4998, 207.4653, 
    207.4786, 207.5533, 207.6645, 207.7844, 207.8859, 207.9594, 208.0172, 
    208.0702,
  207.1546, 207.3197, 207.4754, 207.5958, 207.5844, 207.5099, 207.4438, 
    207.4428, 207.5235, 207.6435, 207.7736, 207.8839, 207.9626, 208.0219, 
    208.0754,
  207.2341, 207.3893, 207.5529, 207.6803, 207.6807, 207.6047, 207.5345, 
    207.5314, 207.6185, 207.7484, 207.8815, 207.9846, 208.0542, 208.1039, 
    208.1485,
  207.2816, 207.4403, 207.5903, 207.7037, 207.6821, 207.6017, 207.5317, 
    207.549, 207.648, 207.7893, 207.9202, 208.0062, 208.0501, 208.0768, 
    208.1099,
  207.2536, 207.4296, 207.5965, 207.7076, 207.7036, 207.6309, 207.5618, 
    207.5858, 207.6952, 207.8424, 207.9678, 208.0321, 208.046, 208.0471, 
    208.0656,
  207.1967, 207.3694, 207.5385, 207.6315, 207.6533, 207.605, 207.557, 
    207.5912, 207.6864, 207.8139, 207.9127, 207.9478, 207.9303, 207.9109, 
    207.9232,
  207.1348, 207.2856, 207.4384, 207.5245, 207.5168, 207.4804, 207.4795, 
    207.559, 207.6781, 207.7933, 207.8668, 207.8745, 207.8392, 207.7989, 
    207.8069,
  207.1174, 207.2342, 207.3239, 207.3717, 207.348, 207.3254, 207.3544, 
    207.4372, 207.5815, 207.6992, 207.7542, 207.7597, 207.7257, 207.7008, 
    207.7155,
  207.586, 207.6467, 207.676, 207.7377, 207.8056, 207.8739, 207.9362, 
    207.982, 208.018, 208.0493, 208.0698, 208.0814, 208.0792, 208.0812, 
    208.0779,
  207.4034, 207.5209, 207.5624, 207.558, 207.556, 207.5726, 207.6173, 
    207.6773, 207.7416, 207.8093, 207.8646, 207.9027, 207.9219, 207.9339, 
    207.9384,
  207.2784, 207.4561, 207.5616, 207.5897, 207.5762, 207.5593, 207.568, 
    207.6092, 207.6687, 207.7331, 207.7924, 207.8267, 207.8407, 207.8366, 
    207.8356,
  207.2712, 207.3933, 207.4904, 207.5462, 207.5208, 207.4647, 207.4303, 
    207.448, 207.4985, 207.5547, 207.6069, 207.6348, 207.6479, 207.6561, 
    207.673,
  207.2609, 207.405, 207.5334, 207.6176, 207.608, 207.5489, 207.4895, 
    207.4806, 207.517, 207.5576, 207.5908, 207.6029, 207.6043, 207.6138, 
    207.6354,
  207.3224, 207.4405, 207.5377, 207.6121, 207.5962, 207.5453, 207.4907, 
    207.4826, 207.5178, 207.5575, 207.5784, 207.5744, 207.5635, 207.5642, 
    207.5839,
  207.353, 207.4742, 207.5751, 207.6575, 207.6616, 207.6047, 207.5305, 
    207.504, 207.5378, 207.5992, 207.6515, 207.67, 207.6644, 207.6546, 
    207.6593,
  207.3453, 207.4586, 207.5722, 207.6465, 207.6825, 207.6736, 207.6273, 
    207.6096, 207.6227, 207.6687, 207.7175, 207.7386, 207.7284, 207.7103, 
    207.7136,
  207.3778, 207.4624, 207.5514, 207.6204, 207.6062, 207.6441, 207.6792, 
    207.7474, 207.8119, 207.8569, 207.8937, 207.9011, 207.8772, 207.8456, 
    207.8383,
  207.478, 207.5144, 207.5467, 207.6008, 207.5916, 207.625, 207.7077, 
    207.8212, 207.9398, 208.0125, 208.0295, 208.0315, 208.0126, 207.9943, 
    207.9933,
  209.5917, 209.5951, 209.5372, 209.5031, 209.4684, 209.4302, 209.4014, 
    209.3673, 209.3127, 209.2178, 209.0832, 208.9117, 208.7379, 208.5686, 
    208.4095,
  209.4265, 209.5455, 209.5075, 209.4069, 209.3013, 209.215, 209.1638, 
    209.1379, 209.1181, 209.0717, 208.992, 208.8685, 208.7231, 208.5789, 
    208.4461,
  209.4159, 209.6035, 209.6348, 209.5495, 209.3813, 209.2011, 209.0713, 
    208.9966, 208.9554, 208.9139, 208.8513, 208.7569, 208.6551, 208.5587, 
    208.4821,
  209.5896, 209.6648, 209.6863, 209.6063, 209.4109, 209.1834, 208.9893, 
    208.8756, 208.8108, 208.7642, 208.6901, 208.594, 208.5029, 208.4334, 
    208.3956,
  209.6739, 209.7449, 209.7708, 209.7339, 209.587, 209.3817, 209.1643, 
    209.0118, 208.934, 208.8763, 208.7916, 208.6704, 208.5338, 208.4155, 
    208.3333,
  209.7155, 209.7946, 209.8077, 209.7863, 209.644, 209.4498, 209.2262, 
    209.0641, 208.9799, 208.9212, 208.832, 208.6972, 208.5476, 208.423, 
    208.3436,
  209.6547, 209.7364, 209.7467, 209.7511, 209.6602, 209.5127, 209.3273, 
    209.1771, 209.1004, 209.0593, 208.9925, 208.8631, 208.6991, 208.554, 
    208.4656,
  209.5757, 209.6491, 209.6704, 209.6613, 209.58, 209.4526, 209.3059, 
    209.2066, 209.1381, 209.1109, 209.0687, 208.9693, 208.8224, 208.6748, 
    208.5726,
  209.5185, 209.5741, 209.5974, 209.5849, 209.4423, 209.3092, 209.2067, 
    209.1679, 209.1554, 209.145, 209.1205, 209.0551, 208.9481, 208.8268, 
    208.7278,
  209.5033, 209.5237, 209.5081, 209.4771, 209.3697, 209.2373, 209.1613, 
    209.1544, 209.1926, 209.197, 209.1507, 209.0943, 209.0098, 208.9119, 
    208.8269,
  208.7589, 208.8332, 208.8785, 208.9366, 208.9939, 209.0439, 209.0583, 
    209.0087, 208.8957, 208.7438, 208.6125, 208.5108, 208.4389, 208.3903, 
    208.345,
  208.7206, 208.9591, 209.0105, 208.9805, 208.9749, 208.9774, 208.9742, 
    208.9313, 208.8481, 208.7394, 208.6407, 208.5692, 208.5296, 208.4951, 
    208.4549,
  208.8856, 209.1851, 209.3254, 209.3197, 209.2468, 209.1569, 209.1022, 
    209.0476, 208.97, 208.8671, 208.7615, 208.6821, 208.641, 208.6111, 
    208.5661,
  209.1854, 209.4218, 209.5783, 209.6229, 209.6039, 209.4715, 209.3445, 
    209.2373, 209.1406, 209.0224, 208.9009, 208.7934, 208.7141, 208.649, 
    208.5834,
  209.5209, 209.6863, 209.8106, 209.8984, 209.918, 209.8441, 209.7076, 
    209.5728, 209.4829, 209.382, 209.2488, 209.0978, 208.9644, 208.8492, 
    208.7435,
  209.8441, 209.999, 210.0965, 210.235, 210.2756, 210.206, 210.0609, 
    209.9066, 209.8114, 209.7193, 209.5796, 209.3978, 209.2229, 209.0755, 
    208.938,
  210.034, 210.2432, 210.3589, 210.4811, 210.6122, 210.6111, 210.4993, 
    210.3625, 210.2574, 210.1631, 210.0327, 209.8375, 209.6352, 209.4437, 
    209.2846,
  210.218, 210.4439, 210.5961, 210.7002, 210.8109, 210.83, 210.776, 210.7106, 
    210.6149, 210.5323, 210.4171, 210.2519, 210.0599, 209.8736, 209.7024,
  210.3843, 210.6142, 210.8202, 210.9756, 210.9648, 210.9544, 210.9288, 
    210.9135, 210.8427, 210.7388, 210.6305, 210.5031, 210.3599, 210.2064, 
    210.0475,
  210.5172, 210.7623, 210.9383, 211.0895, 211.1614, 211.1874, 211.1654, 
    211.1123, 211.0558, 210.9624, 210.8136, 210.6864, 210.5448, 210.3988, 
    210.2482,
  207.2536, 207.3285, 207.4199, 207.5959, 207.7952, 207.9931, 208.1539, 
    208.2517, 208.2968, 208.3173, 208.324, 208.3258, 208.3316, 208.3458, 
    208.3607,
  207.0897, 207.3952, 207.5587, 207.6099, 207.6685, 207.7838, 207.942, 
    208.0791, 208.1735, 208.235, 208.2686, 208.2868, 208.2906, 208.2858, 
    208.2717,
  207.0823, 207.4742, 207.7388, 207.8612, 207.8594, 207.8676, 207.9313, 
    208.017, 208.0885, 208.1498, 208.1864, 208.2204, 208.2567, 208.2923, 
    208.3186,
  207.1374, 207.53, 207.8817, 208.0512, 208.1147, 208.0705, 208.0488, 
    208.0667, 208.0922, 208.0951, 208.0813, 208.0749, 208.1042, 208.1512, 
    208.2041,
  207.1706, 207.4873, 207.8812, 208.1549, 208.2192, 208.2336, 208.2159, 
    208.2123, 208.2144, 208.205, 208.1553, 208.1052, 208.09, 208.1281, 
    208.1841,
  207.3678, 207.5959, 207.9212, 208.2966, 208.4293, 208.4205, 208.3686, 
    208.3295, 208.3244, 208.3104, 208.2401, 208.1378, 208.0778, 208.0777, 
    208.1135,
  207.5192, 207.7563, 207.9948, 208.3206, 208.6288, 208.7354, 208.6942, 
    208.6032, 208.5398, 208.5044, 208.4367, 208.3236, 208.219, 208.172, 
    208.168,
  207.7457, 207.9807, 208.2034, 208.4398, 208.7596, 208.9143, 208.9661, 
    208.9283, 208.8163, 208.7398, 208.6625, 208.5556, 208.429, 208.3307, 
    208.2752,
  207.9909, 208.193, 208.4489, 208.7456, 208.9435, 209.1023, 209.1913, 
    209.2492, 209.1715, 209.0403, 208.9359, 208.8446, 208.7377, 208.6173, 
    208.5069,
  208.2318, 208.4227, 208.6268, 208.9507, 209.2139, 209.4333, 209.5216, 
    209.5215, 209.5034, 209.4005, 209.2267, 209.1278, 209.0231, 208.9175, 
    208.7926,
  207.5095, 207.5643, 207.3852, 207.2794, 207.2186, 207.1904, 207.1791, 
    207.1614, 207.1136, 207.0497, 206.9636, 206.8764, 206.798, 206.7482, 
    206.7206,
  207.3255, 207.565, 207.5287, 207.4012, 207.2341, 207.1253, 207.0572, 
    207.0183, 206.9754, 206.9132, 206.832, 206.7464, 206.6703, 206.6129, 
    206.576,
  207.2708, 207.6019, 207.7373, 207.7447, 207.5364, 207.3319, 207.1919, 
    207.091, 207.0095, 206.9168, 206.8242, 206.735, 206.6579, 206.5975, 
    206.5539,
  207.2076, 207.5519, 207.8141, 207.9627, 207.868, 207.6602, 207.4432, 
    207.2821, 207.1546, 207.0298, 206.9018, 206.7799, 206.6832, 206.6118, 
    206.5527,
  207.1926, 207.3964, 207.7203, 208.0457, 208.0381, 207.9198, 207.7391, 
    207.5843, 207.4549, 207.3203, 207.163, 207.0027, 206.8699, 206.7735, 
    206.7032,
  207.316, 207.4174, 207.5871, 207.9941, 208.1224, 208.0723, 207.9291, 
    207.8047, 207.7255, 207.637, 207.4904, 207.3046, 207.1247, 207.0023, 
    206.9194,
  207.3259, 207.4589, 207.5452, 207.8593, 208.1743, 208.2483, 208.1813, 
    208.0374, 207.9478, 207.8982, 207.7994, 207.6204, 207.4224, 207.2755, 
    207.188,
  207.2576, 207.3964, 207.5354, 207.7262, 208.0905, 208.2571, 208.3224, 
    208.3111, 208.1809, 208.1142, 208.0464, 207.9064, 207.7049, 207.5293, 
    207.414,
  207.1495, 207.2433, 207.395, 207.6126, 207.8148, 208.1107, 208.2876, 
    208.47, 208.4652, 208.3782, 208.2931, 208.1927, 208.0424, 207.8781, 
    207.7454,
  207.1106, 207.1844, 207.2751, 207.4508, 207.6133, 207.8778, 208.1497, 
    208.3425, 208.5072, 208.521, 208.3962, 208.3105, 208.1931, 208.078, 
    207.9731,
  209.3265, 209.5369, 209.5142, 209.5038, 209.5182, 209.5667, 209.6289, 
    209.6981, 209.7472, 209.778, 209.793, 209.8018, 209.8114, 209.8181, 
    209.8166,
  208.8313, 209.2584, 209.3716, 209.3886, 209.3607, 209.3679, 209.4034, 
    209.4618, 209.5255, 209.5767, 209.6089, 209.6259, 209.6405, 209.6436, 
    209.6473,
  208.3611, 208.822, 209.0184, 209.2116, 209.248, 209.2661, 209.3013, 
    209.3495, 209.4043, 209.4511, 209.476, 209.4863, 209.4859, 209.4869, 
    209.4825,
  208.1841, 208.5048, 208.7037, 208.9507, 209.0712, 209.148, 209.209, 
    209.2903, 209.3752, 209.4384, 209.4561, 209.4376, 209.4032, 209.3733, 
    209.3532,
  207.867, 208.1395, 208.3039, 208.6033, 208.7457, 208.8516, 208.9326, 
    209.0333, 209.1542, 209.2614, 209.3056, 209.2919, 209.2623, 209.2377, 
    209.2206,
  207.634, 207.8485, 207.9591, 208.3151, 208.5024, 208.612, 208.6734, 
    208.7686, 208.8948, 209.0124, 209.0596, 209.0366, 208.9953, 208.9736, 
    208.9775,
  207.2736, 207.4738, 207.5817, 207.8902, 208.195, 208.3752, 208.4637, 
    208.509, 208.5741, 208.6643, 208.7194, 208.7019, 208.6644, 208.6559, 
    208.6842,
  207.0494, 207.1573, 207.2568, 207.4891, 207.8033, 208.043, 208.169, 
    208.2698, 208.281, 208.3481, 208.4101, 208.4225, 208.3939, 208.3907, 
    208.4259,
  206.9071, 206.9457, 207.0128, 207.2462, 207.3948, 207.6816, 207.8629, 
    208.0281, 208.0427, 208.028, 208.0536, 208.1082, 208.1426, 208.1839, 
    208.2401,
  206.9181, 206.9019, 206.8691, 207.0147, 207.1524, 207.4236, 207.6706, 
    207.785, 207.8667, 207.9014, 207.855, 207.9157, 207.9634, 208.0409, 
    208.0994,
  210.6956, 210.9047, 210.8468, 210.7883, 210.7032, 210.6437, 210.6236, 
    210.6158, 210.5927, 210.531, 210.4317, 210.31, 210.192, 210.0865, 209.9788,
  210.2982, 210.5889, 210.5523, 210.525, 210.4082, 210.3119, 210.2617, 
    210.2432, 210.2246, 210.1684, 210.0801, 209.96, 209.8448, 209.7458, 
    209.6587,
  210.0208, 210.3293, 210.2675, 210.2846, 210.1693, 210.0745, 210.0176, 
    210.0016, 209.9849, 209.9298, 209.8327, 209.7012, 209.5766, 209.4712, 
    209.395,
  209.8692, 210.108, 210.0254, 210.0559, 209.9359, 209.8396, 209.7819, 
    209.7817, 209.7879, 209.7543, 209.6625, 209.5223, 209.3913, 209.2939, 
    209.2278,
  209.6765, 209.8997, 209.8328, 209.8569, 209.7259, 209.6514, 209.6024, 
    209.6124, 209.6314, 209.6124, 209.5224, 209.3855, 209.2523, 209.1683, 
    209.1217,
  209.5488, 209.7174, 209.6671, 209.69, 209.536, 209.4226, 209.376, 209.4053, 
    209.4449, 209.4355, 209.3437, 209.2001, 209.0581, 208.9788, 208.944,
  209.3701, 209.519, 209.4967, 209.4829, 209.3498, 209.2231, 209.1681, 
    209.1798, 209.1996, 209.1884, 209.0976, 208.9593, 208.81, 208.7238, 
    208.6898,
  209.1966, 209.3252, 209.2854, 209.245, 209.1024, 208.9602, 208.8728, 
    208.9036, 208.8718, 208.8485, 208.7712, 208.6531, 208.5127, 208.3954, 
    208.3306,
  208.8922, 208.965, 208.962, 208.9433, 208.6793, 208.4995, 208.4751, 
    208.5315, 208.5033, 208.4238, 208.3452, 208.2571, 208.1613, 208.0619, 
    207.9815,
  208.5924, 208.6103, 208.5459, 208.5164, 208.297, 208.1393, 208.1106, 
    208.1269, 208.16, 208.0922, 207.9614, 207.8979, 207.8268, 207.7611, 
    207.6871,
  210.6361, 210.698, 210.6809, 210.7583, 210.8883, 211.035, 211.1503, 
    211.2111, 211.2191, 211.206, 211.2086, 211.2271, 211.262, 211.2851, 
    211.2792,
  210.1152, 210.2628, 210.2205, 210.2444, 210.3129, 210.4104, 210.5061, 
    210.5556, 210.5775, 210.5721, 210.5725, 210.5887, 210.6249, 210.6554, 
    210.6594,
  209.8469, 210.0262, 209.9434, 209.9362, 209.9489, 209.9993, 210.0568, 
    210.0881, 210.0954, 210.081, 210.0666, 210.0729, 210.1017, 210.1256, 
    210.1247,
  209.6565, 209.7727, 209.6879, 209.6777, 209.6669, 209.6786, 209.675, 
    209.6722, 209.6607, 209.636, 209.6133, 209.6121, 209.6324, 209.6589, 
    209.6666,
  209.4934, 209.6097, 209.5114, 209.4813, 209.4698, 209.4858, 209.4572, 
    209.4179, 209.3813, 209.3462, 209.3089, 209.2832, 209.2832, 209.2991, 
    209.3092,
  209.3464, 209.4559, 209.3865, 209.3634, 209.2984, 209.2744, 209.2448, 
    209.2138, 209.173, 209.125, 209.0704, 209.0188, 208.9867, 208.9828, 
    208.9876,
  209.181, 209.3065, 209.2729, 209.2401, 209.1685, 209.1274, 209.0661, 
    209.032, 209.0018, 208.9745, 208.9324, 208.8769, 208.8225, 208.7983, 
    208.7953,
  209.0136, 209.1309, 209.1051, 209.0725, 209.0317, 208.9632, 208.8864, 
    208.8365, 208.7602, 208.7312, 208.698, 208.6572, 208.606, 208.5555, 
    208.5323,
  208.8196, 208.919, 208.9541, 208.9305, 208.7711, 208.6387, 208.6347, 
    208.6422, 208.5912, 208.527, 208.4774, 208.4317, 208.3835, 208.3243, 
    208.269,
  208.6356, 208.6997, 208.6942, 208.6935, 208.5271, 208.4397, 208.3916, 
    208.3304, 208.3368, 208.2541, 208.1705, 208.1457, 208.1015, 208.0638, 
    208.004,
  209.915, 209.8755, 209.9088, 210.0814, 210.2634, 210.4024, 210.4751, 
    210.4974, 210.4946, 210.4964, 210.5098, 210.541, 210.5771, 210.6037, 
    210.6106,
  209.5095, 209.5409, 209.5306, 209.6225, 209.7701, 209.9243, 210.031, 
    210.089, 210.1122, 210.1258, 210.1466, 210.1734, 210.2079, 210.2365, 
    210.2503,
  209.2056, 209.3289, 209.288, 209.3376, 209.4333, 209.5591, 209.6718, 
    209.7452, 209.7884, 209.8116, 209.8354, 209.863, 209.9015, 209.9311, 
    209.9529,
  209.0222, 209.0844, 209.0417, 209.1012, 209.1597, 209.2419, 209.3319, 
    209.4014, 209.4475, 209.4768, 209.4988, 209.5267, 209.5642, 209.6065, 
    209.6396,
  208.8542, 208.9216, 208.891, 208.9283, 208.9566, 209.0304, 209.1008, 
    209.1637, 209.2127, 209.2382, 209.2514, 209.2689, 209.302, 209.343, 
    209.3853,
  208.7352, 208.8221, 208.7917, 208.8269, 208.8168, 208.8469, 208.892, 
    208.9562, 209.0055, 209.031, 209.0315, 209.0288, 209.0458, 209.0835, 
    209.1351,
  208.6586, 208.7367, 208.7297, 208.77, 208.7387, 208.7417, 208.7438, 
    208.7948, 208.8384, 208.8646, 208.8702, 208.8596, 208.8554, 208.8675, 
    208.8986,
  208.6427, 208.7293, 208.7247, 208.7168, 208.714, 208.6918, 208.6772, 
    208.6838, 208.6754, 208.7101, 208.7289, 208.7281, 208.7114, 208.6972, 
    208.7024,
  208.5861, 208.6883, 208.7498, 208.754, 208.6316, 208.5626, 208.5929, 
    208.6412, 208.5961, 208.5622, 208.5781, 208.596, 208.6005, 208.581, 
    208.5596,
  208.5084, 208.608, 208.6872, 208.7127, 208.6086, 208.5726, 208.5876, 
    208.5505, 208.5676, 208.5138, 208.4644, 208.477, 208.4844, 208.487, 
    208.4595,
  210.5541, 210.6079, 210.5413, 210.5728, 210.5867, 210.5885, 210.5621, 
    210.5214, 210.4584, 210.3782, 210.2834, 210.1777, 210.0656, 209.9546, 
    209.8426,
  210.1664, 210.3113, 210.226, 210.2255, 210.2232, 210.2323, 210.228, 
    210.2115, 210.1881, 210.1518, 210.0933, 210.0246, 209.9399, 209.8439, 
    209.7432,
  209.6825, 209.9476, 209.8882, 209.9284, 209.9267, 209.9285, 209.9249, 
    209.924, 209.925, 209.9214, 209.8998, 209.8624, 209.8132, 209.7516, 
    209.677,
  209.2639, 209.4084, 209.3789, 209.4684, 209.4657, 209.4669, 209.4662, 
    209.4763, 209.4943, 209.5178, 209.5258, 209.5158, 209.4926, 209.4633, 
    209.4253,
  208.7878, 208.9209, 208.9167, 209.0222, 209.0232, 209.0618, 209.0747, 
    209.095, 209.1276, 209.1615, 209.1819, 209.1875, 209.1853, 209.1852, 
    209.1845,
  208.4363, 208.4908, 208.5042, 208.6254, 208.6147, 208.6524, 208.6543, 
    208.6844, 208.7256, 208.7718, 208.7963, 208.8034, 208.8066, 208.8218, 
    208.8461,
  208.1195, 208.1393, 208.1603, 208.2542, 208.2794, 208.3236, 208.3297, 
    208.363, 208.385, 208.4202, 208.4496, 208.4627, 208.4639, 208.4824, 
    208.516,
  207.8453, 207.8727, 207.8773, 207.9221, 207.9642, 207.9967, 208.0077, 
    208.0402, 208.0413, 208.0689, 208.0793, 208.0898, 208.0849, 208.0913, 
    208.1157,
  207.5524, 207.6102, 207.6464, 207.6561, 207.5871, 207.5902, 207.6533, 
    207.7052, 207.6937, 207.6959, 207.7064, 207.7216, 207.7271, 207.7261, 
    207.7304,
  207.2834, 207.3372, 207.3789, 207.3963, 207.3101, 207.3207, 207.3688, 
    207.3387, 207.3326, 207.2972, 207.2823, 207.3094, 207.323, 207.3476, 
    207.3577,
  209.671, 209.8101, 209.9261, 210.0119, 210.0739, 210.1169, 210.1374, 
    210.1407, 210.1237, 210.0902, 210.0368, 209.9748, 209.901, 209.8367, 
    209.7797,
  209.3674, 209.4559, 209.5311, 209.5787, 209.633, 209.6847, 209.7353, 
    209.7694, 209.7911, 209.8042, 209.8054, 209.7909, 209.7502, 209.693, 
    209.6227,
  209.056, 209.1944, 209.2771, 209.3335, 209.3855, 209.4367, 209.5009, 
    209.5618, 209.6105, 209.6463, 209.6638, 209.6672, 209.6541, 209.6253, 
    209.5802,
  208.925, 208.9798, 209.0116, 209.0423, 209.0625, 209.0967, 209.1481, 
    209.2137, 209.2802, 209.3374, 209.3738, 209.3926, 209.399, 209.3963, 
    209.3813,
  208.7802, 208.8178, 208.8355, 208.869, 208.8879, 208.926, 208.9657, 
    209.0205, 209.0834, 209.1378, 209.1775, 209.2055, 209.2312, 209.2536, 
    209.2689,
  208.7597, 208.7652, 208.7408, 208.7596, 208.7473, 208.7745, 208.8219, 
    208.8826, 208.9443, 208.9905, 209.0132, 209.0226, 209.0389, 209.0719, 
    209.1111,
  208.6635, 208.7105, 208.7095, 208.7249, 208.7268, 208.7268, 208.7446, 
    208.7971, 208.858, 208.9124, 208.9438, 208.962, 208.9847, 209.0233, 
    209.0763,
  208.5742, 208.6475, 208.6648, 208.6814, 208.7295, 208.7647, 208.777, 
    208.8087, 208.8206, 208.8524, 208.867, 208.8763, 208.89, 208.926, 208.9852,
  208.4237, 208.503, 208.5627, 208.6042, 208.5845, 208.6078, 208.6878, 
    208.7728, 208.8102, 208.8329, 208.8611, 208.8822, 208.8899, 208.9045, 
    208.9362,
  208.3112, 208.3651, 208.4149, 208.4795, 208.4715, 208.525, 208.5919, 
    208.6137, 208.6596, 208.6745, 208.6832, 208.7288, 208.7562, 208.7852, 
    208.8122,
  208.0487, 208.1061, 208.1605, 208.2122, 208.2654, 208.3104, 208.3468, 
    208.3751, 208.3948, 208.4072, 208.4008, 208.3762, 208.3437, 208.3095, 
    208.2801,
  208.0071, 208.0279, 208.0699, 208.0924, 208.1306, 208.1719, 208.2222, 
    208.2622, 208.2969, 208.3273, 208.3561, 208.3854, 208.4057, 208.4111, 
    208.4017,
  207.8416, 207.9162, 207.9904, 208.0431, 208.0979, 208.1483, 208.2029, 
    208.253, 208.2989, 208.3389, 208.3747, 208.4096, 208.4488, 208.4843, 
    208.5118,
  207.7282, 207.7733, 207.8415, 207.9055, 207.9646, 208.018, 208.0731, 
    208.1296, 208.1831, 208.2261, 208.2647, 208.3, 208.3373, 208.377, 208.4166,
  207.5678, 207.6178, 207.6928, 207.7597, 207.83, 207.9037, 207.9744, 
    208.0381, 208.0967, 208.1436, 208.1826, 208.2173, 208.2529, 208.2908, 
    208.3278,
  207.4073, 207.4769, 207.5541, 207.6201, 207.6772, 207.7424, 207.8197, 
    207.8959, 207.9615, 208.0131, 208.0516, 208.0825, 208.1168, 208.1576, 
    208.199,
  207.2189, 207.3172, 207.3935, 207.452, 207.5236, 207.6041, 207.6779, 
    207.7616, 207.8317, 207.8892, 207.9332, 207.9618, 207.9913, 208.0284, 
    208.0726,
  207.1013, 207.1978, 207.25, 207.2748, 207.3527, 207.4327, 207.5007, 
    207.579, 207.6355, 207.7072, 207.7707, 207.8174, 207.8478, 207.8789, 
    207.9158,
  207.0391, 207.0979, 207.1503, 207.1713, 207.1632, 207.2102, 207.3143, 
    207.4072, 207.4575, 207.5044, 207.5672, 207.6319, 207.6797, 207.7174, 
    207.7544,
  207.0226, 207.0471, 207.0607, 207.081, 207.0527, 207.1092, 207.1961, 
    207.2189, 207.2725, 207.3104, 207.3506, 207.4235, 207.4843, 207.5305, 
    207.5647,
  206.1377, 206.0445, 205.9411, 205.846, 205.7751, 205.7208, 205.6855, 
    205.679, 205.6867, 205.6997, 205.7218, 205.7414, 205.7686, 205.8028, 
    205.8446,
  206.2893, 206.2124, 206.1271, 206.0143, 205.9244, 205.8455, 205.7875, 
    205.7493, 205.7397, 205.7417, 205.7514, 205.7652, 205.7837, 205.8172, 
    205.8525,
  206.4252, 206.3672, 206.2922, 206.1977, 206.1176, 206.0361, 205.9677, 
    205.9074, 205.8624, 205.8425, 205.8394, 205.8543, 205.8701, 205.89, 
    205.9192,
  206.5372, 206.4835, 206.415, 206.3349, 206.2666, 206.1969, 206.1309, 
    206.0683, 206.0084, 205.9632, 205.932, 205.9217, 205.9318, 205.9507, 
    205.976,
  206.6219, 206.5827, 206.5321, 206.4593, 206.4002, 206.3468, 206.297, 
    206.2438, 206.1907, 206.1365, 206.0896, 206.0516, 206.0354, 206.042, 
    206.0622,
  206.6886, 206.6622, 206.6258, 206.5742, 206.5237, 206.4731, 206.4323, 
    206.3928, 206.3501, 206.304, 206.2563, 206.2116, 206.1752, 206.1615, 
    206.1694,
  206.7087, 206.7111, 206.6938, 206.6521, 206.6236, 206.5944, 206.5641, 
    206.5378, 206.5088, 206.4753, 206.4339, 206.39, 206.3522, 206.3279, 
    206.3236,
  206.6838, 206.7209, 206.7154, 206.6811, 206.6822, 206.6705, 206.6698, 
    206.6631, 206.6424, 206.6291, 206.6092, 206.5737, 206.5357, 206.5076, 
    206.4955,
  206.609, 206.6666, 206.7067, 206.6916, 206.6638, 206.6653, 206.7085, 
    206.7373, 206.7431, 206.7386, 206.7434, 206.7414, 206.7245, 206.6995, 
    206.6835,
  206.5208, 206.5785, 206.6325, 206.6618, 206.6562, 206.6939, 206.7435, 
    206.7614, 206.7921, 206.801, 206.8134, 206.8419, 206.8549, 206.8595, 
    206.8518,
  206.2088, 206.153, 206.0822, 206.0354, 205.9993, 205.954, 205.8826, 
    205.782, 205.6622, 205.5326, 205.3981, 205.2617, 205.124, 204.9915, 
    204.868,
  206.2343, 206.2005, 206.1337, 206.0492, 206.0129, 205.9761, 205.9341, 
    205.8685, 205.7845, 205.6816, 205.569, 205.4495, 205.3288, 205.2021, 
    205.0846,
  206.2932, 206.2803, 206.2103, 206.1158, 206.0587, 206.0175, 205.9842, 
    205.927, 205.8602, 205.7835, 205.7066, 205.6163, 205.5114, 205.3963, 
    205.2831,
  206.3533, 206.3357, 206.2801, 206.1994, 206.1357, 206.0858, 206.0472, 
    205.999, 205.9394, 205.8721, 205.8049, 205.7433, 205.6688, 205.581, 
    205.4784,
  206.4044, 206.3905, 206.3522, 206.2752, 206.2241, 206.1847, 206.1457, 
    206.1016, 206.0444, 205.9765, 205.9125, 205.8546, 205.8002, 205.737, 
    205.6619,
  206.4587, 206.4459, 206.412, 206.3559, 206.3083, 206.2703, 206.2437, 
    206.2144, 206.1727, 206.1117, 206.0445, 205.9779, 205.9229, 205.8709, 
    205.8149,
  206.5275, 206.5154, 206.4735, 206.4156, 206.3779, 206.3471, 206.3214, 
    206.3097, 206.2958, 206.2617, 206.208, 206.1358, 206.0706, 206.0089, 
    205.9544,
  206.6027, 206.5954, 206.5542, 206.483, 206.4528, 206.4191, 206.3986, 
    206.3873, 206.371, 206.3659, 206.3507, 206.3062, 206.2523, 206.19, 206.131,
  206.6608, 206.659, 206.6437, 206.5772, 206.5096, 206.4704, 206.4678, 
    206.4684, 206.4427, 206.4253, 206.424, 206.4128, 206.3856, 206.3462, 
    206.3016,
  206.7084, 206.7071, 206.6891, 206.6504, 206.607, 206.5776, 206.558, 
    206.5468, 206.5345, 206.5105, 206.4983, 206.5062, 206.4976, 206.4719, 
    206.4438,
  206.2244, 206.3322, 206.4024, 206.4176, 206.4347, 206.426, 206.4203, 
    206.3701, 206.3076, 206.2404, 206.1808, 206.1155, 206.04, 205.9621, 
    205.8884,
  206.175, 206.2785, 206.3535, 206.387, 206.4372, 206.4287, 206.4586, 
    206.4387, 206.3986, 206.3327, 206.2695, 206.2055, 206.132, 206.0523, 
    205.9765,
  206.1863, 206.2908, 206.3608, 206.391, 206.4297, 206.4286, 206.4709, 
    206.4921, 206.481, 206.4355, 206.3868, 206.3375, 206.28, 206.2093, 
    206.1329,
  206.2162, 206.2791, 206.3728, 206.4075, 206.4292, 206.4109, 206.4532, 
    206.4904, 206.5017, 206.4769, 206.4469, 206.414, 206.3779, 206.3267, 
    206.2625,
  206.272, 206.318, 206.3787, 206.3934, 206.4133, 206.4194, 206.4666, 
    206.5133, 206.5256, 206.4995, 206.4599, 206.4307, 206.4024, 206.3707, 
    206.3252,
  206.3091, 206.4035, 206.4427, 206.446, 206.4253, 206.4247, 206.471, 
    206.5198, 206.5523, 206.5378, 206.4985, 206.4652, 206.4374, 206.4132, 
    206.3802,
  206.3509, 206.4234, 206.4329, 206.4301, 206.4328, 206.4342, 206.4623, 
    206.5081, 206.5518, 206.5551, 206.5369, 206.4978, 206.4667, 206.443, 
    206.4241,
  206.351, 206.428, 206.4572, 206.46, 206.4571, 206.45, 206.4825, 206.5156, 
    206.5262, 206.5396, 206.5419, 206.528, 206.5018, 206.4786, 206.4618,
  206.306, 206.3806, 206.448, 206.4528, 206.4092, 206.4068, 206.4628, 
    206.507, 206.5074, 206.4986, 206.5188, 206.5391, 206.5362, 206.5233, 
    206.5084,
  206.2843, 206.3297, 206.3607, 206.4093, 206.4256, 206.4288, 206.4618, 
    206.4801, 206.5034, 206.4815, 206.4803, 206.521, 206.5397, 206.5408, 
    206.5312,
  207.3869, 207.3636, 207.4485, 207.5054, 207.5495, 207.5863, 207.6264, 
    207.6587, 207.6971, 207.7342, 207.7495, 207.729, 207.6741, 207.6086, 
    207.5526,
  207.1861, 207.2718, 207.3603, 207.3606, 207.3792, 207.384, 207.4303, 
    207.4822, 207.5418, 207.5816, 207.603, 207.6005, 207.56, 207.4966, 
    207.4231,
  207.1737, 207.3349, 207.362, 207.375, 207.3315, 207.2915, 207.3231, 
    207.3813, 207.4431, 207.4847, 207.4989, 207.4857, 207.454, 207.396, 
    207.326,
  207.2269, 207.3218, 207.3782, 207.3904, 207.3478, 207.283, 207.2803, 
    207.332, 207.3994, 207.4342, 207.4381, 207.4236, 207.4014, 207.3704, 
    207.3181,
  207.3376, 207.3707, 207.4208, 207.4247, 207.3748, 207.3359, 207.3037, 
    207.3443, 207.3908, 207.4128, 207.3967, 207.3643, 207.3388, 207.3195, 
    207.2887,
  207.3633, 207.4214, 207.4581, 207.5019, 207.445, 207.4118, 207.3912, 
    207.4301, 207.4757, 207.479, 207.4382, 207.3884, 207.3493, 207.3233, 
    207.3033,
  207.3623, 207.493, 207.5209, 207.549, 207.5234, 207.4882, 207.4786, 
    207.513, 207.5357, 207.5325, 207.4902, 207.4318, 207.3816, 207.3436, 
    207.3226,
  207.3537, 207.4654, 207.5461, 207.5644, 207.598, 207.6063, 207.6099, 
    207.6689, 207.6648, 207.6656, 207.6241, 207.5729, 207.5128, 207.4621, 
    207.4218,
  207.376, 207.4796, 207.5675, 207.6344, 207.5792, 207.6173, 207.7007, 
    207.7819, 207.8112, 207.7983, 207.7614, 207.7237, 207.6807, 207.6323, 
    207.5786,
  207.4451, 207.5163, 207.5416, 207.5916, 207.5657, 207.6069, 207.7322, 
    207.8333, 207.9016, 207.9147, 207.8544, 207.8093, 207.7663, 207.72, 
    207.669,
  208.9707, 208.9676, 208.9302, 208.9133, 208.841, 208.7342, 208.6169, 
    208.5402, 208.5167, 208.5178, 208.5192, 208.4879, 208.4038, 208.2775, 
    208.14,
  208.9985, 209.0626, 209.0481, 209.0213, 208.9193, 208.7904, 208.6576, 
    208.5683, 208.5329, 208.5223, 208.5018, 208.4441, 208.3389, 208.2037, 
    208.0733,
  209.1181, 209.1936, 209.1724, 209.1465, 209.0265, 208.871, 208.7184, 
    208.6153, 208.573, 208.5606, 208.5326, 208.4549, 208.326, 208.1689, 
    208.0314,
  209.2321, 209.2957, 209.284, 209.2592, 209.1414, 208.9736, 208.8115, 
    208.7031, 208.6547, 208.6361, 208.5972, 208.4985, 208.354, 208.1854, 
    208.0533,
  209.3359, 209.3878, 209.3768, 209.3568, 209.2392, 209.0798, 208.9216, 
    208.8139, 208.7685, 208.7455, 208.6954, 208.5916, 208.4451, 208.2927, 
    208.1758,
  209.4562, 209.4832, 209.4534, 209.4383, 209.3154, 209.1482, 209.0038, 
    208.9134, 208.8877, 208.8719, 208.812, 208.6938, 208.5366, 208.3974, 
    208.3064,
  209.5448, 209.5661, 209.5179, 209.477, 209.3576, 209.1945, 209.0577, 
    208.9783, 208.9638, 208.9634, 208.9049, 208.7805, 208.6194, 208.4825, 
    208.4144,
  209.5861, 209.5994, 209.5348, 209.4685, 209.3475, 209.1917, 209.0643, 
    209.0038, 208.9881, 209.002, 208.9715, 208.8658, 208.7205, 208.5818, 
    208.5196,
  209.5888, 209.5942, 209.5355, 209.4633, 209.3022, 209.1496, 209.0523, 
    209.0111, 208.987, 208.9673, 208.9346, 208.8467, 208.7437, 208.6435, 
    208.6057,
  209.5801, 209.5638, 209.4825, 209.395, 209.2464, 209.1202, 209.0504, 
    209.0237, 209.0353, 208.9958, 208.9283, 208.8421, 208.7544, 208.6953, 
    208.6818,
  208.8559, 208.9088, 208.9097, 208.8638, 208.8008, 208.7346, 208.6934, 
    208.6948, 208.7373, 208.8051, 208.8842, 208.9563, 209.009, 209.0412, 
    209.0603,
  208.9446, 209.0102, 209.009, 208.9598, 208.8971, 208.837, 208.8052, 
    208.8119, 208.8495, 208.9047, 208.9532, 208.9851, 208.997, 208.9971, 
    209.0011,
  209.041, 209.1432, 209.1638, 209.1395, 209.0895, 209.0452, 209.023, 
    209.0295, 209.0587, 209.0953, 209.1148, 209.1102, 209.0803, 209.0527, 
    209.0372,
  209.207, 209.2951, 209.2989, 209.2735, 209.2246, 209.1802, 209.1576, 
    209.1596, 209.1842, 209.2085, 209.2124, 209.188, 209.143, 209.1066, 
    209.0951,
  209.3787, 209.4964, 209.4977, 209.4764, 209.4223, 209.3665, 209.3311, 
    209.3175, 209.3352, 209.3516, 209.3543, 209.3225, 209.2834, 209.2546, 
    209.2638,
  209.5554, 209.6933, 209.7052, 209.6754, 209.6035, 209.5265, 209.4772, 
    209.4563, 209.473, 209.4889, 209.4925, 209.466, 209.4339, 209.4191, 
    209.4479,
  209.6977, 209.8501, 209.8833, 209.8637, 209.8077, 209.7374, 209.6896, 
    209.6803, 209.7134, 209.7402, 209.7497, 209.7185, 209.6818, 209.6685, 
    209.6973,
  209.8197, 209.9745, 210.0074, 210.0002, 209.9471, 209.903, 209.8742, 
    209.9021, 209.9566, 210.0093, 210.0279, 210.0014, 209.9565, 209.9294, 
    209.9418,
  209.8885, 210.032, 210.0788, 210.0977, 210.0307, 210.0021, 210.0218, 
    210.0952, 210.1847, 210.2429, 210.2673, 210.2454, 210.2042, 210.1617, 
    210.158,
  209.9482, 210.0699, 210.0911, 210.1087, 210.0693, 210.0603, 210.0982, 
    210.179, 210.2884, 210.3515, 210.3537, 210.3253, 210.2793, 210.243, 
    210.2285,
  208.6814, 208.6975, 208.6636, 208.5963, 208.5096, 208.442, 208.4185, 
    208.4088, 208.4094, 208.3952, 208.3694, 208.3534, 208.3337, 208.3114, 
    208.2847,
  208.8568, 208.9296, 208.9057, 208.8213, 208.7179, 208.6387, 208.6047, 
    208.5972, 208.5972, 208.5784, 208.5418, 208.5032, 208.4692, 208.445, 
    208.4272,
  209.0041, 209.0957, 209.085, 209.0164, 208.9219, 208.851, 208.8231, 
    208.8198, 208.8192, 208.8009, 208.7579, 208.7095, 208.6725, 208.6472, 
    208.6237,
  209.2484, 209.2989, 209.2885, 209.2174, 209.1267, 209.0431, 209.0031, 
    208.9976, 209.0045, 208.9937, 208.9623, 208.9238, 208.8925, 208.8656, 
    208.8398,
  209.5396, 209.5859, 209.5602, 209.4674, 209.3579, 209.2643, 209.2237, 
    209.2214, 209.2308, 209.2251, 209.1976, 209.1655, 209.1448, 209.1306, 
    209.118,
  209.8503, 209.8947, 209.8481, 209.7568, 209.6364, 209.534, 209.4883, 
    209.4971, 209.5192, 209.5142, 209.472, 209.42, 209.3817, 209.3652, 
    209.3583,
  210.1349, 210.1802, 210.1496, 210.0417, 209.9281, 209.8228, 209.7637, 
    209.7697, 209.7865, 209.783, 209.7338, 209.6681, 209.6088, 209.5775, 
    209.5674,
  210.3275, 210.3817, 210.3685, 210.2634, 210.1429, 210.0298, 209.9739, 
    209.9889, 210.0131, 210.0136, 209.966, 209.8987, 209.832, 209.787, 
    209.7615,
  210.4338, 210.493, 210.5234, 210.4577, 210.2941, 210.184, 210.157, 
    210.1745, 210.1898, 210.1731, 210.1333, 210.0753, 210.0252, 209.9875, 
    209.9691,
  210.4816, 210.5405, 210.5552, 210.5132, 210.3931, 210.2916, 210.2485, 
    210.2899, 210.3235, 210.3086, 210.2573, 210.2128, 210.1792, 210.1646, 
    210.1642,
  210.9156, 210.8719, 210.7451, 210.5851, 210.4288, 210.2891, 210.1879, 
    210.1053, 210.0256, 209.9392, 209.8498, 209.7633, 209.6751, 209.5845, 
    209.4918,
  211.021, 211.0618, 210.9955, 210.8716, 210.7361, 210.6086, 210.5157, 
    210.4447, 210.3682, 210.2783, 210.174, 210.0637, 209.9495, 209.833, 
    209.7262,
  211.1145, 211.2323, 211.2286, 211.1615, 211.06, 210.9531, 210.8685, 
    210.8116, 210.7565, 210.6795, 210.5694, 210.448, 210.319, 210.1976, 210.09,
  211.1599, 211.2814, 211.3247, 211.3094, 211.263, 211.1938, 211.1237, 
    211.0746, 211.0317, 210.9584, 210.8433, 210.7074, 210.5677, 210.4423, 
    210.335,
  211.1207, 211.2099, 211.2746, 211.3253, 211.331, 211.2887, 211.2296, 
    211.1884, 211.1577, 211.0984, 210.9819, 210.8356, 210.6873, 210.5695, 
    210.4775,
  211.0257, 211.1498, 211.2132, 211.3105, 211.3718, 211.3805, 211.3478, 
    211.3273, 211.3204, 211.2718, 211.1529, 210.9954, 210.8439, 210.7308, 
    210.6441,
  210.8237, 210.9813, 211.0507, 211.1266, 211.2839, 211.3503, 211.3735, 
    211.3817, 211.3954, 211.3703, 211.2804, 211.1395, 210.993, 210.8721, 
    210.774,
  210.6887, 210.7968, 210.8266, 210.8633, 211.0236, 211.1479, 211.2412, 
    211.3305, 211.3632, 211.3667, 211.3094, 211.1891, 211.0492, 210.9174, 
    210.8084,
  210.5749, 210.6617, 210.671, 210.6756, 210.6982, 210.8438, 211.0266, 
    211.1626, 211.2243, 211.2163, 211.187, 211.1209, 211.0155, 210.9053, 
    210.8023,
  210.4465, 210.5368, 210.4961, 210.4508, 210.4907, 210.6177, 210.8295, 
    211.0273, 211.1308, 211.1314, 211.0638, 211.0073, 210.9089, 210.8046, 
    210.6984,
  211.2656, 211.2911, 211.3216, 211.3428, 211.3591, 211.3698, 211.3909, 
    211.4124, 211.4173, 211.4174, 211.3944, 211.3522, 211.3036, 211.245, 
    211.1667,
  211.001, 211.1722, 211.2633, 211.3071, 211.3155, 211.3134, 211.3225, 
    211.3409, 211.3374, 211.326, 211.2931, 211.2416, 211.1814, 211.1117, 
    211.0407,
  210.9098, 211.1668, 211.3241, 211.4592, 211.5, 211.5122, 211.5213, 
    211.5376, 211.5462, 211.5393, 211.499, 211.4455, 211.3739, 211.2947, 
    211.2077,
  210.8473, 211.0693, 211.2762, 211.4679, 211.5807, 211.6176, 211.6412, 
    211.6685, 211.7033, 211.7159, 211.6957, 211.6337, 211.5607, 211.4716, 
    211.3725,
  210.8361, 210.9695, 211.176, 211.4138, 211.5757, 211.6432, 211.6821, 
    211.7197, 211.7591, 211.7889, 211.77, 211.711, 211.6228, 211.5176, 
    211.4107,
  210.8344, 210.9463, 211.0612, 211.3161, 211.5442, 211.6949, 211.7654, 
    211.8327, 211.8824, 211.9145, 211.8816, 211.8035, 211.6964, 211.5831, 
    211.4686,
  210.8627, 210.9556, 211.0162, 211.1298, 211.4048, 211.6225, 211.7727, 
    211.8601, 211.9378, 211.9588, 211.92, 211.8255, 211.7015, 211.574, 
    211.4475,
  210.9781, 211.0474, 211.0695, 211.0697, 211.2739, 211.4974, 211.6902, 
    211.8464, 211.9395, 211.9917, 211.9422, 211.8353, 211.6893, 211.5438, 
    211.3956,
  211.0612, 211.1111, 211.0947, 211.0891, 211.0917, 211.2775, 211.53, 
    211.7143, 211.8356, 211.8858, 211.8724, 211.7699, 211.6181, 211.4571, 
    211.2967,
  211.142, 211.1789, 211.1234, 211.0789, 211.0636, 211.1213, 211.3134, 
    211.5234, 211.6705, 211.7375, 211.714, 211.6316, 211.4663, 211.2943, 
    211.1237,
  209.8754, 209.96, 210.0385, 210.1466, 210.2245, 210.2787, 210.3424, 
    210.4052, 210.46, 210.5015, 210.5199, 210.5263, 210.5249, 210.5204, 
    210.5142,
  209.6707, 209.8337, 209.9216, 210.0152, 210.0543, 210.0697, 210.0994, 
    210.1357, 210.1752, 210.2057, 210.2292, 210.2465, 210.2637, 210.2731, 
    210.2734,
  209.5716, 209.8004, 209.9225, 210.0287, 210.0541, 210.0531, 210.0667, 
    210.0866, 210.1161, 210.1394, 210.149, 210.1358, 210.1182, 210.1037, 
    210.0955,
  209.4562, 209.638, 209.7636, 209.8739, 209.9233, 209.9351, 209.932, 
    209.9486, 209.9726, 209.988, 209.9865, 209.9648, 209.9323, 209.895, 
    209.8612,
  209.3402, 209.4742, 209.6012, 209.7323, 209.8015, 209.8531, 209.8818, 
    209.9049, 209.9274, 209.9359, 209.9109, 209.8616, 209.8083, 209.7657, 
    209.724,
  209.1817, 209.3182, 209.4382, 209.5795, 209.6616, 209.7197, 209.7715, 
    209.8091, 209.854, 209.8751, 209.8415, 209.7588, 209.6762, 209.6195, 
    209.5859,
  209.0226, 209.1565, 209.2738, 209.3829, 209.5773, 209.6849, 209.7582, 
    209.789, 209.8373, 209.8903, 209.8814, 209.7926, 209.681, 209.6052, 
    209.5815,
  208.9326, 209.0579, 209.1753, 209.3085, 209.5009, 209.6436, 209.7201, 
    209.7938, 209.8183, 209.8773, 209.9186, 209.8697, 209.7639, 209.6607, 
    209.6085,
  208.8434, 208.9378, 209.0553, 209.2696, 209.3342, 209.5859, 209.7905, 
    209.9447, 209.9846, 209.9641, 209.9937, 210.0063, 209.9475, 209.8465, 
    209.7661,
  208.7685, 208.8286, 208.9261, 209.0964, 209.2994, 209.5659, 209.8877, 
    210.1341, 210.2346, 210.1849, 210.1147, 210.1341, 210.1034, 210.0275, 
    209.9211,
  208.7064, 208.7591, 208.7578, 208.7078, 208.6529, 208.6085, 208.5921, 
    208.6044, 208.6397, 208.6849, 208.7241, 208.7565, 208.776, 208.7879, 
    208.7995,
  208.5143, 208.6222, 208.6724, 208.6484, 208.6063, 208.5827, 208.5805, 
    208.6167, 208.6683, 208.7277, 208.7823, 208.8236, 208.8508, 208.8663, 
    208.88,
  208.4443, 208.5619, 208.6204, 208.6072, 208.5768, 208.5601, 208.5813, 
    208.6424, 208.7177, 208.7903, 208.8496, 208.8929, 208.9276, 208.953, 
    208.9739,
  208.3839, 208.4709, 208.518, 208.5177, 208.4951, 208.4843, 208.5138, 
    208.588, 208.6803, 208.7643, 208.8276, 208.8761, 208.9148, 208.9549, 
    208.988,
  208.2793, 208.3816, 208.414, 208.4192, 208.4091, 208.4229, 208.466, 
    208.5534, 208.6542, 208.7466, 208.8077, 208.8495, 208.8872, 208.9347, 
    208.987,
  208.235, 208.3163, 208.3113, 208.3045, 208.282, 208.3049, 208.3684, 
    208.4728, 208.5847, 208.6812, 208.7433, 208.782, 208.818, 208.8732, 
    208.9413,
  208.1775, 208.2685, 208.2485, 208.2125, 208.1903, 208.2209, 208.2829, 
    208.3961, 208.5143, 208.6158, 208.6853, 208.7269, 208.762, 208.8165, 
    208.8926,
  208.1686, 208.2524, 208.2244, 208.1613, 208.1358, 208.158, 208.2241, 
    208.3293, 208.4183, 208.5056, 208.5717, 208.6237, 208.6662, 208.7194, 
    208.7939,
  208.206, 208.2707, 208.2605, 208.2147, 208.1439, 208.1549, 208.2499, 
    208.3562, 208.4186, 208.4452, 208.4693, 208.5075, 208.5469, 208.5863, 
    208.6368,
  208.291, 208.3314, 208.3185, 208.2952, 208.2595, 208.3211, 208.4075, 
    208.4627, 208.5115, 208.5055, 208.4646, 208.4687, 208.4872, 208.5105, 
    208.5281,
  209.7924, 209.8261, 209.8238, 209.7894, 209.7362, 209.6741, 209.613, 
    209.5456, 209.4705, 209.3821, 209.2819, 209.1787, 209.072, 208.9724, 
    208.8878,
  209.8165, 209.8622, 209.8528, 209.7995, 209.7493, 209.702, 209.657, 
    209.6252, 209.5966, 209.546, 209.4824, 209.4051, 209.3137, 209.2168, 
    209.1292,
  209.8147, 209.9094, 209.9304, 209.8891, 209.8418, 209.8024, 209.7741, 
    209.769, 209.7589, 209.7372, 209.7041, 209.6534, 209.5967, 209.5338, 
    209.4645,
  209.7742, 209.8715, 209.9106, 209.8886, 209.8615, 209.8295, 209.8182, 
    209.8221, 209.8288, 209.823, 209.8061, 209.7703, 209.7305, 209.6944, 
    209.6583,
  209.6563, 209.7842, 209.8554, 209.8617, 209.8645, 209.8578, 209.8667, 
    209.8832, 209.8936, 209.8895, 209.8677, 209.8316, 209.8033, 209.7827, 
    209.7623,
  209.5082, 209.6519, 209.7305, 209.768, 209.7828, 209.79, 209.8193, 
    209.8599, 209.8854, 209.8922, 209.8729, 209.8338, 209.8003, 209.777, 
    209.7589,
  209.3303, 209.4788, 209.5617, 209.5973, 209.6258, 209.6547, 209.6991, 
    209.7647, 209.813, 209.8359, 209.827, 209.7928, 209.7591, 209.7288, 
    209.7054,
  209.1752, 209.3066, 209.3898, 209.425, 209.4529, 209.479, 209.5367, 
    209.6165, 209.6712, 209.7071, 209.7034, 209.6794, 209.6515, 209.6236, 
    209.5971,
  209.0509, 209.1646, 209.2586, 209.2941, 209.2912, 209.319, 209.39, 
    209.4709, 209.5172, 209.5307, 209.5253, 209.5125, 209.5029, 209.4839, 
    209.4629,
  208.9766, 209.086, 209.1343, 209.176, 209.2069, 209.2514, 209.3073, 
    209.3363, 209.3743, 209.382, 209.3601, 209.3486, 209.3425, 209.3371, 
    209.3195,
  208.6999, 208.7405, 208.7538, 208.7459, 208.7282, 208.7125, 208.7274, 
    208.7724, 208.8278, 208.8767, 208.9077, 208.9158, 208.9146, 208.9061, 
    208.8781,
  208.6326, 208.731, 208.7895, 208.7581, 208.7057, 208.6605, 208.6414, 
    208.6504, 208.6756, 208.7145, 208.75, 208.7881, 208.8278, 208.8574, 
    208.8694,
  208.7071, 208.7713, 208.8261, 208.8417, 208.7864, 208.7347, 208.7073, 
    208.7013, 208.7014, 208.7177, 208.722, 208.738, 208.7666, 208.7954, 
    208.8273,
  208.873, 208.908, 208.9542, 208.9598, 208.9372, 208.8709, 208.83, 208.8072, 
    208.8087, 208.8052, 208.783, 208.7641, 208.75, 208.7522, 208.7745,
  209.0932, 209.0789, 209.113, 209.1373, 209.0997, 209.0432, 208.9906, 
    208.9667, 208.9608, 208.9467, 208.9191, 208.8908, 208.8638, 208.8526, 
    208.8576,
  209.3096, 209.3108, 209.294, 209.3433, 209.3395, 209.2923, 209.2208, 
    209.1658, 209.1454, 209.1207, 209.0889, 209.045, 209.0015, 208.9781, 
    208.9794,
  209.4042, 209.447, 209.4711, 209.5069, 209.5891, 209.5522, 209.495, 
    209.4275, 209.3851, 209.3376, 209.2828, 209.2243, 209.1669, 209.1267, 
    209.1028,
  209.4139, 209.476, 209.537, 209.5951, 209.7175, 209.7364, 209.7288, 
    209.7045, 209.6665, 209.6174, 209.5536, 209.4762, 209.3985, 209.3331, 
    209.2769,
  209.3572, 209.4347, 209.5246, 209.6231, 209.6751, 209.7916, 209.8535, 
    209.8782, 209.8585, 209.8089, 209.7345, 209.6431, 209.5644, 209.4965, 
    209.4301,
  209.2829, 209.3775, 209.4466, 209.5569, 209.66, 209.8116, 209.9038, 
    209.9937, 209.9703, 209.9261, 209.8483, 209.7846, 209.7231, 209.6679, 
    209.5959,
  208.756, 208.6155, 208.4986, 208.3793, 208.2662, 208.153, 208.0608, 
    207.9708, 207.88, 207.7912, 207.7015, 207.6266, 207.5584, 207.5111, 
    207.4831,
  208.7823, 208.7252, 208.628, 208.5019, 208.3647, 208.2365, 208.124, 
    208.0097, 207.8933, 207.7723, 207.6456, 207.5352, 207.4509, 207.3917, 
    207.3423,
  208.9275, 208.8879, 208.8306, 208.7376, 208.5908, 208.4271, 208.3026, 
    208.1978, 208.0852, 207.954, 207.8048, 207.6658, 207.5391, 207.4405, 
    207.3665,
  209.0757, 209.0795, 209.0975, 209.0172, 208.9157, 208.7332, 208.5754, 
    208.457, 208.3587, 208.2468, 208.1038, 207.9339, 207.7723, 207.6395, 
    207.5335,
  209.1696, 209.2066, 209.2833, 209.3, 209.1945, 209.0252, 208.8265, 
    208.6749, 208.5645, 208.4699, 208.3495, 208.2066, 208.0582, 207.9196, 
    207.7793,
  209.226, 209.3293, 209.3957, 209.5151, 209.5069, 209.3812, 209.1843, 
    208.9933, 208.8608, 208.7481, 208.6197, 208.4734, 208.3229, 208.1812, 
    208.0488,
  209.224, 209.3386, 209.4467, 209.6305, 209.7979, 209.7794, 209.6626, 
    209.4438, 209.2563, 209.0879, 208.9194, 208.7347, 208.5681, 208.4138, 
    208.2843,
  209.3419, 209.34, 209.3983, 209.5418, 209.848, 209.9996, 209.9848, 
    209.8669, 209.682, 209.504, 209.307, 209.0946, 208.8879, 208.7021, 
    208.5515,
  209.5165, 209.4819, 209.4396, 209.5419, 209.7139, 210.0288, 210.172, 
    210.1774, 210.0523, 209.8762, 209.6771, 209.4679, 209.2395, 209.0404, 
    208.8722,
  209.7009, 209.6412, 209.5499, 209.538, 209.701, 209.9416, 210.2357, 
    210.3482, 210.362, 210.2621, 210.0718, 209.872, 209.6253, 209.4119, 
    209.2232,
  210.3077, 210.3582, 210.4239, 210.4779, 210.5305, 210.5705, 210.598, 
    210.629, 210.6472, 210.6661, 210.6868, 210.7129, 210.7428, 210.7961, 
    210.852,
  209.94, 210.1071, 210.2422, 210.3043, 210.3221, 210.3167, 210.3169, 
    210.3224, 210.3309, 210.3316, 210.3252, 210.3068, 210.2878, 210.2736, 
    210.2656,
  209.7152, 209.9403, 210.11, 210.2269, 210.2386, 210.2085, 210.1917, 
    210.2047, 210.2297, 210.2476, 210.246, 210.2308, 210.2052, 210.1708, 
    210.1284,
  209.5732, 209.7967, 209.9817, 210.1232, 210.1878, 210.1796, 210.1596, 
    210.1787, 210.2217, 210.2547, 210.263, 210.2486, 210.2286, 210.2078, 
    210.1771,
  209.5196, 209.684, 209.8677, 210.0511, 210.1289, 210.145, 210.1184, 
    210.1137, 210.1433, 210.1751, 210.1882, 210.1737, 210.1555, 210.1475, 
    210.1378,
  209.5388, 209.6636, 209.804, 210.0101, 210.1615, 210.2426, 210.2506, 
    210.2307, 210.2284, 210.2279, 210.2024, 210.1611, 210.121, 210.0998, 
    210.0892,
  209.5274, 209.6599, 209.7914, 209.9433, 210.1793, 210.3329, 210.4222, 
    210.426, 210.4061, 210.3832, 210.3472, 210.2991, 210.248, 210.2102, 
    210.1814,
  209.6222, 209.7156, 209.8085, 209.9011, 210.1458, 210.3497, 210.4769, 
    210.5331, 210.5235, 210.5005, 210.4792, 210.4436, 210.4039, 210.3595, 
    210.3174,
  209.8482, 209.9201, 209.9632, 210.0407, 210.1503, 210.3761, 210.5807, 
    210.6653, 210.6644, 210.6449, 210.6299, 210.6062, 210.569, 210.516, 
    210.4527,
  210.1187, 210.1818, 210.1938, 210.206, 210.3208, 210.4998, 210.7598, 
    210.9043, 210.9774, 211.0055, 210.995, 210.9774, 210.9348, 210.8819, 
    210.818,
  210.6645, 210.6658, 210.7262, 210.8196, 210.9394, 211.0532, 211.1736, 
    211.3071, 211.4515, 211.591, 211.7334, 211.8699, 212.0138, 212.1515, 
    212.2444,
  210.4733, 210.5237, 210.6017, 210.6606, 210.7194, 210.7829, 210.8493, 
    210.9368, 211.0435, 211.1601, 211.2821, 211.401, 211.5212, 211.6358, 
    211.7258,
  210.4073, 210.4892, 210.5748, 210.6614, 210.7123, 210.7461, 210.7794, 
    210.8228, 210.878, 210.9435, 211.0069, 211.0694, 211.1401, 211.2179, 
    211.2918,
  210.3796, 210.4337, 210.5175, 210.6072, 210.6969, 210.7469, 210.7683, 
    210.7879, 210.8199, 210.8554, 210.8798, 210.8932, 210.9128, 210.9441, 
    210.9852,
  210.3413, 210.3817, 210.4424, 210.5409, 210.6311, 210.6915, 210.7088, 
    210.7132, 210.727, 210.742, 210.7488, 210.737, 210.7312, 210.7415, 
    210.7582,
  210.3539, 210.3837, 210.3965, 210.487, 210.5923, 210.6706, 210.6782, 
    210.6551, 210.634, 210.6253, 210.6087, 210.5808, 210.5485, 210.5349, 
    210.5381,
  210.3479, 210.3704, 210.372, 210.3812, 210.5222, 210.6264, 210.6897, 
    210.6761, 210.6476, 210.6304, 210.6171, 210.5908, 210.5522, 210.519, 
    210.492,
  210.4255, 210.4362, 210.4304, 210.408, 210.4916, 210.593, 210.664, 
    210.6894, 210.6594, 210.6327, 210.6156, 210.5923, 210.5612, 210.521, 
    210.4826,
  210.4783, 210.5154, 210.503, 210.4936, 210.4533, 210.5683, 210.6859, 
    210.7469, 210.7279, 210.6868, 210.6515, 210.6173, 210.5827, 210.541, 
    210.4946,
  210.5552, 210.6261, 210.6199, 210.5736, 210.565, 210.6545, 210.8083, 
    210.8866, 210.9241, 210.9258, 210.8817, 210.8449, 210.8083, 210.7724, 
    210.7313,
  210.6919, 210.7662, 210.8481, 210.9149, 211.0018, 211.0862, 211.1624, 
    211.2486, 211.3514, 211.4592, 211.5629, 211.6676, 211.7784, 211.894, 
    212.0072,
  210.4872, 210.5901, 210.6828, 210.7369, 210.8027, 210.8656, 210.9192, 
    210.974, 211.0406, 211.1169, 211.1924, 211.2662, 211.3472, 211.4384, 
    211.5356,
  210.4118, 210.5455, 210.6476, 210.6988, 210.7575, 210.8058, 210.8413, 
    210.8697, 210.9046, 210.9478, 210.998, 211.0458, 211.1019, 211.1702, 
    211.2492,
  210.3868, 210.4794, 210.5627, 210.6157, 210.6783, 210.7256, 210.7593, 
    210.7854, 210.8157, 210.8509, 210.8878, 210.9245, 210.9695, 211.029, 
    211.1018,
  210.2995, 210.4077, 210.5003, 210.5688, 210.6324, 210.6759, 210.7114, 
    210.7418, 210.7686, 210.8065, 210.8422, 210.8752, 210.9124, 210.9636, 
    211.0272,
  210.2238, 210.3204, 210.3929, 210.4553, 210.5195, 210.5653, 210.61, 
    210.6541, 210.6973, 210.7508, 210.7969, 210.8252, 210.8486, 210.8844, 
    210.9384,
  210.0962, 210.1885, 210.2356, 210.2942, 210.3762, 210.4416, 210.5004, 
    210.5521, 210.5949, 210.6589, 210.7266, 210.7768, 210.8047, 210.8325, 
    210.873,
  210.0383, 210.1106, 210.1294, 210.1636, 210.232, 210.2992, 210.3939, 
    210.5046, 210.5656, 210.6296, 210.6992, 210.7517, 210.7732, 210.7791, 
    210.7996,
  209.9277, 210.0178, 210.0328, 210.0586, 210.0767, 210.1501, 210.3106, 
    210.4702, 210.5643, 210.6103, 210.6668, 210.7197, 210.7453, 210.752, 
    210.7562,
  209.8421, 209.9301, 209.9292, 209.9138, 209.9293, 209.9963, 210.2355, 
    210.4592, 210.6436, 210.7148, 210.7362, 210.7775, 210.8049, 210.8214, 
    210.83,
  211.5671, 211.6026, 211.6424, 211.6655, 211.6846, 211.7009, 211.7142, 
    211.729, 211.7474, 211.7728, 211.7996, 211.819, 211.831, 211.8312, 
    211.8219,
  211.535, 211.5967, 211.6252, 211.6405, 211.6638, 211.6841, 211.7043, 
    211.7215, 211.7426, 211.7646, 211.7849, 211.7912, 211.7814, 211.756, 
    211.7177,
  211.4601, 211.5764, 211.6206, 211.6487, 211.6852, 211.7167, 211.7472, 
    211.7767, 211.811, 211.8452, 211.8697, 211.8779, 211.8628, 211.8252, 
    211.7664,
  211.4326, 211.5076, 211.5391, 211.5646, 211.6018, 211.6397, 211.6764, 
    211.7186, 211.7641, 211.8098, 211.8438, 211.8566, 211.8505, 211.8215, 
    211.7715,
  211.3081, 211.3955, 211.443, 211.4812, 211.5165, 211.5553, 211.5943, 
    211.6374, 211.6882, 211.7381, 211.772, 211.7793, 211.7672, 211.7387, 
    211.6942,
  211.1965, 211.2726, 211.3118, 211.3548, 211.3853, 211.4083, 211.4405, 
    211.4838, 211.5376, 211.59, 211.6201, 211.6117, 211.5871, 211.5607, 
    211.5325,
  211.0367, 211.1067, 211.1438, 211.1889, 211.2334, 211.2595, 211.2838, 
    211.3218, 211.3721, 211.4267, 211.4596, 211.4469, 211.4045, 211.3613, 
    211.3271,
  210.901, 210.9566, 210.9767, 211.0137, 211.0493, 211.0681, 211.0853, 
    211.1159, 211.1454, 211.1941, 211.2447, 211.2552, 211.2155, 211.1588, 
    211.1183,
  210.7287, 210.7746, 210.7931, 210.837, 210.8484, 210.861, 210.8926, 
    210.9274, 210.9496, 210.9594, 210.9945, 211.0296, 211.0224, 210.9806, 
    210.9409,
  210.5868, 210.6122, 210.6154, 210.6465, 210.6827, 210.72, 210.7619, 
    210.7861, 210.8159, 210.81, 210.7989, 210.8215, 210.8348, 210.7982, 
    210.7468,
  211.756, 211.7987, 211.8261, 211.831, 211.7992, 211.7542, 211.6877, 
    211.6076, 211.5232, 211.4399, 211.3707, 211.3103, 211.2578, 211.2041, 
    211.1617,
  211.6189, 211.6889, 211.7013, 211.6982, 211.6595, 211.6111, 211.5516, 
    211.4824, 211.4094, 211.3336, 211.2591, 211.1909, 211.1292, 211.0683, 
    211.0125,
  211.4187, 211.5246, 211.5553, 211.5787, 211.5553, 211.5171, 211.4681, 
    211.4175, 211.3673, 211.3126, 211.2487, 211.1777, 211.106, 211.0334, 
    210.9617,
  211.2282, 211.3112, 211.3397, 211.3667, 211.3625, 211.3514, 211.3183, 
    211.2865, 211.2599, 211.2285, 211.1796, 211.1139, 211.0402, 210.9679, 
    210.8931,
  210.9241, 211.0308, 211.0844, 211.1301, 211.1476, 211.1737, 211.1737, 
    211.1661, 211.161, 211.1506, 211.1146, 211.0512, 210.9801, 210.9135, 
    210.8465,
  210.6573, 210.7464, 210.8005, 210.8638, 210.89, 210.924, 210.9529, 
    210.9734, 210.9955, 211.0084, 210.99, 210.9367, 210.873, 210.8179, 
    210.7727,
  210.3605, 210.4471, 210.4988, 210.5642, 210.6132, 210.6633, 210.7027, 
    210.7399, 210.7839, 210.8248, 210.8341, 210.7999, 210.7495, 210.7089, 
    210.6902,
  210.1241, 210.1926, 210.2305, 210.2851, 210.3373, 210.3872, 210.4291, 
    210.4778, 210.5181, 210.5724, 210.6174, 210.6208, 210.595, 210.5693, 
    210.5694,
  209.8791, 209.9346, 209.9763, 210.0418, 210.0641, 210.1115, 210.1695, 
    210.2305, 210.2769, 210.3106, 210.3674, 210.4116, 210.4245, 210.4207, 
    210.4355,
  209.6996, 209.7429, 209.7656, 209.8183, 209.8652, 209.9196, 209.9659, 
    210.0073, 210.062, 210.0937, 210.1267, 210.1898, 210.236, 210.2565, 
    210.2772,
  211.3962, 211.5836, 211.7104, 211.6697, 211.5704, 211.4636, 211.3701, 
    211.3043, 211.27, 211.2736, 211.2978, 211.3235, 211.3317, 211.3126, 
    211.2626,
  211.0911, 211.3293, 211.5958, 211.6821, 211.639, 211.5309, 211.4324, 
    211.3573, 211.3116, 211.2951, 211.2971, 211.2941, 211.2777, 211.2376, 
    211.1769,
  210.8899, 211.1799, 211.49, 211.6682, 211.6843, 211.6021, 211.5286, 
    211.4711, 211.4399, 211.4261, 211.4205, 211.4097, 211.3855, 211.3399, 
    211.2823,
  210.6417, 210.8758, 211.2149, 211.4665, 211.5918, 211.5783, 211.541, 
    211.5167, 211.5158, 211.5153, 211.5087, 211.4842, 211.4499, 211.4011, 
    211.346,
  210.3666, 210.5383, 210.834, 211.1328, 211.2916, 211.3664, 211.3896, 
    211.4192, 211.4555, 211.483, 211.4854, 211.4644, 211.43, 211.3929, 
    211.3521,
  210.2071, 210.3437, 210.4802, 210.7184, 210.8942, 211.0062, 211.0863, 
    211.1743, 211.2639, 211.3365, 211.3654, 211.3592, 211.3302, 211.3032, 
    211.2791,
  209.9942, 210.1215, 210.2219, 210.3633, 210.522, 210.6609, 210.7781, 
    210.9014, 211.0233, 211.1189, 211.161, 211.1616, 211.1401, 211.1266, 
    211.1174,
  209.7131, 209.8507, 209.9258, 210.0184, 210.1377, 210.254, 210.3793, 
    210.5133, 210.6346, 210.7374, 210.8031, 210.8294, 210.8304, 210.8359, 
    210.8503,
  209.3888, 209.5193, 209.6, 209.687, 209.7658, 209.8786, 210.0029, 210.1398, 
    210.2602, 210.3519, 210.4221, 210.4724, 210.4969, 210.5161, 210.542,
  209.0496, 209.1726, 209.2375, 209.323, 209.4197, 209.5242, 209.6281, 
    209.7487, 209.8658, 209.9494, 210.0063, 210.0688, 210.1172, 210.158, 
    210.1941,
  209.769, 209.903, 210.0127, 210.1011, 210.1813, 210.256, 210.3309, 
    210.3996, 210.4532, 210.5017, 210.5372, 210.5643, 210.575, 210.5818, 
    210.5855,
  209.6156, 209.7043, 209.7906, 209.8699, 209.9644, 210.0506, 210.128, 
    210.1988, 210.2516, 210.2874, 210.3143, 210.3315, 210.3481, 210.3611, 
    210.3694,
  209.5276, 209.6556, 209.7685, 209.8572, 209.9461, 210.0202, 210.0999, 
    210.1689, 210.2316, 210.2728, 210.2968, 210.3067, 210.3078, 210.3063, 
    210.3027,
  209.4723, 209.5726, 209.6987, 209.7963, 209.8922, 209.954, 210.0249, 
    210.0872, 210.1453, 210.1841, 210.2041, 210.2125, 210.2126, 210.2076, 
    210.2007,
  209.4316, 209.5165, 209.6638, 209.7995, 209.9126, 209.9846, 210.0435, 
    210.094, 210.1387, 210.1689, 210.183, 210.1826, 210.1759, 210.1652, 
    210.1512,
  209.4365, 209.4757, 209.5883, 209.7384, 209.846, 209.9358, 210.0095, 
    210.065, 210.1045, 210.1317, 210.1407, 210.138, 210.1294, 210.1182, 
    210.1036,
  209.3867, 209.4218, 209.5089, 209.6398, 209.7663, 209.8749, 209.9557, 
    210.0181, 210.0533, 210.0752, 210.0853, 210.0886, 210.0889, 210.0885, 
    210.0876,
  209.2872, 209.3689, 209.4401, 209.5314, 209.6472, 209.7366, 209.8245, 
    209.8973, 209.931, 209.9577, 209.9705, 209.9754, 209.9706, 209.9684, 
    209.9744,
  209.1006, 209.1989, 209.2777, 209.3577, 209.4493, 209.549, 209.6531, 
    209.7222, 209.7563, 209.7808, 209.8037, 209.8246, 209.8322, 209.8356, 
    209.8441,
  208.898, 208.9827, 209.0529, 209.1451, 209.2332, 209.3311, 209.4109, 
    209.4603, 209.5104, 209.5325, 209.5556, 209.5927, 209.6115, 209.6195, 
    209.6279,
  209.3663, 209.5056, 209.5697, 209.6277, 209.6684, 209.7306, 209.8141, 
    209.8894, 209.957, 210.0178, 210.0712, 210.1217, 210.1635, 210.1914, 
    210.2034,
  209.0971, 209.2035, 209.2905, 209.3352, 209.3719, 209.4045, 209.469, 
    209.5433, 209.6139, 209.6706, 209.7149, 209.7543, 209.7878, 209.8139, 
    209.8339,
  208.9158, 209.0037, 209.0921, 209.1467, 209.1868, 209.2123, 209.2725, 
    209.3385, 209.4052, 209.453, 209.4872, 209.52, 209.5439, 209.5641, 
    209.5809,
  208.7262, 208.7732, 208.8866, 208.9637, 209.0143, 209.0209, 209.0598, 
    209.1104, 209.161, 209.1958, 209.215, 209.2361, 209.2564, 209.2786, 
    209.2973,
  208.5413, 208.579, 208.6831, 208.7821, 208.8688, 208.9122, 208.9304, 
    208.9603, 208.9939, 209.0175, 209.0281, 209.0366, 209.0485, 209.0702, 
    209.0905,
  208.3973, 208.4122, 208.4751, 208.605, 208.6939, 208.7451, 208.7966, 
    208.815, 208.8413, 208.8559, 208.8612, 208.8652, 208.873, 208.8878, 
    208.8983,
  208.2301, 208.2592, 208.2947, 208.3725, 208.5409, 208.6117, 208.6703, 
    208.695, 208.7225, 208.7351, 208.7407, 208.7488, 208.7573, 208.7702, 
    208.7779,
  208.0533, 208.0921, 208.1401, 208.1745, 208.3182, 208.4756, 208.5347, 
    208.5913, 208.604, 208.6208, 208.625, 208.6429, 208.6508, 208.66, 208.6677,
  207.8675, 207.9174, 208.0036, 208.0124, 208.0858, 208.2999, 208.4125, 
    208.4985, 208.5326, 208.5511, 208.5619, 208.5804, 208.5893, 208.6045, 
    208.6106,
  207.7378, 207.7787, 207.8366, 207.8958, 207.984, 208.1544, 208.2672, 
    208.3408, 208.4188, 208.4532, 208.4908, 208.5226, 208.5379, 208.5582, 
    208.5643 ;

 time = 0.5, 1.5, 2.5, 3.5, 4.5, 5.5, 6.5, 7.5, 8.5, 9.5, 10.5, 11.5, 12.5, 
    13.5, 14.5, 15.5, 16.5, 17.5, 18.5, 19.5, 20.5, 21.5, 22.5, 23.5, 24.5, 
    25.5, 26.5, 27.5, 28.5, 29.5, 30.5, 31.5, 32.5, 33.5, 34.5, 35.5, 36.5, 
    37.5, 38.5, 39.5, 40.5, 41.5, 42.5, 43.5, 44.5, 45.5, 46.5, 47.5, 48.5, 
    49.5, 50.5, 51.5, 52.5, 53.5, 54.5, 55.5, 56.5, 57.5, 58.5, 59.5, 60.5, 
    61.5, 62.5, 63.5, 64.5, 65.5, 66.5, 67.5, 68.5, 69.5, 70.5, 71.5, 72.5, 
    73.5, 74.5, 75.5, 76.5, 77.5, 78.5, 79.5, 80.5, 81.5, 82.5, 83.5, 84.5, 
    85.5, 86.5, 87.5, 88.5, 89.5, 90.5, 91.5, 92.5, 93.5, 94.5, 95.5, 96.5, 
    97.5, 98.5, 99.5, 100.5, 101.5, 102.5, 103.5, 104.5, 105.5, 106.5, 107.5, 
    108.5, 109.5, 110.5, 111.5, 112.5, 113.5, 114.5, 115.5, 116.5, 117.5, 
    118.5, 119.5, 120.5, 121.5, 122.5, 123.5, 124.5, 125.5, 126.5, 127.5, 
    128.5, 129.5, 130.5, 131.5, 132.5, 133.5, 134.5, 135.5, 136.5, 137.5, 
    138.5, 139.5, 140.5, 141.5, 142.5, 143.5, 144.5, 145.5, 146.5, 147.5, 
    148.5, 149.5, 150.5, 151.5, 152.5, 153.5, 154.5, 155.5, 156.5, 157.5, 
    158.5, 159.5, 160.5, 161.5, 162.5, 163.5, 164.5, 165.5, 166.5, 167.5, 
    168.5, 169.5, 170.5, 171.5, 172.5, 173.5, 174.5, 175.5, 176.5, 177.5, 
    178.5, 179.5, 180.5 ;

 time_bnds =
  0, 1,
  1, 2,
  2, 3,
  3, 4,
  4, 5,
  5, 6,
  6, 7,
  7, 8,
  8, 9,
  9, 10,
  10, 11,
  11, 12,
  12, 13,
  13, 14,
  14, 15,
  15, 16,
  16, 17,
  17, 18,
  18, 19,
  19, 20,
  20, 21,
  21, 22,
  22, 23,
  23, 24,
  24, 25,
  25, 26,
  26, 27,
  27, 28,
  28, 29,
  29, 30,
  30, 31,
  31, 32,
  32, 33,
  33, 34,
  34, 35,
  35, 36,
  36, 37,
  37, 38,
  38, 39,
  39, 40,
  40, 41,
  41, 42,
  42, 43,
  43, 44,
  44, 45,
  45, 46,
  46, 47,
  47, 48,
  48, 49,
  49, 50,
  50, 51,
  51, 52,
  52, 53,
  53, 54,
  54, 55,
  55, 56,
  56, 57,
  57, 58,
  58, 59,
  59, 60,
  60, 61,
  61, 62,
  62, 63,
  63, 64,
  64, 65,
  65, 66,
  66, 67,
  67, 68,
  68, 69,
  69, 70,
  70, 71,
  71, 72,
  72, 73,
  73, 74,
  74, 75,
  75, 76,
  76, 77,
  77, 78,
  78, 79,
  79, 80,
  80, 81,
  81, 82,
  82, 83,
  83, 84,
  84, 85,
  85, 86,
  86, 87,
  87, 88,
  88, 89,
  89, 90,
  90, 91,
  91, 92,
  92, 93,
  93, 94,
  94, 95,
  95, 96,
  96, 97,
  97, 98,
  98, 99,
  99, 100,
  100, 101,
  101, 102,
  102, 103,
  103, 104,
  104, 105,
  105, 106,
  106, 107,
  107, 108,
  108, 109,
  109, 110,
  110, 111,
  111, 112,
  112, 113,
  113, 114,
  114, 115,
  115, 116,
  116, 117,
  117, 118,
  118, 119,
  119, 120,
  120, 121,
  121, 122,
  122, 123,
  123, 124,
  124, 125,
  125, 126,
  126, 127,
  127, 128,
  128, 129,
  129, 130,
  130, 131,
  131, 132,
  132, 133,
  133, 134,
  134, 135,
  135, 136,
  136, 137,
  137, 138,
  138, 139,
  139, 140,
  140, 141,
  141, 142,
  142, 143,
  143, 144,
  144, 145,
  145, 146,
  146, 147,
  147, 148,
  148, 149,
  149, 150,
  150, 151,
  151, 152,
  152, 153,
  153, 154,
  154, 155,
  155, 156,
  156, 157,
  157, 158,
  158, 159,
  159, 160,
  160, 161,
  161, 162,
  162, 163,
  163, 164,
  164, 165,
  165, 166,
  166, 167,
  167, 168,
  168, 169,
  169, 170,
  170, 171,
  171, 172,
  172, 173,
  173, 174,
  174, 175,
  175, 176,
  176, 177,
  177, 178,
  178, 179,
  179, 180,
  180, 181 ;

 zsurf =
  1.522432, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  122.465, 2.830728, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  113.0215, 29.31339, 0.004701966, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  140.0874, 33.71546, 1.141547, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  141.9684, 87.21121, 14.52402, 0.1304746, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  165.7051, 185.2302, 111.1391, 5.227489, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  172.6293, 232.1111, 238.8028, 89.74486, 0.6524738, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  149.5705, 217.5222, 183.4477, 142.7244, 6.651272, 0.2006134, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  253.9191, 270.7406, 160.8987, 135.4378, 83.93595, 3.422685, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  248.2018, 381.5977, 396.3867, 296.0411, 147.8827, 85.51294, 0.2661929, 0, 
    0, 0, 0, 0, 0, 0, 0 ;
}
