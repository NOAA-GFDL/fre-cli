netcdf tracer_level.0003-0003.scale_salt_emis {
dimensions:
	bnds = 2 ;
	lat = 18 ;
	lon = 29 ;
	time = UNLIMITED ; // (1 currently)
variables:
	double bnds(bnds) ;
		bnds:long_name = "vertex number" ;
	double lat(lat) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_N" ;
		lat:axis = "Y" ;
		lat:bounds = "lat_bnds" ;
	double lat_bnds(lat, bnds) ;
		lat_bnds:long_name = "latitude bounds" ;
		lat_bnds:units = "degrees_N" ;
		lat_bnds:axis = "Y" ;
	double lon(lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_E" ;
		lon:axis = "X" ;
		lon:bounds = "lon_bnds" ;
	double lon_bnds(lon, bnds) ;
		lon_bnds:long_name = "longitude bounds" ;
		lon_bnds:units = "degrees_E" ;
		lon_bnds:axis = "X" ;
	float scale_salt_emis(time, lat, lon) ;
		scale_salt_emis:_FillValue = 1.e+20f ;
		scale_salt_emis:missing_value = 1.e+20f ;
		scale_salt_emis:units = "unitless" ;
		scale_salt_emis:long_name = "scale salt emis" ;
		scale_salt_emis:interp_method = "conserve_order1" ;
		scale_salt_emis:cell_methods = "time: mean" ;
	double time(time) ;
		time:units = "days since 0001-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "NOLEAP" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bnds" ;
	double time_bnds(time, bnds) ;
		time_bnds:units = "days since 0001-01-01 00:00:00" ;
		time_bnds:long_name = "time axis boundaries" ;

// global attributes:
		:title = "cm5_c96_am5f7c1r0_b06_piC_galb_noiceinit_alb" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:code_release_version = "2024.02" ;
		:git_hash = "b86d27037f755a82c586e55073dd575245c144b1" ;
		:creationtime = "Fri Dec  6 16:33:51 2024" ;
		:hostname = "pp211" ;
		:history = "Tue Aug 12 16:39:03 2025: ncks -d lat,,,10 -d lon,,,10 tracer_level.0003-0003.scale_salt_emis.nc reduced/tracer_level.0003-0003.scale_salt_emis.nc\n",
			"fregrid --standard_dimension --input_mosaic C96_mosaic.nc --input_file 00030101.atmos_tracer --interp_method conserve_order1 --remap_file .fregrid_remap_file_288_by_180.nc --nlon 288 --nlat 180 --scalar_field bk,pk,radon,ssalt1_emis,ssalt2_emis,ssalt3_emis,ssalt4_emis,ssalt5_emis,ssalt1_setl,ssalt2_setl,ssalt3_setl,ssalt4_setl,ssalt5_setl,ssalt1_wet_dep,ssalt2_wet_dep,ssalt3_wet_dep,ssalt4_wet_dep,ssalt5_wet_dep,ssalt1_dvel,ssalt2_dvel,ssalt3_dvel,ssalt4_dvel,ssalt5_dvel,ssalt1_ddep,ssalt2_ddep,ssalt3_ddep,ssalt4_ddep,ssalt5_ddep,scale_salt_emis,time_bnds --output_file out.nc" ;
		:comment = "FMS time averaging, version 3.0, precision=double" ;
		:NCO = "netCDF Operators version 5.2.4 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 bnds = 1, 2 ;

 lat = -89.5, -79.5, -69.5, -59.5, -49.5, -39.5, -29.5, -19.5, -9.5, 0.5, 
    10.5, 20.5, 30.5, 40.5, 50.5, 60.5, 70.5, 80.5 ;

 lat_bnds =
  -90, -89,
  -80, -79,
  -70, -69,
  -60, -59,
  -50, -49,
  -40, -39,
  -30, -29,
  -20, -19,
  -10, -9,
  0, 1,
  10, 11,
  20, 21,
  30, 31,
  40, 41,
  50, 51,
  60, 61,
  70, 71,
  80, 81 ;

 lon = 0.625, 13.125, 25.625, 38.125, 50.625, 63.125, 75.625, 88.125, 
    100.625, 113.125, 125.625, 138.125, 150.625, 163.125, 175.625, 188.125, 
    200.625, 213.125, 225.625, 238.125, 250.625, 263.125, 275.625, 288.125, 
    300.625, 313.125, 325.625, 338.125, 350.625 ;

 lon_bnds =
  0, 1.25,
  12.5, 13.75,
  25, 26.25,
  37.5, 38.75,
  50, 51.25,
  62.5, 63.75,
  75, 76.25,
  87.5, 88.75,
  100, 101.25,
  112.5, 113.75,
  125, 126.25,
  137.5, 138.75,
  150, 151.25,
  162.5, 163.75,
  175, 176.25,
  187.5, 188.75,
  200, 201.25,
  212.5, 213.75,
  225, 226.25,
  237.5, 238.75,
  250, 251.25,
  262.5, 263.75,
  275, 276.25,
  287.5, 288.75,
  300, 301.25,
  312.5, 313.75,
  325, 326.25,
  337.5, 338.75,
  350, 351.25 ;

 scale_salt_emis =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9102966, 0.8604305, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1,
  0.329, 0.329, 0.3290007, 0.3315968, 1, 1, 0.3309978, 1, 1, 1, 1, 1, 
    0.6208647, 0.3294797, 0.329, 0.329, 0.329, 0.329, 0.329, 0.329276, 0.329, 
    0.3290021, 0.3290004, 0.330379, 0.3307733, 0.329, 0.329, 0.329, 0.329,
  0.3386644, 0.3357917, 0.3389455, 0.3396149, 0.3379605, 0.3640754, 
    0.3550712, 0.4008825, 0.3609604, 0.3559966, 0.3571183, 0.383464, 
    0.3729959, 0.5966685, 0.6344737, 0.5845091, 0.5592052, 0.4601717, 
    0.5475214, 0.5538313, 0.5541232, 0.5801978, 0.5961217, 0.5794385, 
    0.3903645, 0.4029928, 0.3903408, 0.3554128, 0.3365177,
  0.6154826, 0.597862, 0.5751273, 0.5852602, 0.5833346, 0.5825846, 0.5886685, 
    0.6805927, 0.6506971, 0.6590164, 0.6883829, 0.6964859, 0.709233, 
    0.7163035, 0.7045639, 0.730353, 0.7358185, 0.7266539, 0.7136763, 
    0.6923197, 0.6860583, 0.671795, 0.6797336, 1, 0.6834327, 0.6568024, 
    0.6383022, 0.6433075, 0.5856381,
  0.7484106, 0.7501605, 0.7949758, 0.8223435, 0.7829797, 0.7724049, 
    0.7622003, 0.7516952, 0.7398153, 0.7408993, 0.7465547, 0.7594556, 
    0.8103017, 0.784839, 0.9609539, 0.7993691, 0.7903514, 0.7758853, 
    0.7637093, 0.7603381, 0.7548351, 0.753917, 0.7611391, 1, 0.7938136, 
    0.7862911, 0.7801703, 0.7643793, 0.7606145,
  0.8620348, 0.8279294, 1, 1.099958, 1.028549, 1.011317, 0.9811019, 
    0.9223393, 0.8845235, 1.044466, 1, 1, 1, 0.9854294, 0.9902083, 1.013269, 
    0.9803775, 0.9627616, 0.9714314, 1.017264, 1.044754, 0.9800581, 
    0.8855591, 0.9054438, 1, 1.05192, 0.9417324, 0.9519039, 0.918153,
  0.9676554, 1.226261, 1, 1.573946, 1.470492, 1.390419, 1.309265, 1.257113, 
    1.288275, 1.495601, 1, 1, 1.454796, 1.446811, 1.451686, 1.407355, 
    1.389763, 1.40057, 1.372461, 1.272648, 1.111311, 0.9689834, 0.9122677, 
    1.058119, 1, 1, 1.254582, 1.107046, 0.9991981,
  1.449109, 1.730362, 1, 1, 1.679766, 1.680167, 1.708227, 1.696623, 1.819634, 
    1.852053, 1.730685, 1.772489, 1.780189, 1.924791, 1.950311, 1.96034, 
    1.842463, 1.697886, 1.559782, 1.438065, 1.325435, 1.23943, 1.253205, 1, 
    1, 1, 1.527694, 1.501806, 1.418771,
  1.885194, 1, 1, 1, 1.681952, 1.846654, 1.876529, 1.965161, 1.062158, 1, 
    2.020741, 2.059572, 2.050028, 2.030409, 1.931856, 1.811471, 1.692983, 
    1.569441, 1.463127, 1.361672, 1.270097, 1.257399, 1.523213, 1, 1, 
    1.62786, 1.546755, 1.59479, 1.71973,
  1, 1, 1, 1, 1.556403, 1.742658, 1.73079, 1.810057, 1.859463, 1.791407, 
    1.773229, 1.794324, 1.782783, 1.791246, 1.761106, 1.750035, 1.733799, 
    1.723065, 1.765922, 1.761489, 1.749357, 1.718022, 1.115057, 1.500256, 
    1.662446, 1.614624, 1.55093, 1.523607, 1,
  1, 1, 1, 1.776287, 1, 1.458252, 1, 1.687797, 1, 1.553278, 1.539948, 
    1.551988, 1.544229, 1.472581, 1.425158, 1.442701, 1.422392, 1.257713, 
    1.163319, 1.222614, 1.565377, 1.332283, 1.660072, 1.629048, 1.466053, 
    1.323689, 1.232029, 1.166357, 1,
  1, 1, 1.051448, 1, 1.120371, 1, 1, 1, 1, 1, 1.014807, 1.149917, 1.062867, 
    1.03825, 0.9943351, 0.9353057, 0.9404357, 0.9489446, 0.9050004, 
    0.8518944, 1, 1, 1.046042, 1.204078, 1.16586, 1.139209, 1.043896, 
    0.9688502, 1.158291,
  0.9262565, 0.9403858, 0.8772196, 0.8883365, 1, 1, 1, 1, 1, 1, 1, 0.8088989, 
    0.7782525, 0.7361909, 0.7584515, 0.7434983, 0.7489386, 0.7622078, 
    0.7779982, 1, 1, 1, 1, 0.7574108, 0.8775922, 0.8307835, 0.8268527, 
    0.8324881, 0.8301814,
  0.723639, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9944623, 0.5308298, 0.5707077, 
    0.6004254, 0.6139314, 0.6375204, 0.6771399, 0.7158762, 1, 1, 1, 1, 1, 
    0.6412042, 0.6805701, 0.736725, 0.7472577, 0.7417752,
  0.6963347, 1, 0.5617622, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.6569986, 0.4602332, 
    0.5047401, 0.4521323, 1, 0.5046378, 1, 1, 1, 0.9683141, 0.4370593, 
    0.9520392, 0.5492584, 0.5789813, 0.6917861, 0.715255, 0.7130584,
  0.4766365, 0.6180748, 0.4473523, 0.4517508, 0.4095937, 0.348612, 0.3941887, 
    1, 1, 1, 1, 0.9372528, 0.7757074, 0.4311774, 0.3912068, 0.3561752, 
    0.4353301, 0.4016452, 0.3700163, 0.3465343, 1, 0.3650447, 0.4138954, 
    0.6497492, 0.4050392, 0.9794201, 1, 0.3490314, 0.3629941,
  0.329, 0.329, 0.3323479, 0.329, 0.3298017, 0.330596, 0.329, 0.3293555, 
    0.3296299, 0.3318305, 0.3290766, 0.3314459, 0.3325869, 0.3351538, 
    0.334858, 0.3332629, 0.3304953, 0.3364313, 0.3375536, 0.3352008, 
    0.3298441, 0.344496, 0.3550921, 0.3309542, 0.6685761, 0.9744557, 1, 
    0.4219843, 0.329 ;

 time = 912.5 ;

 time_bnds =
  730, 1095 ;
}
